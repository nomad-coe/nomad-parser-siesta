H   F�`)�Z#@                        ���+BY@                        I�p�^+@H      6       P         �   ��F=�0=\�<�@<P�P��z>��Fx�@�������1����Fx��z>�dO�X�X@<�]�<^�0=��F=�h.=��<�A����½ЮT�.k��!S��1j��-����%���6�YKb�sZ��bС�X����C��*���D�������С��Z��DLb���6��%�࿿.��h3j��T�=m����T�܇½�L���<�e.=�   �   ��0=��=�0�< �9������5��s��cn��$跽3���跽Hn���s��P�5����� C�9�2�<��=��0= �=䎛<O��F���]OP�h���rc�cf��Z���hܿ���!�3�O�]��o���*���y�����������Hz��+��!p��2�]��3�U��jܿ�[��!f��d�q���BRP�Kž�,Z��<��<^�=�   �   TM�<h�^<��ڱ�7���#�������;:��� �2:����}��m#�����������^<�P�<8B�<x�V<ٽ��;��_�C�����+����Y�9"���ѿ���΢*���Q��s|�ؓ�*���!�����:!��|����ؓ�et|�_�Q���*�R��7�ѿ;#����Y�w��袰� �C��?���㽼�V<0=�<�   �   �w�Eμ��m�Lǽ�v���8��^���{�󅇾�Ҋ�텇���{��^��8��v��ǽ��m��Bμ�A��K<�!;��μ�.��X�0�������F�?:�������O�����LZ?��Rd�����i�������}���ǰ����������Sd�[?�d���P�� ���.;����F�L��䶟��0�U2����μ � ;HB<�   �   (X5�T`B�j�C�k0���🾸r��1<Ѿ�9߾���9߾&<Ѿ�r����U0��6�C�$B����V5�������f�,���'��H�������侠�.�r{�R|��B#߿ϟ��`)�!H���e����ٸ���݋�������< f��H�ra)�b��T$߿J}���s{��.���4������Y
��<���X�f�l����   �   )�ҽ��&�$4s��ꤾЇҾL���U��"��-�:|0��-��"��U�5����Ҿ�ꤾ�3s���&�^�ҽ�w��k��[�OǇ��A�jg����]�t�U������>�����͵�`�*��NB�V�yjc��&h��jc�qV�3OB���*�N�����|?��������U��^����,!g��C� ʇ��_��n��w��   �   4|8�����.^��5�����x >�J�Y�QZo�.}����.}�HZo�<�Y�i >������^��v����{8�k�r�����Y��I���Խ�8��5���h�T�.�<;r������ɿ�b�S#��� ��/�2�9��=�T�9�]�/�� ��#�uc��ɿ�����<r���.��j�g7��h�8�b�Խ;L���Y������k��   �   _M����; ����6�]b�݅��2��뉦������Ͳ�����剦��2��݅�Ib�t�6�	����;,M��Ez9�z�罄e������7�� I��j�,(��|��T?��~�@���+�ĿZ��Ϣ��L�(��=q�B���L������ۄĿ򠡿@�~�V?�}��)����j�K�������g����罺z9��   �   K�ʾ�3�67B�c�x�8���m@����ʿeݿD�����@��^ݿ�ʿb@��*���I�x�7B�y3��ʾQ����I*�V/ӽ'Γ��̓�=*ӽE*�����0�ʾ60��2B�A�x�:���=��L�ʿ�ݿH�����p���ݿ��ʿ�=��ǀ��^�x�4B�(1���ʾ"���G*�F-ӽ�Γ��ϓ��0ӽJ*������   �   �~��X?���~����x�Ŀ��٤��N�j��|s�g���N�Ӥ���h�Ŀ	�����~��X?��~�3,��q�j�XL�������a��6�罔t9�I��&�;���%�6�4b�1څ�j/������7���kʲ�W���Ɔ���/���څ�b��6�Y����;XJ���v9�X��5d���s	���L��j�p,���   �   ��.�X?r�<����ɿ f�T%�פ ���/�ř9�w=�9���/�Τ �K%�f��ɿ*���6?r�b�.�im��8����8���ԽfJ��ĐY�����b�_u8����dX��������>���Y��To�F(}�%�x(}�Uo�{�Y�=>�b�_����Y��-���7w8�!e�a�����Y��K��
�Խd�8�"9���m��   �   ��U����A��񿜷��*�:QB��V�hmc�x)h�dmc��V�0QB�t�*������A��������U�`�L���"g�D��ȇ�Y�*d�"w���ҽ��&�:+s�R夾E�Ҿ�����Q���"�3-��w0�X-���"��Q�����4�Ҿ@椾�,s���&�E�ҽ�w��g�\�ʇ��D�	#g����9`��   �   Pu{�X~���%߿K���b)�RH�Hf����j���ߋ�g������;f�DH��b)�=���%߿@~��'u{��.�� 便������8	�����H�f��o��(H5��㩽�;�V}C��+��&럾�l���5Ѿ�2߾0�,3߾�5Ѿm���럾G,���~C�=�1橽(L5��v����f�����C
��4������;!��.��   �   �;�������Q�����[?��Td� ���Ը�����씣����͸�������Td��[?�	���Q�������;��4�F����"���˰0�$1���μ�F!;0e<@�T'μ,�m�ǽOp�|8��^���{�G���'Ί�i���c�{�A^��|8�>q��ǽ��m�,.μ@e꺸Z<�"!;�μ2��8�0�\������Z�F��   �   w#����ѿ����*��Q�Vu|�-ٓ�Q���4"��"���0"��J���$ٓ�@u|��Q��*����{�ѿ_#����Y�v��������C�B>��$ܽ�X�V<�I�<@]�< �^<H��v��������+����v4�"� ��4����2��X��/���D��x��h�^<�X�<xE�<�V<T߽�?�� �C����������Y��   �   �[��jܿT����3�W�]�Gp��S+���z��<��N���8���z��I+��<p��C�]��3�C���iܿ�[���f�pd�˝��0QP�gþ��R�����<��=��0=H�=>�< ��9P䵼�5��n���h���ⷽ���ⷽ�i���o���5��赼 ��9`9�<�=��0=��=`��<�U��%ľ��QP�����d��f��   �   D.����s%�m�6��Kb��Z���С������C��)����C�������С��Z���Kb�Z�6�b%�m�+.��q2j��S�l���T�u�½�E��x�<8h.=��F=��0=4_�<�@<����M��y>�Fx���������K���.Gx�Z{>�`Q��@@<�Z�<��0=��F=zf.=X�<�H��-�½~�T�Ul���S��2j��   �   [��iܿ���)�3�@�]��o��i*���y�� ��.�����y��_*���o��,�]��3�����hܿ[���f��c�ǜ���OP������N��l��<\�=�0=��=`>�< ɋ9,䵼�5��n���h���ⷽ���ⷽ�i���o���5��赼 ��9�9�<n�=�0=��=$��<�Q��l¾�>PP�����c��f��   �   "��Ϸѿv��v�*��Q��r|��ד�^��� ������ ��V���wד��r|��Q�e�*�g����ѿ"����Y���ʠ��	�C��:���ӽ��V<M�<L_�<��^<���F��������2��&��~4�+� ��4����<��\��*����� ����^<�Z�<�H�<��V<׽��;��s�C����)����Y��   �   �9��I����N����aY?��Qd�ڠ��L���R������N���E���Ҡ��uQd�QY?����N��0����9��b�F����s���C�0��,��h�μ �!;�n< �麜%μ��m��ǽHp�|8��^���{�M���+Ί�p���l�{�H^��|8�8q��ǽZ�m�p,μ 8��c<�]!;X�μ{-����0����������F��   �   �p{�`{���!߿����_)��H���e�1��k����ۋ�i���&����e��H��_)����!߿H{���p{���.�A侎���������������f�Tj���F5�i㩽�;�H}C��+��'럾�l���5Ѿ3߾9�63߾6Ѿ m���럾D,���~C��<��婽�J5�8q��P�f�ؖ�������ʦ���侲�.��   �   ��U���=����𿍴���*��LB��V��gc��#h��gc��V��LB���*��������<���󒿞�U�q\�4
���g�w?���~Q�^_�&	w���ҽ��&�+s�I夾B�Ҿ�����Q���"�7-��w0�[-���"��Q�����1�Ҿ8椾�,s�@�&�^�ҽ�w�$c��T�'ć�@�,g�s
���\��   �   z�.��8r�����ɿ`��!��� ��/�Ɣ9�U=�Ô9��/��� ��!��_��ɿ�����8r�Y�.�f��3����8���ԽsD���Y������`��t8�����QX��������>���Y��To�K(}�(�|(}�Uo��Y�?>�a�V����Y������v8��c� ����Y� F����Խ��8�4��Vf��   �   -z�\R?���~�+�����ĿY�����J���o����J���J�忓�Ŀ�����~�<R?�z�P%���~j��E�V���`���'^������s9��H���;�� �6�3b�2څ�j/������:���nʲ�Z���Ȇ���/���څ�b� �6�Q��~�;$J���u9��罗`��I���� ��lF�Xj��%���   �   ��ʾ�-��/B�[�x��}��F:���ʿ�ݿ������|���ݿ�ʿ<:���}��?�x��/B��-���ʾ'����@*��#ӽDƓ�YǓ��&ӽ D*������ʾ)0��2B�>�x�:���=��N�ʿ�ݿL�����t���ݿ��ʿ�=��Ȁ��]�x�4B�1���ʾ����F*�*ӽ�ɓ�ȓ��$ӽ~A*�a����   �   F��
�;�����6� b��ׅ��,��p���褯��Ʋ�夯�i����,���ׅ��b���6������;�E���o9����W[������� ���G�,�j��'���{��T?��~�>���,�Ŀ[��Т��L�)��?q�D���L������܄Ŀ򠡿=�~�
V?��|��)����j��I����ͥ���\�����;p9��   �   \p8������S��`���= ��>�A�Y�uOo��"}�D񀿱"}�jOo�3�Y�p>�* �<����S�������o8��Y�=�����Y�D��M�Խ��8��5���h�G�.�8;r������ɿ�b�S#��� ��/�3�9��=�U�9�^�/�� ��#�tc��ɿ�����<r���.��j�7��D�8���Խ�F��*�Y������Z��   �   ��ҽ��&�9$s��ा�{ҾF����M���"���,�s0���,���"��M�/����{Ҿ�ा�#s�J�&�ΰҽT�v�zX�N���B@��g�����]�l�U������>�����͵�`�*��NB�V�|jc��&h��jc�sV�4OB���*�N�����{?��������U��^����G g�BB��Ň�R�f[�p w��   �   B<5��۩��6��vC��'��\柾g���/Ѿw,߾t��q,߾/Ѿ	g��J柾�'���vC�\6�V۩��:5��Y��(�f�t������,��J����侖�.�r{�R|��B#߿ϟ��`)�!H���e����ٸ���݋�������= f��H�ta)�b��U$߿K}���s{���.���㨊�t����������f�$^���   �    ��tμ��m�	ǽ�j�|u8�^���{��|���Ɋ��|��x�{��^�_u8��j��ǽ��m��μ���؆<��!;�|μG,����0�㴟�
���F�>:�������O�����LZ?��Rd�����h�������}���ǰ����������Sd�[?�d���P�����.;����F�>�������0��/��Ȇμ��!;8}<�   �   �f�<_<������ ���$������/�}� ��.� ����������̗�(��8
_<@j�< U�< �V<XϽ�J:����C�נ��#����Y�9"���ѿ���͢*���Q��s|�ؓ�+���!�����:!��|����ؓ�ft|�`�Q���*�R��9�ѿ<#����Y�q��Ƣ����C�%>�� ڽ�0�V<(P�<�   �   ��0=��=�D�< �9�ص���5��j��Hd���ݷ�i뾽yݷ�3d���j����5��׵� [�9�F�<��=��0=��=���<LJ��{���#OP�X���nc�bf��Z���hܿ���"�3�O�]��o���*���y�����������Hz��+��!p��3�]��3�V��jܿ�[��"f��d�`���RP��ľ�pU�����<�=�   �   ��I=�4=h��<اT<�}廀,ۼ��5��Hn�������a����l���2�tԼ`\ƻ��d<.l=�8=N=r6=�׼<�֟��A����N��纾h
�u�e�.���ܿ*��ɂ3�.�]�f��G5���V���������o���`a��㪆�yh^�z&4���� ݿ@ѣ���f�����#��$~P�.@���ש�P��<��1=�   �   �T4=l�=$r�< 7�:@觼�g-��}�|❽0α�1q���)������h�y�n�)�\ȟ� �/;DԹ<��=�k8=��'=X��<�������_TJ�T.���*�Ba�UU���}ؿ,>�q0��Y�ۘ��̯����������uI�����������͚��σ��"Z�1�����Xٿ�����b�C��x^���(L�����TҪ��դ<�h#=�   �   (��<�r<0�׻^&��~�혹�:�w2��9�W��V���~
���뽷l��r(z��}�P?���<xQ�<��< �{<����W���>��o��<���U�J��hοֈ�~�'���M��gw����������<��;���!*��������w�+N�V(����:�οlؘ�0wV�̈���0�?��������j<���<�   �    �ȹ�W��>e�C����!���4��{Y�r�v�����ȇ��h����u��JX�W+3�ڹ	���b`��̶� �5: 4<���;\���Ѯ��~f+�<���������B�K�������0+��n2��<� $`��	��W���8L�����?*���w�������_�m<�IX�����"��
��p�C��v �ￜ�g�,����pG��@�{;�u#<�   �   �>-�B㤽��?�Qs}�������Zc;D۾��߾��ھ��̾�;��8���{�|�=�]���5��ڐ(��U�� v<��ݼ���}���C��F߾>+���v�����Ñۿ�r	�ֵ&���D�z�a���z�z�������ׅ��wz��na��jD�r�&��d	���ۿ�Ȩ��^w�a�+���'쇾+������u��L�T����   �   �ͽG#�ȅn������ξ���S��,; ��*��M-���)����Q�"���C�;&頾n�l���!�0�ʽʪi�`��D��[)���
���Ja�7�;��&R�F����=��he�6���<(�WB?��{R��Z_���c��_�r�Q�p�>��'��;���^������5:R�����c���)b�.����Ȃ��
��C���m��   �   w4��H��L���~�A$;��FV��k��	y��}���x���j�r�U�RT:�����Q���黾���"3��:܉�xrM�n
v���ͽ�4��ؕ����+�9n�.���(ƿ���$�R��-��6���9��Q6���,�������.ￚ�ſ᜿�m��{+�.��R���4�n�νtbx��$P�}���,��   �   態��Nʾ8z
��3��^��߃��������x꯿���ߛ��_j���T����]��3�<�	��Zɾ�׊��O4�		ཽ命�8}�)u���=
�m#e�Q�����@$<���z�==��(���ڡ�§���C�a����$\���
��������&��ﴞ��y��;���,F��ve�S
�\稽�~�-ܒ�xb��D5��   �   D;Ǿ���>?��3u��K�������ǿ��ٿ^W�J&鿵忥Sٿl&ǿ ������M9t��f>��A���ƾ�˃���%��̽�̍��ہ̽�&�/-��>6ǾV��?��.u��H��L���v�ǿ��ٿqS�b"����'PٿF#ǿH���,���r5t��c>��?�c�ƾ�Ƀ�'�%�~̽n͍�F�*�̽�&��0���   �   a
�(<�4�z�@��h������ȫ���E�����
�>^���
������Ῡ������F�y���;�����H��Qe�UT
�[稽�~�ג�2Z��>5�����Iʾ�v
���3�У^��܃��핿���-篿̱��͘���g��3R����]��3���	��Vɾ�Ԋ�L4���n䑽l;}�My���A
�<)e������   �   �+�=n��0���+ƿJ���%�RT�e-���6�m�9�<T6���,�j��9���0￬�ſ�✿��m�]}+���������4�ލν�^x�zP�[v���"�Gp4������B����y�;��AV�\�k�*y�U�}��x���j��~U�:P:����&L��K廾j���3�I�-ى�tqM��v���ͽ�4��ە�����   �   cR�U���*@��hh����?(��D?�Z~R��]_���c��_���Q�b�>���'��<�����������;R�����d��J+b������ǂ�H�v9���m�ͽ1@#��|n�����/�ξ����8���6 �C *�vI-�X�)�����M�����ܼ;�䠾��l��!�2�ʽ�i�b������+����@Oa���������   �   ��v�񛨿,�ۿt	���&���D��a�d {����f���Vم�zz��pa�lD���&��e	�Ϩۿ�ɨ��_w�H�+��	ྮ쇾V������k�8�K����/-��ؤ��
� {?��i}�h������\;��ھ�߾�ھ��̾86��w���{��=�]���.����(��I��8m<�P�ݼ)���Z��7F���I߾@+��   �   ����ʦ��`-���3��<�&`��
�������M��.���+���x��������_�W<��X��������
����C�w �,���O�,���� ?��`�{;0�#< �¹,:���+e�(����~~4�SsY���v�����}Ç�Cd��p�u�:CX��$3�a�	��羽�`�p����M7:�-4< ��;����	���Li+�n⛾3�����B��   �   <K���ο�����'���M�Riw����������=��J���+����������w��N��(����}�ο�ؘ�NwV�ʈ��~����?����\�� �j<��<���<@�r<�?׻"�r�~������t��,�64��������y
�}���d��z�s�0�����<�X�<$�<��{<PƦ��Z��`>��q�����ӖU��   �   @V���~ؿ�>��q0��Y�v���{���m���\���J��2�������͚��σ��"Z�1�y���Xٿ���R�b�����]���'L�����,˪��ܤ<�l#=VY4=��=�< '�:ק�|^-�B}�ݝ��ȱ��k���$��筜��y�J�)����� �/;�ڹ<�=�l8=4�'=؝�<h��蚶��VJ��/��,���a��   �   ����ܿ���7�3���]�Xf���5�����o�� ������?���"a�������g^�&4�W� ݿ�У���f�+���"���|P��=���Щ����<(�1=��I=�4=x��<�T<�r�*ۼ��5�Hn�������z���0l���2�XԼ�eƻ��d<�j=8=@N=N6=�Ҽ<lݟ��C��e�N��躾*�j�e��   �   �U���}ؿ@>�%q0�ږY�������g���F����H���������͚��΃��!Z�J1�����Wٿ���D�b�%���\��8&L�����ƪ��ߤ<�m#=�Y4=N�=|�<�*�:�֧�|^-�J}�ݝ��ȱ��k���$����y�N�)�������/;,۹<Z�=(m8=�'=���<4���=���9UJ��.��]+��a��   �   �I��,ο���(�'��M��fw�븐� ����;��-���)���ߢ� ���U�w��N�7(������ο6ט�IuV�^���|���?�h
���
����j<t��<��<��r<�<׻��P�~������t��,�<4��������y
�����d��z��r������<�Z�<L�<��{<8����W���>��o��:��ԔU��   �   ޥ��_���P*���1�<��"`����D����J��d���(��rv���ށ���_��<��V�ʑ��T�����4�C�u �������,����l3���'|;��#< *¹h8��,+e�����y~4�UsY���v�����Ç�Hd��}�u�BCX��$3�`�	��羽F`�趶���7:�64<PϞ; ��������e+��ߛ�M���/�B��   �   ~�v������ۿ�q	���&�b�D���a�$�z���f���oօ��tz�Vla�nhD��&�<c	��ۿ�ƨ�W[w���+��྇釾.��4����]开�K�x���j--�mؤ�i
�{?��i}�g������\;��ھ�߾"�ھ��̾>6��|���{���=�>��.���(�LD��8\<���ݼ����>��C���D߾3=+��   �   }R�#���%<��xc����n;(�j@?�YyR�+X_���c�_���Q��>��'��9�� �����~���6R����_��}$b�Ŭ����������4���m�) ͽ�?#��|n�����)�ξ����;���6 �F *�zI-�]�)�����M�����ڼ;�䠾��l���!�U�ʽ(�i����T��6&��B���Ha������   �   !�+��6n�x,���&ƿK��x"�FP���,���6�k�9�^O6�8�,�a������*￦�ſ�ޜ���m�fx+�b�������~4�քνSx��P��s��p!��o4�m|���7����y�;��AV�^�k�.y�[�}��x���j��~U�<P:���� L��:廾K��)3����։��iM��v��|ͽ�4��֕�q���   �   ���!<�A�z�0;��������U����A�H��]��Y���
�����,��� ��$���U�y���;�#���A����d��M
��ި���~�gӒ��W�">5�}����Hʾ�v
���3�ͣ^��܃��핿���.篿б��И���g��4R����]��3���	��Vɾ�Ԋ�iK4�������J0}��p��8;
��e��}���   �   �2Ǿ��?��*u�SF������R�ǿ2�ٿ�O忄���^Lٿ�ǿ����?���i0t��_>�5<�9�ƾ�Ń�-�%��̽�č��ꍽ�~̽�&��,��6ǾH��?��.u��H��K���v�ǿ��ٿtS�g"����+PٿH#ǿK���-���r5t��c>��?�>�ƾIɃ�.�%�J	̽`ȍ��덽�|̽&��*���   �   �~���Dʾ t
�L�3���^�kڃ��ꕿ����ꬿ�㯿h���}���vd��WO��u�]�C3�
�	�QɾwЊ�eE4�u�߽�ۑ�0+}��p��x<
��"e����m�5$<�|�z�<=��(���ء�ħ���C�b����&\���
��������(����y�y�;����E���e��Q
��⨽��~�1Ғ��SὋ:5��   �   Uk4�6놾&�������fv�g;��<V�6�k���x���}�b�x�H�j��yU��K:�e��%E���߻����x3�&�*Љ��aM�"�u�}ͽW4�(ؕ�����+��8n�.���(ƿ���$�R��-��6���9��Q6���,�������.ￛ�ſ᜿��m��{+��������4�͉ν@Wx��P��p�����   �   <�̽�:#�vn�0���ξ�������2 ���)��D-�ݿ)�����I�[z��u�;`ߠ�ˠl�д!��vʽ��i�<�����$������Ia���)��R�D����=��fe�5���<(�WB?��{R��Z_���c��_�u�Q�q�>��'��;���^������/:R����ac��)b�L����Ă�T���0��m��   �   L#-�Ѥ�p��t?��a}����������V;$�ھC�߾{�ھY�̾A0������{��=��~��#��Xu(�-���;<�t�ݼ����b���C���E߾>+���v�������ۿ�r	�յ&���D�y�a���z�{�������ׅ��wz��na��jD�s�&��d	���ۿ�Ȩ��^w�Y�+�l��뇾��K��La�@�K�|����   �    ־�l$���e�>�����x4��kY�]�v����������_����u�;X�z3��	��ܾ� �_�̙���y::Y4<@�;����Z����e+����������B�J�������1+��m2��<� $`��	��W���8L�����@*���w�������_�o<�IX�����"��
��l�C��v �������,�=���8��@0|;��#<�   �   <��< �r<��ֻR�4�~������k��'��.���P��Qt
�M�뽎[���
z��d�P���P&�<|j�<�!�<H�{<����:V��Q>��o��2���U�J��iοֈ�~�'���M��gw����������<��;���"*��������w�-N�X(����:�οnؘ�0wV�ň��~����?����T����j<���<�   �   �Z4=H�=腱<���:�˧��W-�2}��؝��ñ��f���������y��)�����b0;��<��=�q8=$�'=��<���Q���%TJ�E.���*�@a�UU���}ؿ,>�q0��Y�ۘ��̯����������vI�����������͚��σ��"Z�1�����Xٿ�����b�?��j^��e(L�̂���ͪ�4ܤ<@m#=�   �   V�V=*�A=�=���< ׺Tm����O��q�x�{���n�F�J������� ��9Ă�<�=�OJ=ns_=BrH=���<x2J�4��&�>��	��V��YY�Yޚ�feѿ׭��x*�y�Q��|�-��F��ͳ��<���ҳ��6��zv���}�,�R�D�+���cӿ�(���V[�9��=Z��UnB�n����r�0X�<X�?=�   �   VB=�}%=���<`9�;��n��`�z�]������n���x��)���;���W��	��{M���<{�<@;.=�J=؆:=�)�<��L�����^�:�K���4��htU��=����Ϳ��j�'�Z�M��w�-����U���������I����`���(���[x��N���(�;e���Ͽ�s��
WW�������0E>�pr����t����<��1=�   �   67=<��<�У���ۼ�x_�e����ؽ�����7�03�Uz�����5սe���%V�вȼ�L�:83�<�=�=��< uX�b����/�Q�����d J�����Ŀ Y��%u�m C�iSi�����������������y����އ�d�i�)�C�N �k���Aſ����K�����P��U2�?a��ب~�dE�<��=�   �   �s�;����G��F�� �7�'���J�'�f�%x���}��6w���d�ǄH���$�'����Ω��<�X�v��e�;,~�<�2<��y�*'���o�f������f8�!����r��/��=��_�2�"T��u��Ԉ�����(��dS������t�C�S�پ2��!��F뿄4��.>��%�9����}D���4 �/���������<�Ip<�   �   *L���������12��Xm�@���L��ڕ��pxξp�Ҿm�;�q���˫�"ܑ���i���.���R��4����,��j���<��L�v���R#|���Ѿ�!�#?j�:a���Bѿ��N����:���U��l�1^|�Ԁ�l�{�A l�>U��T:�v����hѿv����k�F�"��`Ӿ��~��?
��~�����߻0`O��   �   �����&�(_��\��!Iþ�r!	�����!�$��� �}�������,��.X��V�[��,�����F��fἔ����^����7Q�qy���r��!G��a��0O��Q��|	��_ �q�5�ڹG��S�YqW��R���F���4�_���k�|������Z���\G���L���R�]E�6ae�P\��l4���N��   �   &z'�>�|�&'���쾝P�@�1�R�K�_�_���l���p��l�ʸ^�*%J�, 0����������y�z�$��ɽ}o�0�,���S�*ָ�uH&��:��^Sܾ�k"�69b����������|������$���-��0��C-�$�;�.�����������a��<"��bܾI����&'��亽�tX�,2��v��ν�   �   ł��¾�O�ާ*���S��{��͎�zD������2}��~P��*���~܍��y�*�Q��#)��������x���;&�{Xʽ0��\D[�ɕ���adU�p���wE���d2��Wn�:���"۸��lؿ,�����	����r��F������ֿ^���p����
m�&�1��]��J6���$U��l��1���
 ^��с��ͽ(��   �   �������[5��2i�{-�����������Ͽ��ڿ Q޿�8ڿq�ο�w���E������mg��4�Y4��}����u�}��Ƿ���x�}y������\�]Fw�檻�d��W5��-i��*��t���D���p�Ͽ��ڿEM޿h5ڿ�ο�t���B������ig�
4�+2��z����u��z��ŷ��x�\�y�����ma�NMw��   �   �J��Oh2�	\n�츗�B޸�Apؿ�/�����$����	t�bH������ֿǕ��kÖ�m���1��`���8���'U�:o��3���@�]��́���̽H(������������*�̞S�&�z��ʎ�FA��=����y��VM��:����ٍ�By�2�Q�Q )�Q��M���
v��f8&��Tʽ����F[�͕�,&���iU�m����   �   �n"�=b�쥕�f��;�\������$��-�X�0��E-�$������V����r��B�a�M>"�4eܾ����5('�J庽`qX�\2���u�<�ͽ�s'���|��!���쾠L���1�M�K��_�2�l�B�p�v�k�ٳ^�� J�C0����������_�y�*�$�x�ɽ2wo�:�,���S��ڸ�vL&��=���Wܾ�   �   �$G��c���Q��.��+	��a ���5�U�G���S��sW���R���F�v�4�ن��l�]��b���[��{^G�(��oM��U�R��E潮^e�P��H �"�N�����` ��_�|W���Bþ�	����L� ��$��� ����E������T����[�.(�b���6|F�_�t����^���B<Q��|���t��   �   &Bj�c��2Eѿ*������:�Q�U���l��`|�fՀ���{�sl�U�V:�#w�����iѿ`���Jk�$�"�bӾ��~��?
���~�������߻x3O�=�3�������7*2��Om����IF������	rξ
�Ҿ>�;�k��Pƫ��ב��i���.�0��lK��p����,��Y���?���v��	��'|���ѾU�!��   �   �����t��C��}���2��#T��u��Ո���q���T�������t�p�S���2�F"��G�#5���>����9����D���4 ��������0�<(kp<@̚;�厼G�/<��� ��'���J���f�Gx���}�'.w���d��}H�X�$������Ʃ���<���v����;<��<X2<�z�8*���r�}������h8��   �   B���3Ŀ�Z��0v��C��Ti����ħ�����������3���4߇�,�i���C�� �׫��JAſ>��� �K����oP���T2��_��X�~��N�<��=�>=�<@`����ۼ�h_�\����ؽ����U2��-�!u�	���,ս����V�T�ȼ@I�:�>�<�=��=��<؀X�]���/��R��R��3"J��   �   u>����Ϳ���)�'�D�M���w�����*V��7���s	������a��()���[x�'�N���(�,e�v�Ͽ�s���VW�]����)D>��p����t�$��<��1=�B=��%=p��<�s�; �n��W��~]�s����i���s��9$��Y7���	W��	�8eM�H <d��<6=.=�J=��:=8&�<x�L�F���l�:�ς��B���uU��   �   �ޚ�	fѿ3��8y*��Q���|�M-��s��ͳ��<���ҳ��6��Bv����}���R�ߑ+�����ӿW(���U[����*Y���lB�$	���r�x]�<x�?=8�V=ޱA=>=h��<@�ֺ k����^O�`q�V�{�ܦn���J�@��𿙼 5�9T��<~�=NJ=�q_=<pH=���<�?J�� ����>��
���V��ZY��   �   �=����Ϳ��s�'�P�M���w�����8U��/���c������`��T(��wZx�(�N�<�(��d��Ͽ�r���UW���$����B>��n��0�t����<��1=pB=Z�%=���<pt�;��n��W��~]�v����i���s��B$��`7���	W��	��dM�` <���<�=.=h�J=T�:=�(�<h�L�����0�:�ہ������tU��   �   �����Ŀ�X���t���B��Ri�&����� ��	������p����݇�ȓi�ڄC�> ������?ſ𒑿�K����N��)R2��\���~��S�<��=�?=p�<@R���ۼ�h_�\����ؽ���X2��-�*u�	���,ս����V��ȼ S�:�?�<�=2�=� �< qX�J����/�*Q�����N J��   �   ����Ar��Z�꿧����2�� T� u��ӈ�w������R�����ĉt�^�S�N�2�e ��D��2���<���9����,B��C1 ���L�����<�tp<�ך;�㎼~
G�<��� ��'���J���f�Nx��}�4.w���d��}H�[�$�����mƩ���<���v���;h��<�2<��y��%��]o�����1��f8��   �   �=j�V`���Aѿ �D��o�:�:�U���l��[|��Ҁ���{���k��U��R:�it����jfѿ�����k��"��]Ӿ�~��;
���~�P��d߻`(O�J;�����/���*2��Om����JF������rξ�ҾF�;�k��Vƫ��ב�
�i���.����K�����X�,�9���2����v����!|�[�Ѿ/�!��   �   A G��`���M��x��R	�6^ ���5���G��}S��nW���R�[�F�o�4�n���i���῀���X���YG�����H����R�?=�^Se�\A����(�N����� ��_�nW���Bþ�	����N� ��$��� ����I������ T��Ǝ[��'�����vyF�,V�T����^�d���5Q��w��qq��   �   j"��6b���������~���+���$���-���0�DA-��$�,�T�����2��|����a��9"�O^ܾℌ��!'��ܺ��eX��2�"�u���ͽ?s'�l�|��!���쾛L���1�N�K�	�_�4�l�E�p�}�k�߳^�� J�F0����������*�y���$�!�ɽ�ro��,���S�LҸ�F&�9���Pܾ�   �   �A��Xb2�nTn�B����ظ��iؿ�(����������o��D����ֿH���þ��zm���1��W��2���U��b���^�]�NɁ�e�̽�(�����p�������*�ǞS�#�z��ʎ�GA��>����y��[M��=����ٍ�Gy�3�Q�P )�L��7����u���7&�zRʽ���@<[��ĕ�����`U������   �   ����-��T5�A*i�e(��ˁ��?����Ͽ<�ڿ�I޿�1ڿy�οaq���?�����eg�4��.��u��0�u��t�b�����x�"sy�{����[��Ew�����U��W5��-i��*��r���D���p�Ͽ��ڿIM޿l5ڿ�ο�t���B������ig�
4�#2�mz�� �u��y�y·�`�x��ty�����UY��Aw��   �   <�������]	�w�*�њS�t�z�2Ȏ�T>������v��J��}���֍��y�_�Q�4)�����＾�q���1&��Jʽ��R7[��ĕ�N���cU�,���PE���d2��Wn�8��� ۸��lؿ,���������r��F������ֿa���q����
m�"�1�v]��6��*$U�j������$�]�+ȁ���̽((��   �   �n'�H�|�w����OI�Ɠ1��~K��_��l���p��k���^��J��0������l����y�^�$���ɽ�eo�.�,��S��Ҹ�RG&�q:��*Sܾ�k"�-9b����������{������$���-��0��C-�!$�=�/����������ݮa��<"��bܾ�����%'�]ẽjX�,2���u�I�ͽ�   �   R� _�ES���=þ��	����%� �$�k� �q��h�����
���N��q�[�j!����jF� B���*�^����7Q�.y��yr��!G��a��.O��M��{	��_ �q�5�ڹG��S�ZqW��R���F���4�`���k�~������Z���\G����K��,�R��B潠Xe��B��p���N��   �   �1����������#2�9Hm�����A������kξ��Ҿ��;�e������ґ��i��.����BA����Ȱ,�0����(����v����"|�U�Ѿ�!�?j�7a���Bѿ��N����:���U��l�2^|�Ԁ�n�{�C l�@U��T:�v����hѿu����k�>�"��`Ӿ\�~��>
�z�~��� U߻�O��   �   �
�;�Ў���F��3��� ���'���J��{f��x�R�}��%w�L�d��uH�N�$�^���򻩽<�<��v�0��; ��<*2<p�y��$��9o�.������f8�����r��/��<��^�2�"T��u��Ԉ�����(��eS������t�D�S�ھ2��!��F뿅4��->��!�9����ID���3 ����������<�p<�   �   JC=��<�Z��Ȅۼ\_��T��a�ؽr���5-�z(��o�����*#ս���D	V�,�ȼ ��: R�<�=�=�)�<�bX�����!/��P�����` J�����Ŀ Y��$u�l C�iSi�����������������x����އ�f�i�)�C�O �m���
Aſ����K����vP���T2��_��x�~��R�<��=�   �   4B=*�%=���<@��;�n�"Q��v]�����d���n��$��\2�� W�J�	�HEM��<��<�B.=�J=<�:=0�<��L�ҧ��$�:�<���0��dtU��=����Ϳ��j�'�Z�M��w�.����U���������I����`���(���[x��N���(�<e���Ͽ�s��
WW��������D>��q��x�t�l��<.�1=�   �   �_k=��W="^'=ls�<�&�;0a.��"׼$t���<��F���8������ü ����&<��<��5=Jf=��y=�qd=��=�����ׄ��&�Q䜾���F�2������c�������?��6e��i���ו�����������������2<f��A��:�\�����¿�ԏ�,I�������+��Ǎ�����b�=κU=�   �   ��W=@==��= �p<���ɼ-+��Qb��e��E����}��P"[��>!�X���2򺨔�<B=
�K=Ff=^cW=^=@V̺9����"�F���G���7�B���ѽ��e���a��o<���`�訂�����p��7F���j������6���&�a��=��������2���L��`E�k�2����(�k������D =8�H=�   �   LT=l��<��;�@���H-�HL��8&��Kܽ���˒���h��׽������������R�p4<@��<&�*=�;/=(��< ��<�q�Z?��H��+s�@y8�����M����������2�H�T���u��U��c1����������-����u�9�T�X�3����b������:����G�����(����û���<�� =�   �   `\S< ���Է�����h�ܽ4��~3�-M��]��8b���[�<�J��40�O �z�Խ?v������[����<0�<���<`U��vhX����ہ���پ�(��s�#��;�ؿ��~$�
)B�	�^��{w�.��c����փ�y�v��;^��A��$�\���gٿj���t���)��ܾ)����`g����`�<$׵<�   �   ��ȼ�p�Iҽ���3�S�P|��=���鮾L����{���߹�\��?,��� ����N��.0ɽ0�_�(#�� t�8 }�;Й�D�=���V�_�Bl��JQ��vV��������;�Ә�*,���C���W��'e���i�-�d���V��B�m;+��+�l��cE���铿fvW�`T��S���Kc��<�tJ� .?� �;``U��   �   L���J���nF���������eL׾2����K
����͈��=�C	�M���jKԾǩ��y+��gA����������P(���ӈ�J#(��h��MX8�����������5��K|� /��	Eѿ:X��	���'��[7�!�A�E�,A�mF6�-]&�������pп{ԥ��9|�D6�X����͞��:��3Ľz2�h靼@O������   �   �����a��Π��o־+;��]"��a:�B&M���X�/�\�30X��K�x�8�1k ��X��Ӿ2󝾾K]�x���ϧ�N�7���� ������D��9|z�3LǾ���AO�|���ge�� �ӿ����,��')��& ���"�{��6+��|
�js��^"ҿ�A������ΏN�����`ǾQ{�*�KÛ���%� ;��A�:魽�   �   �i�/b��gq�y��&�A�h�f��^������P����6��K/��z쎿�+��Td��?�0���>�奄�f�W}�������G��K&��/q�_�ؽ��<������徚�"�-�Z��������� 
ȿ��������A��@��� �`B����߿$ƿ����\q��]�X�D�!�½侇���'Z<�:�ؽ&�s��m*��M������.��   �   j������%���U�7���Ta��Y��|���ʿcLͿbfɿ�Ѿ�����˙��S��X�S��$�2���ǧ�9Z�
����.�B��cC�w��|W��N\��e�����[�%��U�����Z^������~ʿ�HͿcɿ}ξ��|��1ə��Q���S�M$�(��ŧ�L5Z������H�B��iC��|���[�`U\��   �   �����"�Y�Z�B���䚪�Cȿ��῝���vC��B�}� ��E����߿�&ƿ����3s��E�X�v�!���侞����\<���ؽ"�s�&i*��M�]���W)���i�D]�� k����A�B�f��[���ݏ�>����3��[,���鎿,)���d�4�?�3��B:뾞멾�f�z�������G��M&�7q��ؽۺ<����   �   �	��EO�����h���ӿl�����3+��( �׷"�z��-��~
�"v���$ҿ�C��,����N�_���bǾ�S{�t��Û�|�%��3�yA��୽�����a��ɠ��i־x7��Y"��\:�M!M���X��\�J+X���K�Q�8��g ��U��Ӿ^
F]�y���ʧ��7�ع󼘘��������z�@PǾ�   �   i�5�dO|�>1���GѿR[������'�.^7�m�A�ME�OA�SH6��^&��� ����qп�ե��;|�E6�U���'Ϟ�S�:�`4Ľ	2��ݝ�x<�� ���z��,���fF����D����E׾����G
����Ʉ��9�}?	������EԾ����'��aA���������Nw�!��xԈ��'(��m��E\8����������   �   �yV�̂������>�R���,���C���W�L*e�S�i�]�d���V���B��<+��,�� �F���꓿�wW�-U��T���Lc�==�pJ��?�@F;��T�t�ȼFp��ҽ���ғS��w��'8���㮾b���v���ٹ��V��q'�������N�b�U'ɽ�_���� D�8���;�����=�)��]�_�Ao��dS��   �   }	s��$��&�ؿ��o$��*B���^��}w�O��~����׃�0�v�*=^��A�Ҋ$����hhٿ����t�	�)���ܾN)��z�Dg��������<��<��S<����x������ŵܽ����v3�T�L��]�m0b���[��J�8.0���ՄԽhn��v������'�<��<ȏ�<0g��$nX�w��݁���پ�(��   �   ��������=������2���T�&�u��V��L2��w���U���.��|�u���T�΍3�\��Fc�@���Ҏ:����#��g������`û@��<d� =d[=$��<	�;H'���9-��C����}�۽���Ĉ���^��׽����������xR��04<���<��*=�</=��< ����q��A��J���u��z8��   �   �Ë�ҽ��f���b��p<���`�q�������Jq���F���j��C���b���U�a�&�=������������K���_E��j������(�Wi������� = �H=��W=E==n�=H�p< ަ���ȼ�#+�.Hb��`��{���ey���[�J7!���� ��蜔<$=��K=�f=cW=�=��̺������"�����9�����B��   �   �2�������d��F�� �?�7e��i���ו��������������溅��;f��A�e:�����X�¿*ԏ�SI�������+��ō��s����=�U=�ak=R�W=�_'=v�<�0�;�\.�� ׼js��<��F���8� ��0�ü �����%<h�<T�5=�f=��y=�od=��=@���ل�z�&�R圾���ȇF��   �   Ë�5ѽ��e���a��o<���`�����ۑ��ap���E��j��l����߂�0�a�D�=�������3���9K���^E�j�����\(��g������ =��H=p�W=tE==��= �p<�ݦ���ȼ�#+�&Hb��`��~���iy��[�P7!���� ����<T=4�K=��f=�cW=
=@y̺;�����"�̥��������B��   �   �������O�꿸�4�2���T���u�U���0���������-���u���T�.�3���Da쿩���텿�:�e��j�� �������`ûP��<
� =r\=� �<��;�&���9-��C�� ����۽���҈���^��׽���������@xR��14<ȸ�<p�*=l>/=���<`���q�k?��H��(s�+y8��   �   0s��"��u�ؿ^��X}$�(B���^� zw�-��H����Ճ�N�v��9^�Z�A���$�3���eٿ���k�t���)��ܾ�&��V�g��s����<P�<��S<Ё��Ц�m�����ܽ����v3�R�L��]�r0b���[���J�@.0���҄ԽUn�������,*�<��<��<�>��8fX�l�qہ�=�پO(��   �   �uV�5�������:���� ,�Y�C���W��%e���i�ʁd���V�
�B��9+�'*����9C��0蓿�sW�6R�tP��DGc��5～J�?� �;��T� �ȼ$p�Xҽ�����S�{w��%8���㮾g���v���ٹ��V��z'�������N�W�$'ɽJ�_� �� ��8���;���,�=�����_�.k��{P��   �   �5��I|��-��TCѿV�����'�Z7� �A��	E��A�AD6�1[&�������Wmп9ҥ� 6|�A6�����ʞ�D�:�M,Ľh�1��ϝ�h3����z��ڸ��fF�����9����E׾����G
����̈́� :��?	������EԾ����'�� aA�H�������t����Hǈ��(��e��SV8�S��������   �   >��?O�	����c����ӿA������X'��$ ���"�c��0)�{
� p��Vҿ?��{�2�N����D\Ǿ�J{�\�������%��,�ntA�߭�A���a�hɠ�}i־s7��Y"��\:�L!M���X��\�O+X���K�V�8��g ��U��ӾQ�E]���kɧ��}7�d��0��������yz��IǾ�   �   ���f�"�D�Z�襋�����Wȿ���r����?�	?��� ��>��]�߿� ƿ�����n��2�X���!���供���AT<��ؽ��s��^*�(�M�.����(�@�i�]��k����A�=�f��[���ݏ�?����3��],���鎿.)���d�6�?�2��9:뾊멾�f��y����B�G��C&��'q���ؽ��<�Ȓ���   �   �b������%���U�y����[��I
�����*ʿxEͿ�_ɿ˾��y��Dƙ�LO��r�S��$�B�����].Z�y	�%��yB�FZC�t���V�YN\�ae�����P�%�	�U�����Z^������ʿ�HͿcɿ�ξ��|��4ə��Q���S�K$����ħ��4Z������&B��[C�`r��`T��J\��   �   f�i��Y��cf����A��f�gY��
ۏ�R����0��R)���掿d&���d���?�c��4뾧橾@f�)t������G�>?&�x'q���ؽ�<�Д����徍�"�$�Z����������	ȿ��������A��@��� �eB����߿ $ƿ����]q��[�X�A�!����R���lY<���ؽ6�s��a*�&�M������%��   �   N����a��Š��d־f4��U"��X:��M���X�	�\�;&X���K���8�hc �R��ӾRꝾ>]�,�������q7�|�󼴊�P���,���{z��KǾ���AO�x���de����ӿ����+��')��& ���"�}��7+��|
�ns��`"ҿ�A������ʏN����_`ǾP{�&�������%��+�RoA�ڭ��   �   �s��t���`F��w���#@׾f���D
���Ҁ�6��;	�����L?Ծe����"��LYA�+����ꓽ*g��������(�f��pW8�y���������5��K|��.��Eѿ8X�����'��[7�"�A�	E�.A�pF6�/]&�������pп|ԥ��9|� D6�>����͞�P�:�C1ĽX2�4ѝ��,���{��   �   ,�ȼ,�o��ҽ�����S�Os��[3���ޮ�����:p��Թ�"Q��4"�����K�N�`��ɽ�_�� ��8`�;�t���=��轲�_�l��>Q��vV��������;�ј�(,���C���W��'e���i�/�d���V��B�o;+��+�n��eE���铿gvW�WT��S��dKc��:�>J��?� �;`9T��   �    �S<P;����������ܽ���$p3��L��]�l(b���[�8�J�'0��cyԽ�d���t� ����>�<L-�<���<����cX�F��ہ���پ�(��s�#��9�ؿ��~$�)B�	�^��{w�.��d����փ�z�v��;^��A��$�]���gٿk���t���)���ܾ�(���
��g�p�����<|�<�   �   �_=�
�<`F�;����--��<������۽{��~��U��׽���{������8FR�(\4< ��<\�*=�C/=x��<�u�\�q��>��H��s�:y8�����L����������2�H�T���u��U��e1����������-����u�:�T�Y�3����b������:����'��p������xû��<R� =�   �   �W= G==j�=��p<������ȼ�+�@b�~\��ܢ���t���[�p.!�@�������<=�K=��f=�gW=h= ̺������"�7���?���6�B���ѽ��e���a��o<���`�訂�����p��7F���j������5���(�a��=��������3���L��`E�k�%���O(�Uj������N =l�H=�   �   I�=>�r=2�F=Hg=\��< ~;��D�D����z��� �4���������;���<ľ =�H]=
ф=�=�#�=l�@= �M<�7�(%������M���.��'|�*��a�߿�?��`*�Q�I�%|h�����������.Ŋ�̳��=i���J���+�h��
c⿾/������1��羠����P���; \)=*�p=�   �   "�r=z�Z=�4(=��<�k�;�,��Lռ4���Y:�0C��5����8�� ]λ �A<���<�>=�q=B�=XR|=Bm:=��J<�"2���������ݾ�t+�A�w�u<��hܿ�
�Ə'��&F�*d��}�Gʇ����kć���}�!id���F�ݔ(��$�Ƙ޿|0��{�:0.��X�ꆾ����J�Ы�;RD#=�-e=�   �   �<=:i=���<�!_��bڼ>J�*��f1���½�ǽ?���Ĩ�o����7�h��� �;|0�<�i(=�S=��W=fu&=x�><�"�����x�u�L�о�"�!�j�Q��ѿ��t���;�efW���n���~��?��(�~�ҟn��SW�	9<�� ��K�(�ӿz����m�En$���Ծ�k|��v�z9����;v%=�A=�   �    V�<
�;�-���X�3u���񽶣�Je,���:�#�>���8��K)��`���~A��ް@�\C���%<T�<,l=҉=�#<�F���ٽ��[�lż��s�'�V�ד�ӄ����������,��D���X�'jf�[k�)�e��%X���C�'8,���3a��j¿֔���X��9�L�ʢa�^t�t� ���;L4�<��=�   �   �_-�f�)�����z����2�cb�i�����݀������g����+��<���Az\��U,��p��"����U�@���h�_<�7�<@h�;p��w۶���;��i��d� ��;=�F�� V��c�ؿG9�����-� �>��I��tM�Y4I�7�=��-�������6�ؿ{����p���S>�g�M���yT@������X� ��:`<0y<�   �   �i�Q�ս��&��j��Θ��[��zھ� 򾷢 �v����������־ɷ�9!���wc��H ��ʽ�T��^��@щ�@���<�ļ �������h�׾P �x_�����s����b��ѱ�d[#��#,���.�?�+��Q"��������p��6������d_�Cd �6�ؾzz�����#�������������缼�   �   @��e?�&���8������G���K$��"5�޵?��C�v�>�&�3�}G"�D��m�������wj9��z���x��W���c�0K��p�_�F$��bT����#����6�j`t�\~��]h��$�ݿ�$��\1�j5�8l����8�>�����ۿ����KL���r��'6�p_�塬�pgU�<W�g� Gɼ0Ɖ������̄��   �   �&F��ٔ�vо���:'+�KL�(&i����b솿%��\���}�~�f�ZI���(�Ω��J̾lޑ��A�;�齐�{� D �lż6�&��ܩ��@�Uׂ��+Ⱦ"��JA��x�����ʲ�3"ʿA:ܿŇ翊����ڿF#ȿ�Ұ�|e��~u�t?�w��K�ƾ���v���e�� *�H�мTb��P��.���   �   �����Ծ���z"=�k�i�bP�����A���f���ms��m߳��<��h������k�f���:����Ҿ(���87�sԽ<8_�����*��bc�G�׽��9����g�Ծj��g=���i��M��
��'���:���Ip��hܳ�:���e��������f���:����Ҿ���457�kԽ�4_�����\5��~c�7�׽��9��   �   :0Ⱦ%�DNA�Xx�&���Ͳ�l%ʿ�=ܿ?����7����ڿ&ȿ�԰��g��a�u��v?�p���ƾ������h��*�<�мZ��I�����" F�CՔ��оr��$#+��L�!i�!���醿["��wY��*�}��f�0VI�P�(���lF̾Mۑ���A�i���{�B ��żҏ&��⩽9E��ڂ��   �   �����6�odt�À��"k��@�ݿ�'��*3�F7�n�����9����j�ۿ�����M��(�r��)6��`�ѣ���iU��Y�,�g�8Aɼ���,v���Ą��v�p^?�����������{��^G$�H5�D�?�'C�	�>��3��C"����g�u������Ze9��s潚�x��M༘�c��Q��B�_��*�hT������   �   � �R{_�����������������D]#��%,���.��+��S"��������r�f8��>����f_��e ���ؾ�{���������8�� ޷�`Ш�ϼ��i�I�ս��&�w�j�nɘ��U���ھ��� �� �����`����־
ķ�����pc�SC ���ɽ��S��P���g���	����ļZ$������!��5�׾�   �   >=����X����ؿ�:���� .��>���I��vM�(6I���=�G-����l����ؿ�����q���T>��,���PU@�5����V� f�:�%`<(�<�,-�ʂ)�����2�mZb�Gd������{��{���K{��,'���ۃ��r\�pO,�wf��/����I�P^���_<<;�<�]�;���߶���;��l��F� ��   �   t�V��ؓ������������,�z�D�S�X��kf�'k���e� 'X���C�	9,����8b�k¿�֔�t�X�K:���+�a�0t但� ��:�;�>�<��=�h�<j�;���W��j������>^,�F�:���>���8�rE)��Z�����8��¢@�t-��X�%<@!�<6o=`�=x<L��ٽE�[��Ǽ��u��   �    k���ѿ؈�u��;��gW���n�U�~�H@��g�~�ؠn��TW��9<�� ��K���ӿTz��7�m�\n$���Ծ�k|�v��w9����;�)=�A=��<=Nq=$��<`h^�(HڼJ�2"���(���½�ǽu6������/���X�7�఼�g;�=�<bn(=
�S=�W=�t&=��><��"�������u���о"��   �   ��w�X=��iܿ�
�t�'�Y'F�d��}��ʇ�	���ć�l�}�jid���F��(��$���޿V0���{��/.��W⾍醾$��r�J����;nG#=@1e=�r=�Z=�9(=0��<��; �,�<ռ|���P:���B��5�Z������0/λȨA<��<��>=��q=��=R|=�k:=��J<b'2�X�� ��w�ݾ�u+��   �   �(|������߿@�>a*���I�w|h�'����������Ŋ������i���J�l�+���sb�6/�����H�1�� 羼� ���P�`2�;V^)=�p=�I�=r=��F=�h=Ԓ�<��;P�D�܏��z�� �\4輤�������	�;���<�� =�G]=cЄ=M�=�"�=0�@=��M<�7�x&�� ��/O�­.��   �   ��w��<��#hܿ�
���'�s&F��d���}��ɇ�C���Ç��}�?hd���F�+�(�C$���޿�/���{�/.��V⾾膾���J����;�H#=2e=��r=x�Z=":(=���< ��;��,��;ռx���P:���B��5�h��  ��/λ �A<<��<ڿ>= �q=��=�R|=�l:=��J<�$2�N��U��N�ݾ,u+��   �   ��j�!^�ѿć��s�Z�;��eW���n���~��>����~�^�n��RW��7<�� ��J���ӿ�x�� �m��l$�`�Ծhh|�t�4r9���;�+=NA=��<=r=0��<�b^��Gڼ�J�!"���(���½�ǽ6������3���Z�7��߰� j;L>�<�n(=��S=D�W=�v&=��><r"�������u�J�оp"��   �   z�V��֓�!������,����,�˔D�0�X��hf��k�R�e��#X���C��6,����_�i¿�Ԕ�c�X�8��￾��a�yn��� ��b�;LE�<$�=�k�< r�;�����W��j������8^,�H�:���>���8�xE)��Z�����8����@��,����%<�#�<q=R�=.<�D���ٽ �[��ļ�ns��   �   �:=�� ��U���ؿq8������-���>�7�I��rM�b2I�W�=�9-���6���ؿ����No��?Q>�s��n���8P@�h���M� %�:�5`<��<�%-���)�%����2�[Zb�Ad������{��~���Q{��2'���ۃ��r\�rO,�df������I��S����_<LB�<���;��mٶ���;��h���� ��   �   � �/v_��������2��6��k���Y#��!,���.�O�+�P"�։���"n�f4�������a_��a �<�ؾ�w��P��3����p�𩷻𭨻pɼ�� i���ս��&�M�j�^ɘ��U���ھ��� �� �����f����־ķ�����pc�:C �g�ɽ�S��K�� �G���ļ=��C�������׾�   �   �����6��]t��|��Pf����ݿ�!���/��3�ej�"��=6������ۿձ���I��z�r��$6��\�����aU��N�:�g�P-ɼ����pm��_Ä��u�^?�����������u��ZG$�G5�D�?�*C��>��3��C"����g�r������-e9��r�<�x� F���c��>���_�$ �`T�����   �   �(Ⱦ ��GA�zx�z��)Ȳ�qʿ17ܿ{���|�濕�ڿ ȿ�ϰ��b���yu�Fp?�s����ƾC�����]����)�}м�S��G��/��F�Ք��оg��#+��L�
!i����醿\"��yY��.�}��f�4VI�R�(���cF̾7ۑ�0�A�J��X�{� < �`�ļ��&��ة��=�EՂ��   �   �	����Ծ���N=���i�qK��x��S���5���(m��Eٳ�7���b��ښ���f���:�V���Ҿ|���.7��Խ:%_�����T����b�e�׽>�9�m��G�Ծ]��_=���i��M��
��&���:���Jp��kܳ�:���e��������f���:����Ҿu���47��Խ�/_�D�������b��׽��9��   �   \F�	Ҕ��о����+��L��i�'���憿����V��Ԥ}���f��QI�H�(�����@̾�֑��{A����ܲ{��3 ���ļ��&�Yک��?�ׂ��+Ⱦ"�vJA��x�����ʲ�1"ʿ@:ܿƇ翎����ڿH#ȿ�Ұ�e��~u�t?�q��0�ƾ�������c���*� �м R��D������   �   �n�Y?����(������3���C$�$5�ج?��C�z�>���3��?"�J�a�񊶾*��$^9�Ih潒�x� 0༐�c� 8���_�2"�HbT�܊������6�b`t�Y~��Xh�� �ݿ�$��\1�k5�:l����8�C�����ۿ����LL����r��'6�h_������fU�YU�l�g��4ɼ����dd��羄��   �   ��h�ĽսR�&�qj�Ř��P��ھ򾨛 �M��z�����ﾃ�־D������Vhc�N< �x�ɽZ�S�<3�� ؇������ļx��:�����@�׾C ��w_�����o����`��б�d[#��#,���.�@�+��Q"��������p��6������d_�@d ��ؾDz����������y�@���P�������   �   �-��u)�G楽����2��Rb��_�����|v��=���v��#"��>׃�Lj\�H,��Y�������8�0�`<�O�<p��;��鼉ٶ�Q�;��i��V� ��;=�D��V��a�ؿF9�����-� �>��I��tM�Z4I�;�=��-�������7�ؿ}����p���S>�^�*����S@�����R���:�;`<H�<�   �   @v�<���;������W��a�����3���W,�S�:���>���8��>)�HT��潀.���@�l��P	&<(6�<*x=��=H<<�B�T�ٽf�[�Lż��s�"�V�ד�҄����������,��D���X�'jf�^k�*�e��%X���C�)8,���4a��j¿֔���X��9�5�k�a�s�\� ��O�;�E�<��=�   �   ~�<=�v=��<��]��2ڼn�I����� ��Y	½1�ǽ�-��鳨������7��Ű�`;xQ�<�v(=D�S=f�W={&=��><�|"�����8�u�;�о~"��j�O��ѿ��
t���;�efW���n���~��?��)�~�ҟn��SW�	9<�� ��K�(�ӿz����m�Dn$���Ծ�k|�v�jw9����;2+=j	A=�   �   2�r=��Z=�<(=|��<���;��,� /ռ6��
I:�(�B�H5�����︼p�ͻ��A<��< �>=��q=��=.V|=p:=��J<�!2�l�������ݾ�t+�>�w�t<�� hܿ�
�Ǐ'��&F�+d��}�Gʇ����kć���}�"id���F�ߔ(��$�Ș޿}0��{�90.��X�ꆾЀ�>�J�p��;&G#=�1e=�   �   pӎ=�=��g=��3=���<X �<p��;�	���e2��SH�p��@���h�<P��<p�=>�T=Y��=�w�=Σ�=��=hWr=�&�<�O��^˽�QX��K��Ϊ��tW�<���¿ea�]�	"-�\�E�CZ�Vh��Um�S\h�tnZ�J�E�:�-��Y������(Ŀ�2��l�Z�ۤ�������a���ܽ����Lp�<�M=';�=�   �   ��=��x=�L=��=��<��;��t8��@V˼|ؼ 뼼ؖx���]� �8<(v�<��3=fp=ю=ҵ�=`��=�l=L��<DҪ��_ŽZS��r�����S�޺���ݾ�=��w ��>*��B��+V���c�o�h���c�:V��[B��*�l��v�N���m�����V�x���r���y\���ֽ��\3�<�fH=V�=�   �   `�^=��8=�B�<�L4<�%�x��*s=�vvt�*��ՙ��U����e�p�(�L0��@�����<
=��\=�y�=��=xZ=Lj�<�F������E��I�����FtH�al��_���,B�P(
�;�!�$8�4�J��V��H[�k�V��YJ�8��'"���
�P��o'��g���2&K��1�#����EM��Ž��м�ӟ<��7=�b=�   �   �=b�< �����by��q��ϻ��o�{���
�P��L����ܽ�����yZ��sż`�V;���<h%/=:�L=�:=\ �<xjU��5����.��$����6���}��2���ҿ����8)���(�H;9�8�C���G��C�v�8��(�������+ӿ���f����8�{���&�����5��4������{�<�0=��+=�   �   ��;,2��<i�K�Ž
j�>�6�Nc[�Rx�0�������σ�f�s�@XU��z/��_�Pд��G�g�(DO<<��<�V=���<����Y|�Y����9�׾�� �H`����1������F!��f��@$��6-��(0���,��y#�ޖ�!~���H���ɴ���a���!�Meھ�������ڞ��Xi��P}<d��<<�<�   �   ���򝽽0�P>��{����.8����ʾ�ؾ�	ܾʧ־}kȾ����^�����r� ?5��z�����d�� �C:���<p�v<����V5=�9�hA[������/���>�t4~�G�����Ŀ�濈���y�q���9��W����d� ��]俲Uÿ�à��}��y>����1贾Ni^�����[N�(B� <�#<p1���   �   ɮ���U���b����̓ƾ���������"���%�A"�N%�� 	�#
�]���m���XZ�n��s��r�� ���@��;@�P��;�[?���I)��I���پ�/�t�P����¡��>��ٿyf�,����^������X���׿91���������4O�Eh�8پ^`��{*�BH���C�`�׻ X�8X�I���,��   �   ��kt�q����������-��1G�~�Z��Mg��)k��8f���X��D�+�w]�W���V���_m�^*���� 3��h:��c��������i��:�\|T��o���9�O$�KCT��Â�oI��lܮ�^ʾ�E�ȿ2�˿��ǿ�M���
���t���&��^�Q�+q"����ؤ���R�N����j� `�� (黸og��(��[���   �   VEo����������� ���G��Tm��"��H铿7᛿�^��o2��2���B����j�q�D�'�����{���j����
��
�`�5�x�<��2�������p>o����)���� ���G��Om�` ���擿kޛ��[���/����������j��D�Z$�����x����j�������"����5��<��;�u������   �   �s���>�_R$�FGT��ł�	L��D߮�[;�S�ȿ6�˿��ǿuP�����v���(��J�Q�ts"����Lۤ�<�R�B��j�`���黈Rg���(�9S��S��zct��������T���-��-G���Z��Hg�%k��3f�'�X��D��+��Z����AS��{Zm��&����T-�Pa:��r��0��ޱi��B��T��   �   :�پ�2���P�5���3�������ٿ�i�`����a��������U
׿a3�����6�����O�j��پ
b��}*�HJ��*D��r׻ ��8��I���,�j���`O�!�b����ƾ���2������"���%�d"��!�^��}쾠���Hi���RZ�����l��J��`������; �P��B�'E���M)��L���   �   -2���>�8~�f���p�Ŀ> ��� {���l;�pY������ ��_�lWÿVŠ��}�8{>� ���鴾2k^�k��\N�x:�x<�#<�ھ�`��靽�*���=�5�{�󧛾�2��z�ʾ� ؾNܾġ־�eȾ��������Q�r�"95�Vq������u� 7E:T��<x�v<�ݔ��<=�i�F[�洳��   �   $� ��J`�ȉ��5»���㿔"�Gh�LB$�98-��*0�)�,�E{#�����Q�}�������7 a���!��fھ_���:������i��_}<0��<� �< j�; ���i�4�Ž{c���6�[[�l�w�����🇾�ʃ�!�s��PU�t/�
Z�jǴ�G���f�(aO<���<HX=T��<����a|�1\�
��~�׾�   �   ��6�H�}�+4����ҿ����a*���(��<9���C���G�V�C���8�ځ(����
��ӿy��W��O�8�A���������5��4��D���0��<�5=>�+=H�=0w�<в��P��
y�"g��S���i�'����6�������ܽ�����jZ�[ż�5W;��<8*/=��L=6:=��<p|U��9����.�I𛾵'���   �   �uH�pm�������C�$)
�,�!�.8�R�J�;�V��I[�b�V��ZJ��8�C("��
�ȕ��'������f&K��1�!����EM��Ž8�м$ٟ<j�7=��b=�^=��8=�S�<�u4<����켚d=�gt�>�������M����e���(���@z�� /�<�$=\=J{�=y�=�wZ=�e�<�O��#��=E��K������   �   ^�S������޾�F���(?*�pB��,V�f�c��h�J�c�s:V��[B� �*�x��v�9���L���6�V�/��r���x\�k�ֽ��Ｔ8�<�iH=��=��= �x=֦L=�=0!�<��;���)���F˼L�׼�ܼ�h|x�@Z]� �8<d~�<ڽ3=�p=�ю= ��=?��=��l=\��<Lڪ��bŽH\S�t��"���   �   �uW��<���¿�a�b]�Q"-���E�NCZ�3Vh��Um�9\h�DnZ��E���-��Y�#���G(ĿU2����Z�0�����R�a�@�ܽ����u�<�M=<�=2Ԏ=��=�g=�3=@��<<"�< ��;����c2��RH��������0�<܍�<��=T�T=ʕ�=+w�=��=�=hUr=�!�<�V���˽pSX��L��{���   �   c�S�����ݾ�L��r �m>*��B��+V�C�c�ؚh�#�c�e9V�
[B�\�*�����t�a�������0�V�o��	q��Ww\���ֽd��0<�<�jH=K�=�=��x=&�L=F�=�!�<@�;0���(���F˼@�׼�ܼ�x|x��Z]�0�8<|~�<�3=�p=�ю=S��=���=��l=���<�ժ��`Ž�ZS�s��j���   �   tH�7l������A�(
���!��8�o�J�&�V��G[�H�V��XJ�8��&"���
�ғ�&&��Tߋ�u$K�{0�!����BM�$Žt�м�ߟ<��7=&�b=2�^=z�8=U�<`w4<0��`��jd=��ft�3�������M����e���(����w��X/�<%=<�\=�{�=�=�yZ=�k�<�F������E��I������   �   �6���}�2���ҿ�����(���(�2:9���C�.�G���C��8��(�������Xӿ?��е���8�S����~���5��/���r��T��<�8=h�+=��=\y�<P�������y��f��.���i�!����8�������ܽ�����jZ��Zż�:W;H��<D+/=��L=�:= %�<�bU��4��V�.��훾�#���   �   � ��F`�0���
���8��` ��e�z?$�15-�d'0��,�px#�m���|�z��?������a�\�!��aھ���¿����P�h��u}<���<�< x�;l��
i�؞ŽVc���6��Z[�b�w�����򟇾�ʃ�'�s��PU�t/�Z�SǴ��G���f��eO<���<x[=H��<0���U|��W������׾�   �   �.��>�R2~�芡�L�Ŀx�U��+x����98�NV����� �"[�@Sÿ����R}}��v>�����䴾(d^��~�tON����,<P�#<�ľ�f��Y蝽d*���=��{�㧛�}2��s�ʾ� ؾMܾǡ־�eȾ��������P�r�95�"q��p�� s� �E:D��<0�v<���T0=��3?[������   �   g�پ".�&�P�����󟣿���ٿ�c�+����[��w���<���׿�.����������{O�le��پ]��
v*��@���6�@*׻ <�8 �I��,�s���O���b������ƾ���,������"���%�f"��!�a���쾠���Di���RZ����l����@��� Ӊ;�<P��5��;���F)��G���   �   6m��6��L$�`@T�����NG���ٮ��Ǿ�c�ȿ2�˿��ǿ�J�����r���$��h�Q��m"�ҫ��Ԥ�ǷR�����j�|F�����;g���(��Q�����(ct�s������K�|�-�-G���Z��Hg�%k��3f�+�X� �D��+��Z����8S��QZm�:&����*�L:� 1���좼��i��5�xT��   �   �9o�Κ������K� �3�G��Km���䓿�ۛ� Y�� -�����w����j���D�� ����:t��t�j�3��������P�5�p�<��-�����z��>o�᝱������ ���G��Om�] ���擿kޛ��[���/����������j�"�D�Z$�����x��b�j�@����F��ع5���<�"+��~������   �   "���]t�ڋ����k��-��)G�_�Z�Dg�8 k�/f�x�X���D�� +�W����`N���Rm�p �%���p-:�����뢼Ԣi�]9��{T��o��q9�
O$�BCT��Â�kI��kܮ�\ʾ�F�ȿ3�˿��ǿ�M���
���t���&��^�Q�)q"����ؤ���R�	����j� S����軐5g�V�(�M���   �   \����J���b�-��<�ƾB����c����"���%�j"������������}d���JZ�����b��F���n��0�;�P�6�d=���H)�mI��ɞپ�/�j�P��������=��ٿzf�,����^������[���׿<1���������5O�Bh�'پ:`���z*��F��>��D׻ ��8��I�R�,��   �    ���᝽�%���=��~{�~���n-����ʾ��׾�۾��־�_Ⱦ����􍗾��r��15�e�������U輀�H:�̂<��v<�����0=����@[�r����/���>�k4~�C�����Ŀ�濇���y�p���9��W����e� ��]俴Uÿ�à���}��y>���贾�h^�(��xWN�`'��)<0�#<@����   �   `��;P���^�h��Ž�]�,�6��S[�%�w�,섾c���ƃ�\�s��HU��l/��S�]�����F��f��O<���<�a=��<���V|�xX�����׾� ��G`����/������F!��f��@$��6-��(0���,��y#�ޖ�"~���J���ʴ���a���!�>eھ|�����-�����h�Po}<��<�<�   �   N�=��<�`�������x�^�����d���C���|����i�ܽ�맽�XZ��;ż�	X;8�<�3/=��L=�:=�+�<[U��4����.��훾�$����6���}��2���ҿ����8)���(�I;9�8�C���G��C�x�8��(�������,ӿ���g����8�q������+�5��3��D|����<�8=��+=�   �   ��^=r�8=0`�<ؔ4<�������W=�Yt����8����E����e�|�(� ��@��XC�<�-=@�\=�~�=`�=(}Z=�q�<�A�����RE��I�����@tH�`l��_���,B�O(
�;�!�$8�4�J��V��H[�l�V��YJ�8��'"���
�Q��o'��h���2&K��1�����EM��Ž��м�ڟ<��7=��b=�   �   ?�=��x=>�L=H�=T)�<�>�;�l�T���8˼��׼�ͼ� _x�@�\�x�8<`��<4�3=�p=�ӎ=��=��=x�l=ܜ�<�Ϫ�6_Ž�YS��r�����S�ܺ���ݾ�=��w ��>*��B��+V���c�p�h���c�:V��[B��*�l��v�N���n�����V�w���r���y\���ֽ����6�<:iH=�=�   �   ��=@]�=Fa�=X�W=ʝ(=�N�<P�</Q<H�<��<��4<�9�<$��<�`!='W=�j�=�O�=B̯=3��=�h�=_ȓ=�#;=@�;Di��!g"������0�lv�lO��l�̿j�����Jr$�W4�4�>� �B���>��t4���$����|o��Tο
��mxy��4�
�������'.��嚽�-��`=�l=�ʐ=�   �   R��=�z�=Z�k=�;=�+=\T�< �<�g�:@V[�5���]��)�;hʊ<DW�<�]5=n5p=f��=^��=
�=ծ�=�0�=�G:=@$L;|Q{�PE������?�4�-���q������Nɿ�����A�!�8;1��;��?�5};�D1�n�!�6�G����ʿO=����t�߯0��	�}'��c�)�O������N�=Dfh=���=�   �   �G{=��Z=8�%=x��<(<h��x�� (	�0�#�j)�bw�����|��Vs:葛<��=d_]=<�=p�=3�=4�=F7=Pb�;#`��V��7��(�ܾ�0$��Ce�����1���/}�������T(��1��5���1��)(�?��b'��;�e���B���c�g��&�G��&=��2��@$��@R��=�@[=��~=�   �   �`6=>�<8M3<��A��r�F q�h.���M½��ս��ڽ5�н&���t����K� �̼ LX9,��<v 3=��l=��=�~u=t�/=К<��6�����Z{s�RbǾ d���Q��J��j}��jֿD�����^��.#�*&�p�"��W��[��{��Nwֿ�밿����dXS�w?�RJ˾״{�`����]���{�4� =;C=F0Q=�   �   8e�<`�]���Y���ν��	�>(�'�?�-�N���R���K���:��� ��k �����_�4z��8�<~�=�<=.�I=
� =P�X<6���ѽ�N��l�������8���v�휿�1��<�߿����p�	�$�S��!��G	�L���b�޿꙾�������v�RM9�Ԟ�d���U���߽V�$�p��;T�<h=8�=�   �   �i���J�����A�E�C�o�u������B�����A������n�����Xl��9�d��5������ Wo��"�<|==dB=2�<�硼R��+,&�����pھ ���R��t��Ć���2���[ڿ���[��BT�����b��f�ؿ$˿�u��nȅ��iQ�����۾$m����)�����Ѽ�<���<<b�<�8<�   �   .@o�R��A�.���t�Hܞ��4¾�ι��0��}���������2ݾ����d����i��R$�>�̽raJ��66�(^<P�<<q�<�8��Y�����e�]��4��,R��M�+�|d]�h>��ţ������גƿ��п�:Կ�-п:ſQa�����[冿,^[��A*�A���)�����]�/���r�c���>��JB<�p�<0R�;�����   �   d�轑W=�FӉ�Hƹ�K����yr#��&4�\�>���A�r�=�M2�a� �oF�澲d���섾z�4�&�ٽd�R�X[N��7<8>p< ��:h���>���_!��_���B¾���U|.�2ZX��@��Lޑ�%������+���`���J��~R���O}��pU�s,���ϐ������5��U��L��� ��9 �B<@X�;|���l��   �   �{8�����kƾ���`�#�L�C��_� �u�������������rs��]���@�.!��b �
¾Ln���2�Jd̽_6���	�@V<0n<�)'��B��	ս�u8����gƾ�����#�E�C���_�T�u�����K������mns��]���@�\!��` � ¾�k��U�2�9_̽�X6���	�xS<�^<�G'���B��ս�   �   �b���F¾����.�(^X�+C������������������b��*M���T��]S}��sU��,������������7��X����� ��9��B<���;����|l����(Q=�0ω�?���N�뾊��n#��"4�8�>���A�z�=�_I2�� ��C�:��`���鄾�4���ٽ��R�hGN�8><8p<@��:��������d!��   �   �8���V��I�+�h]��@�����~����ƿ{�п�=Կ&0пd<ſqc������憿�`[��C*�7���E���t�]������c��>�xSB<�z�<@��;����d0o��}ཪ�.���t�tמ��.¾��,
��̱���������#-ݾ4���`��1�i��M$��z̽�VJ��6�0^<��<tl�<�O�t$Y�@�����]��   �   Qtھ����R��v��݈��5��^ڿ���^���V���������q�ؿ�̿��v���Ʌ�lkQ����۾tn��r�)� ���x�Ѽ@�<4��<�n�<@48<�h���J�s����:�ҿC��u�A����=�����k<��㌫�Mi�������
l�k 9�U��H���ư���n��-�<@=*B=�+�<����>W��0&�`���   �   t���8�n�v��|3��p�߿������	�J%����O��&H	�$�����޿3�������L�v�{N9����t��4U���߽��$�P�;��<m=R�=Hx�<@]����O���ν��	�7(���?�r�N��R�:�K�ȣ:�9� �f �����x_�\b����<��=D	<=��I=� =��X<�<���ѽ��N��o���   �   �e��Q� L���~���kֿ4��� ��z��9/#�?&�r�"��X�C\��|��Ixֿ�찿!���3YS�@��J˾��{����p�]��M{��� =�>C=�5Q=�g6=�O�<Xy3<�]A�c��q��$��4C½@�ս��ڽ�нp���k��V�K�<�̼ �b9�	�<�3=��l=��=�~u=�/=h�<j7����s��dǾ�   �   2$��Ee����r����~连������U(���1�\5���1�O*(�����'�><�μ��������g�9�&�j��%=�����#�� D���=�C[=p�~=�L{=��Z=��%=���<h+< ������	���#��\)��j���鼈�{� �u:�<��=fd]=�=�=��=3�=�=h7=D�;
)`�'Y��9��Z�ܾ�   �   M�-�R�q����oOɿ�����ɷ!��;1���;�/?��};�ED1���!�6�0G����ʿ==����t���0�E	�'����)�����p����=�hh=���=ׄ�=�|�=~�k=��;=H1=`�<`�<�:�:`�Z�P����[��V�;\Ԋ<�_�<da5=,8p=`��=���=I�=���=0�=�E:=��K;�V{�(G�Ά���A��   �   g�0�=v��O���̿������{r$�,W4�H�>��B���>�lt4���$�J��o���Sο����wy�44�����$���2&.��㚽�-�Vc=��l=_ː==�=�]�=�a�=p�W=Ҟ(=<P�<��<H1Q<�<0�< �4<`9�<$��<L`!=X&W=�j�=jO�=�˯=���=h�=vǓ=$!;=��;?k��xh"�b���?���   �   x�-�:�q�Л���Nɿ���
���!��:1���;�N?��|;�xC1���!��5�$F����ʿ�<��v�t���0��*&��j�)�U���H��2�=�ih=[��='��=�|�=��k=�;=�1=t`�<�<�>�:��Z�� ����[�W�;hԊ<�_�<~a5=D8p=v��=��=}�=���=�0�=�F:= L;�S{��E�����y@��   �   |0$��Ce�����֬���|������T(�Z�1��5�!�1��((�i���&�@:� ���)󘿌�g���&���s;�����l ��!���=�E[=�~=N{=��Z=J�%=��<`-<�}�����	���#��\)�tj���鼈�{� �u:��<&�=�d]=!>�=��=4�=��= 7=�c�;#`��V��7��	�ܾ�   �   }c���Q�)J���|��!iֿ���;�����-#�&�Q�"��V�tZ��y���uֿM갿9���1VS��=��G˾�{�j����]���y�� =�AC=�7Q=Zi6=|R�<�}3<8ZA�vb�q�z$��C½*�ս��ڽ�нm���k��F�K���̼ c9p
�<23=��l=��=H�u=��/=��< �6������zs��aǾ�   �   ш���8���v�윿B0����߿����e�	��"�������E	����,�޿ꗾ�4�����v��J9����	���U��߽(�$��A�;�#�<�p=��=(|�< �\�b�8O����νs�	��6(���?�d�N�ާR�;�K�ɣ:�:� �f ����^x_��a����<��=<=j�I=r� =��X<�2���ѽ��N��k���   �   �nھ����	R��s��P����0���Yڿ���^Y���Q��f��������ؿ�ȿ��r���ƅ�xfQ�+���۾5j��p�)�����LzѼX�<`��<�v�<�?8<��h��J�ȟ���:���C���u�/���v=�����i<��㌫�Oi�������
l�e 9�F���������n��1�<C=�F=X:�<�ޡ�AO��B*&�=���   �   �2��<O��V�+��a]��<��������x�ƿ3�п:8Կ�*п\7ſ�^���
��Dㆿ�Z[��>*�n���m�����]�������c��k>�(tB<���<p��;�z��L.o�"}�X�.���t�Xמ��.¾݆�"
��ɱ���������&-ݾ3���`��$�i��M$�^z̽zUJ��6��'^<�#�<P{�<�#�2Y�����^�]��   �   {]���?¾����y.�$WX�?��7ܑ�Յ��g������t]��PH��P��QK}��lU�,���a�������/�xM�� ��� e�9��B<P��;0����l�����P=�	ω� ���6�뾁��n#��"4�5�>���A�{�=�bI2�� ��C�9��`���鄾��4��ٽؓR��;N�(Q<�Tp<�T�:��������\!��   �   �q8������cƾK���#���C���_��u�I�����&���is���\���@��	!��] ������g��<�2��U̽J6�(V	��<0�<�'���B�OսSu8�����fƾ�����#�=�C���_�R�u�����L������rns��]���@�_!��` �w ¾�k���2�h^̽FV6�Xv	��m<Ѕ<x'�@�B��ս�   �   ���[L=�̉�?���`�뾟�Wk#��4�?�>�j�A�^�=�dE2�R� �'@�H澽[���儾K�4�9�ٽH�R�(N��k<�bp<@g�:�����
��f_!�p_��eB¾���J|.�*ZX��@��Jޑ�#������-���`���J���R���O}��pU�r,���Đ��v����4�xT������ ��9��B< ��;�됼�l��   �   0$o��u�n�.�$�t�eӞ�'*¾g���������(��,���'ݾ���\���i�G$��o̽tEJ��5�xI^<P.�<̀�<H#��Y�������]��4��R��@�+�rd]�d>��£������֒ƿ��п�:Կ�-п:ſTa�����\冿-^[��A*�9������^�]�B���P�c�8�>�hB<��<���;n���   �   @�h���J�����5�t�C�^�u����8��� ��17������Fd������|l� �8�
��ҝ����� �m��D�<�I=RK=�>�<ߡ��P���+&�q��qpھ��}R��t�������2���[ڿ���[��DT�����f��f�ؿ%˿�u��nȅ��iQ�����۾m��~�)�H���@�Ѽ��<���<�z�<pR8<�   �   ���<�t\����G����ν�	��0(���?��~N�5�R���K�d�:�R� ��_ ������e_��B��h <�=~<=��I=�� =ЭX<�2���ѽ��N��l�������8�z�v�휿�1��;�߿����q�	�$�T��#��G	�N���d�޿꙾�������v�OM9�ў�S���U���߽Z�$�� �;� �<�q= �=�   �   m6=�]�<�3<�1A��U�*�p�����9½��սi�ڽQ�н6��Ab����K�g̼ Pp9� �<:3=�l=��=z�u=v�/=�<|�6�/���{s�<bǾ�c���Q��J��j}��jֿD�����_��.#�*&�r�"��W��[��{��Nwֿ�밿����dXS�w?�GJ˾��{�����]� �z� � =�AC=�9Q=�   �   �O{=ީZ=�&=d��<L<�X�Ḽ�	��#��O)�D]��鼠�{� �x:��<Χ= l]=.A�=l�=
6�=t �=�7=`t�;v!`��V��7���ܾ�0$��Ce�����0���/}�������T(��1��5��1��)(�?��c'��;�f���B���c�g��&�A��=�����#���A��ڇ=*E[=��~=�   �   M��=a}�=��k=p�;=�4=�h�<��< �: �Z�χ���Y�`��;|��<(k�<�f5=�<p=���=ۈ�=�=\��=�1�=DI:=@5L;�P{�2E�|����?�1�-���q������Nɿ�����@�!�8;1��;��?�7};�D1�n�!�6�G����ʿP=����t�ޯ0��	�v'��N�)���������=hhh=��=�   �   	��=vc�=��=�o=��K=��)=��=\2�<��<�a�<���<(�=@�;=�\g=�M�=��=d�="��=N��=:�=��=���=40�<�Y�|۽�1\�p˷�P�
���C�����C�� ʿ���Z��%@�pQ���AS��R���F��*˿eQ��k��m�F�a��V��Wlj�����j�<����;�(=�n}=�=�   �   ⃔=6B�=�f}=�X=*0=��	=���<�< R�<<q�<Tת<�>�<��=X�F=9z=L��=�l�=薾=ھ�=�!�=�b�=�G�=4<�<!ۼqԽD	W�� ���G�q@�ql���B��I�ƿ���c�����G���w����j����`����ǿwl��"���=C�}8��F��i�d��F�rg3�`e�;�d)=X�z=f��=�   �   �Є=0�n=��D=��=��<p�"< QZ�P��8�X��>]����@t����&<$U�<\a#=Doc=V�=*��=(��=��=�B�=.}=��<����I���H�~���\� �/$6�ͳs�13���<��W�ݿR�������N�:��6����Ⱥ���޿Hǽ����ִu��i8�������KsT�!�ݽ���4<@+=rkq=F��=�   �   d�R=�G#=��<�>�;��X�t� ��qA�nr�g���k���2��xaU�8i������PQ;�l�<\�5=hz=G|�=t��==��=
�u=�0=��\������0��̗��龚�%��_�����'��l̿�%�Z2�������1��d���ڢ�K$̿Z0���Վ�p/`�`�'����.���;�]���r�l��<:�+=D7`="j=�   �   �=(O<�	:�2�����ʭ��.����	�r!��������`ڽ�[�� �P��i���j�;$�=�<P=T,�=Rm�=z�g=\=�rz�p�}��N�����\ʾd��D��[|��������οj��;���� 7���߿N(Ϳ�N��DJ���|���D���m�̾������$��P#{��D�<��'=r;D=��4=�   �   `��;�%ɼ��t��ʽ���|�6��4Z��u�UL�����G���?�n��^P��q*��Y �������1�x��(��<d�)=��T=�?P=`�=P��;�F,�P��S�m˧�m"���l&�JW��~���d���^�������˿�NϿZj˿ڹ���9��)P�������U�\�%���~���+V�֢�t�G��l ����<�u=\9=\�<�   �   P���Q~��1����6��_q�-��Ci��h¾�fξ�
Ҿ��̾��������=����c��C(�@�޽�q�tᎼpg<<�=b�,=�=�C~<�ǵ�󇡽� ���8�þ����/�Z��@�����Z⠿����V��s���\۟�ȑ������W���-��������7��� �T>��0�Ӽ�"<���<=���<@��:�   �   L�����.O�(f���۶��޾9j �p ����~����:�n����LؾO������,�B�1R���ㄽP\��@qE<D�<�8=��< �|���B�d�W�B�#�����о�f	��+���L�D�i�FW���u��浉��膿��~��fg��J�)�����̾����P>���ٽ�{=�����Lb�< 1�<P��<���;�%��   �   ���Z�S��i��j̾ � �g��o�1���C�kO��R�
N� �A��X/���l���b~ƾrS����J�*���`�v���u�(kn<�D�<��<8�@<𰟼 Ƈ����(}S��e���	̾� �����1���C�tO��R�:N���A��U/��������zƾ�P��T�J��{����v��u��sn<D�<�|�<�@<�ß��̇��   �   ��B�����=�о�i	�L�+�I�L�N�i�hY���w������ꆿ��~�Hjg��J��)�����̾{���.T>�Kڽr�=��Ў��a�<�5�< ��<�9�;��=D������O�b���ֶ��޾#g �%��2��ϑ��7������GؾV���w��*�B��J��(ބ��M��0�E<D�<V7=��<�p}���B�1��   �   
���þr����/�Z��B������䠿c����X������Zݟ��ɑ����A�W�.�D��~���S9��a� �8A��,�Ӽh"< ��<�=���<@��:�����u�������~6�Xq��(��Gd��¾haξ[Ҿ��̾ï�������9��O�c��>(���޽Rsq��ώ�0g<v�=�,=�=1~<�׵�����[� ��   �   {Χ�j&��)o&�NW�O����f���`������K�˿QϿrl˿ǻ���;���Q��P�����U���%�Q��"����-V����8�G��x ���<�x=n>=(�<��;0ɼ>�t��ʽ�����6�*-Z�̢u�H����&�����n��WP��k*��T �3���̶1����<��<��)=��T=�?P=��=P��;lO,���佁S��   �   �_ʾf�^�D��^|�b������οx��P��	��
9쿠��)Ϳ�O��WK��A|�	�D���̾�	�����%��X%{��F�<h�'=d?D=4�4=Z=@:O<��9�������~������	�"�0��Д�����Uڽ�R����P��P����;�=6BP=�-�=�m�=��g=
Y=��z��}� R�*���   �   ��b�%�)
_�T����(���m̿`'� 4��p�������ϥ����O%̿,1���֎�b0`��'�}�쾠.��p;�����r༜��<D�+=X:`=vj= S=RO#=��< ��;��X��� ��aA�rnr��}������B*���QU��Z�Ln�� �Q;T~�<:�5=6mz=~�=s��=r��=Ʒu=t-= �\������0��Η��   �   �� ��%6���s�=4��>����ݿ�������RO�����6�v�������޿�ǽ����I�u� j8���ɀ��LsT�֒ݽ���4<+=�mq=޵�=�҄=4�n=��D=��=�$�<�!#< �W�Є���X�`]��m��5����&<�d�<
h#=�tc=r�=���=%��=��=�B�=p,}=ؾ�<�Ư�HM��\H�J����   �   �H�+r@�m���C���ƿ���б�������Tx�˷����>�����мǿtl������<C�I8��F����d��E�Le3�pu�;�f)=T�z=���=%��=�C�=*j}=�!X=�.0=��	=h��<싣<]�<|�<��<,H�<��=��F=�;z=v��=�m�=h��=��=�!�=Tb�=�F�=T6�<�)ۼ*tԽ^W�6���   �   ��
���C��������fʿ"�쿂��C@��Q���4S��R�����)˿Q������F����U���jj������<�p��;�(=vp}=��=���=d�=���=�o=ƙK=j�)=��=|3�<���<,b�<���<��=��;=^\g=�M�=���=�c�=��=Ʋ�=^9�=@��=ݿ�=+�<4`꼷۽3\�`̷��   �   H�Cq@��l���B��A�ƿ���C��V�����w�#�� ���������ǿ�k��y����;C��7�xE��<�d��C�jb3�p��;Rh)=v�z=���=���=�C�=�j}=�!X=�.0=��	=���<T��<d]�<L|�<��<PH�<��=�F=
<z=���=�m�=���=8��=�!�=�b�=pG�=�9�<�$ۼ?rԽ�	W�8���   �   =� ��#6�g�s��2���<����ݿ����j��N����[5�K��q����޿ƽ�}���u�Sh8�w��~��zpT��ݽ`����4<�+=pq=���=[ӄ=T�n=��D=n�=�%�<0$#< �W�p����X��]�xm� 2���&<,e�<.h#=�tc=��=脦=v��=���=IC�=�.}=|��<����I���H�e����   �   ����%�_�s���&��k̿}$��0�������N������"�濭"̿�.���Ԏ�9-`���'�����+���;�d��tc༌��<2�+=Z=`=�j=�S=�P#=���< ��;؞X�&� �aA��mr�p}������-*��pQU��Z�n�� �Q;�~�<��5=�mz=x~�= ��=x��=�u=(2=p�\�����l�0�!̗��   �   k[ʾ0c���D�Z|������
���
ο���W�����5���߿T&Ϳ�L���H���|�B�D���N�̾Y����[��H {��S�<*�'=CD=�4=�=�AO<X�9��������
���p��	�
�"��Ȕ�����Uڽ�R��z�P�P��0��;B=:CP=�.�=.o�=��g=�^=�Dz��}��M����   �   �ɧ�- ��%k&�XW�Y}�� c���\��ֱ����˿�LϿ!h˿�����7��4N��S�����U���%����W{���&V�{����G�`�����<~=bB=D$�<��;(ɼ��t�(ʽB��M�6��,Z���u� H������ �����n��WP��k*��T ����\�1������<��)=��T=DP=�=`��;B,��佻S��   �   Q��ɪþd����/�t�Y� ?���	��`࠿����KT��2���%ٟ��ő����/�W��-�+������4��Z� �7��0�Ӽ�C"<���<d =���<��:�����t������.~6��Wq�h(��0d���¾[aξUҾ��̾���������9��E�c��>(�ǟ޽�rq�P͎�@"g<4�=L�,=V=�V~<T���E����� ��   �   ��B�������о�d	���+���L���i�ZU���s�������憿��~��bg��J��)�!
���̾y���K>���ٽn=� a���u�< D�<���< Y�;��C��T��,O��a���ֶ��޾g ���.��ϑ��7������GؾR���q���B�TJ���݄�`J����E<x�<�==���< �|� �B�.��   �   ����xS��b���̾�� �V����1�R�C��O�+�R�MN���A�1R/�������uƾ�L���{J��q���v��Lu�h�n<xW�<8��<p�@<ܩ���ć�d���|S��e��k	̾� �����1���C�qO��R�<N���A��U/��������zƾ�P��2�J�|{��r�v� vu�Ђn<tO�<`��<p�@<ġ������   �   (>�����`O��^���Ҷ�2޾cd ����{���o���4�����PBؾx���Z��_�B��?��tՄ��1��ȯE<��<�@=d��<��|���B�>���B�������о�f	���+���L�?�i�EW���u��浉��膿��~��fg��J�)�����̾����P>��ٽ�y=�����Dl�<�?�<���<Pr�;L���   �   ����o��Ѱ��y6�bQq��$���_��¾\ξ��Ѿ)�̾s�������f5��u�c��7(��޽Naq�l����Jg<x�=�,=�=�W~<h��������� �����þ�����/��Z��@�����Y⠿����V��u���^۟�ȑ������W���-����	����7��Ϭ �}=����Ӽ�-"<X��< =�<���:�   �   �>�;�ȼ@�t�/wʽL��]�6�&Z��u��C��z���∁�Q�n�JPP��d*��N �����P�1� ]��ի<��)=x�T=�GP=�=`��;D,�J�佤S�I˧�Q"���l&�AW��~���d���^�������˿�NϿ]j˿ݹ���9��*P�������U�[�%���x~���+V�/��D�G� 6 ����<}=�C=`+�<�   �   �=X\O<Ь9����+���G���Y����	�����������mJڽAH��f�P��0��%�;�=�KP=�1�=�q�=��g=j`=@@z�8�}��N�����\ʾd��D��[|��������οk��<����%7���߿P(Ϳ�N��EJ���|���D���d�̾���J�	$���{��L�<��'=hCD=`�4=�   �   �	S=ZU#=L�<@�;0vX�
� �SA�r^r�u�������!���@U��J�,Q����R; ��< �5=xuz=���=���=I��=~�u=�3=�}\�����ּ0��̗��龒�%��_�
����'��l̿�%�Z2�������2��g���ۢ�L$̿[0���Վ�q/`�_�'����
.���;����`o���<P�+==`=  j=�   �   Ԅ=��n=R�D=n�=P2�< B#< }U�]�@aX���\��A��޵�h'<�w�<�p#=|c=��=���=���=���=�D�=�0}=H��<$���I���H�l���U� �*$6�ʳs�/3���<��V�ݿR�������N�;��6����ʺ���޿Hǽ����ִu��i8�������2sT�͒ݽʻ�P�4<�+=:oq=ڶ�=�   �   ���=MD�=�k}=�#X=|10= 
=l��< ��<�f�<���<<�<�R�<��=��F=V@z=t��=�o�=��=���=#�=�c�=yH�=0>�<�ۼ�pԽ.	W�� ���G�q@�pl���B��I�ƿ���c�����H���w����k����`����ǿwl��"��� =C�|8��F��`�d��F��f3�@l�;Bf)=>�z=���=�   �   �|�=�ʊ=�b�=xqo=�kY=ބE=�6=
A-=rs,=�4=�F=�N`='�=	��=b�=���=i�=�F�=���=@�=|g�=�>�=� I=�a�;�Tq�:���܄�oϾ;#��I��f��d����̺�"�ӿ�B翺��Z3�����X�R�ӿ�O���v��a��9�K�����־kь��'��ئ��w��0Ȕ<�6=<�u=q�=�   �   ��=χ�=h�v=�]=:�C=�,=�=�=@/=��=�j%=��@=�d=~W�=b��=��=�!�={��=���=��=�^�=e��=V"K=�q�;�&g�B�� 聾�B˾S��E��P~��������%-п�v㿬�￢������{�[п�������r
��2,H�5��4�Ѿl����a#��������C�<L�7=~t=�^�=�   �   `v=�j=d�K=�T'=T9=�п<�u�<лB<�s$<��9<���<H��<M=f�==VMt=xL�=p��=���=|<�=X��= �=�ٟ=��P=�E<d�I�4&��r�,$��G%
��k;�=q�T<�������ƿ(oؿ,�*迡�gFؿƿٮ������|r�
 =�:T�ݞľ	)����Nj���o���<<=@4p=�ہ=�   �   \1X=�Y2=ƶ =`ȑ<�K;x������,�V�����8*ڼX^���k}�`YG<�~�<�FB=�=�7�=8�=.y�=/��=���=tEX=���<H&��%潊�W��8��5�����*�9�\�����S���/���&ǿ|�ѿÎտ�ѿ��ƿ�ӵ�T��#���v9]���+�`����j��� c�Zu��~d��޾� ��<XA=�$g=�l=�   �   �=��<���;����B��D�k��#������½,cĽlQ�����(yu��\�h��(<��=�Z=�8�=R��=�8�=��=��^=��<4�ƼN�����5��@���7ھ7��kmB�Iyp�X���ѡ��
�������ܽ��U��2x���.���ˍ�ȿo��)B�Q��%�۾nܖ���=�٩ν���PE�;V_=�C=КV=�GG=�   �   ��<PI����?����o��z������>l.�
�:��J=���5�\#%��M��>۽H����#������֪<��4=	x=QҌ=��=��a= ��<@�5օ��	��r�I���x���N�$�<�L�s������ʗ��(���⢿����w��"����lq��*K���#�r����Z��"Gt��.�
�� S��3�<4�=RA=Ԃ;=� =�   �    G��,��尿{`��FT-�9IY�Z������I���Ú��)���܊���s���I�<��ֽ.�w����hKL<*L=�[=��s="Y^=��=Д�;�X$��ҽL*;�Iӏ�_`ʾ���E'�lG�d�w`z�}:��~��%ʃ�j�x�I b�R?E��$����jǾׯ��\�8�-�ѽP�.� �X9|��<$�,=Ծ5=�=���<�   �   nH-������N������������6�վ�⾻��T����Ѿ;�����&p~�r'>��� �N����׼0�<O=��G=&R=ʨ*=lў< W���]�����$�V�ᄚ���ξ�`�)��Z�3�,�E�a]Q�j�T�.uP��@D��1�����f��Hlɾ����KmN��&���'|�h��+�<�I=*�5=��=H��<P(���   �   a����W���]�B_��
x���A��5�v[�.;��� ��K�B��t��8I侪캾����qP�Ϻ������¼PD<^�=��;=z]5=P��< {�;���|��*S���]�x[���s��r<��2�fX�8��� ��H�q�����D��躾#����lP�V��s�����¼�!D<`�=n�;=>[5=4��< A�;���   �   �����V�d����ξ�c�����3���E��`Q���T��xP�DD�ى1����j���oɾĕ�qN�\,��Z/|�'h�'�<(I=��5=��=H��<⣻F<-������&�N�����1��������վ���_��)���Ѿ�
��D����i~�Y">��� �H���׼H�<�R= �G=vR=�*=�ƞ<�g���c���   �   �.;�L֏�3dʾQ��	'�$oG�s
d�dz�U<������˃���x�*b��AE�%�$����OmǾ±���8�� ҽ(/� 8V9���<�,=��5=�=�͒<���,��禽BV��/N-�7BY�q���
���E��g����%���؊���s���I����ֽ��w��
���hL<Q=��[=��s=�W^=�= c�;jb$�?ҽ�   �   ��r�k���n�����$��L�7 s�q����̗��*���䢿r�������.oq��,K�R�#����O\���It�F0�N��X��P1�<��=l	A=��;=v=@(�<����"��N���f���}������e.�P�:�D=��5�C%�~H�%5۽�?����#��w����<��4=�x=Fӌ=��=��a=��<�+�6ۅ�>��   �   FC���:ھ%���oB��{p��Y��.ӡ�\��9���^޽�fW���y���/���̍���o��*B�]����۾~ݖ���=���ν���@@�;�_=��C=��V=LG=x=<�<�H�;߅�"}�~k����|���%�½/YĽ�G������hu��M���g��4(<��=0�Z=;�=���=J9�=c�=~�^=p��<��ƼQ���}6��   �   �:�����O�*�L�\���������v0��(ǿ��ѿ#�տ_�ѿ��ƿԵ��T������|:]���+�m���sk���c��u��d��߾�$��<�A=�&g=� l=�5X=�_2=н =�ّ< �;�n��򤼌�Z�����ڼ�D��@�|�8�G<��<�MB=��=�9�=��=z�=^��=%��=�BX=L؀<�,�E*���W��   �   &��v&
��l;��>q�G=�� ���ƿ>pؿ--�+迄�.Gؿ�ƿ�ٮ�柔��}r�g =�sT��ľ$)����j��`�o�p�<F<=6p=�܁=dy=��j="�K=�Z'=�?=�߿<셇<��B<p�$<�:<,��<x��<TT=��==�Rt=�N�=.��=��=E=�=���= �=Nٟ=*�P=�5<N�I�H(���r��   �   SD˾�S�,�E��Q~�9	��>����-п�w�G��)����0|�G[п������p
��,H����Ѿ���Fa#�(���X����E�<��7=�t=�_�=��=���="�v=�]=��C=�,=�=��=�3=��=o%=��@=~�d=�X�=���=��=^"�=��=���=��=^�=���=�K=�U�;�+g����遾�   �    pϾ�#���I�$g�������̺�a�ӿ�B����^3�� ���X��ӿYO��zv���`����K�L���־�Ќ���'�6צ�(r��p̔<t 6=��u=�q�=e}�=ˊ=�b�=Lro=�lY=��E=86=�A-=�s,=�4=�F=nN`=��=Ԕ�=�a�=H��=�h�=F�=;��=��=�f�=�=�=f�H=@K�;VXq�i��E݄��   �   <C˾>S�>�E��P~����v����,п�v�D�� ����8{�`Zп7��󯜿�	��#+H�O����ѾE���`#�n���P����I�<8�7=̀t= `�= �=^��=йv=��]=f�C=��,=@=ު=�3= �=8o%=��@=��d=Y�=���=��=t"�= ��=��=<��=p^�=!��=f!K=�f�;�(g����Q聾�   �   �#��%
�:k;��<q��;������Uƿknؿ@+�)迓
�UEؿƿخ�����B{r��=�S��ľ�'��x��f�� xo����<$<=L8p=�݁={=d�j=v�K=�['=�@=H�<`��<��B<@�$<�:<���<ܴ�<�T=��==�Rt=�N�=P��=&��=�=�=��=��=<ڟ=��P=F<b�I�$&���r��   �   8��2�����*�A�\� �������.���%ǿ<�ѿj�տ��ѿ�ƿ ҵ��R������[7]��+�x���uh��[�b��r��vd�����`�<�A=:*g=�#l=�7X=�a2=�� =�ܑ<��;�i������&��hڼDD����|� �G<���<4NB=�=:�=�=�z�=>��=x��=�FX=��<�$�X$潡�W��   �   �?��6ھ2��lB��wp�W��]С�N	�����۽�0T���v��&-��ʍ��o�?'B�Y����۾�ٖ���=���ν���p��;�e=x�C=t�V=LOG=6=(�< Z�;Pۅ�|{��|k������ϗ½�XĽ�G�����xhu��M���g��5(< �=��Z=�;�=^��=Z:�=��=:�^=,��<�Ƽ8�����5��   �   H�r�z���
�����$�G�L��s�Z���=ɗ�'��ᢿ����l����iq�(K�J�#�`���?W��
Bt��*� ����?��HC�<��=�A=ʊ;=�	=X.�<�⧻��@���1e���|������e.�"�:��C=���5�4%�mH�	5۽�?��2�#��s��\�<��4=Xx=nԌ=t�=��a=(��<� �zӅ����   �   g';�Tя��]ʾN��4	'��iG�)d�C]z��8��<|��Oȃ���x���a�0<E�H�$�����fǾ����l�8���ѽN�.� �b9X��<�,=�5=�=Ւ<��6�,�`榽7U���M-��AY�M��x
���E��Y���|%���؊���s�x�I� �v�ֽl�w�\	���lL<�R=�[="�s=]^=ȼ= ��;�R$�Pҽ�   �   ���9�V�N���w�ξ�^������3��E�ZQ���T��qP��=D�ك1�����a���gɾ轕�ugN����t|� �g�?�<R=z�5=ڞ=���< ƣ�V9-�Ø��e���N�������������վ���S��#�� �Ѿ�
��?����i~�F">��� ��G���׼H�<�T=~�G=�R=d�*=�۞<�I��0Y���   �   ~v��{O��]�qX���o��8�`0��U� 5��� ��E�c�����?�j亾?���~fP�(��9�����¼0LD<��=�;=�c5=���<���;d���z���R�7�]�B[��Ws��N<��2�\X��7��� ��H�q�����D��躾����lP�3��
���0�¼�)D<��=<�;=0b5=��<P��;���   �   �1-�b�������N�����`}��[���,�վ}����������Ѿ
��ܫ��b~��>�o� �.?��h�׼�<Z\=��G=�R=d�*=�ٞ<LP��5\��@����V�������ξ�`���P�3�%�E�]]Q�h�T�.uP��@D��1�����f��Clɾ����-mN��&���&|��h��1�<�M=N�5=Ğ=���<p����   �   ��
���,�`ঽ_M���H-��;Y�������lA�����*!���Ԋ���s�a�I�����ֽ��w�0��L<[=F�[=J�s=x_^=`�=���;(V$�nҽ�);�ӏ�5`ʾ��8'��kG�d�u`z�|:��~��&ʃ�m�x�J b�T?E��$����jǾʯ��6�8���ѽ��.� 0[9���<N�,=N�5==�ے<�   �   (7�<����jv�#z���]���s��?���_.���:�R==�J�5��%�[B�*۽ 6����#� �����<|�4=6x=�֌=!�=��a=���<��Յ�F	���r�"���U���B�$�4�L�
s������ʗ��(���⢿����x��"����lq��*K���#�l���yZ��Gt�X.�}��pO���8�<^�=`A=L�;=T=�   �   D =��<��;(Ʌ� p�ok�2��;���U�½OĽ�=�����`Vu�J=�0�g�Xh(<��=��Z=?�=��=Z<�=^�=��^=��<��Ƽm�����5��@��f7ھ+��dmB�Cyp�X���ѡ��
�������ܽ��U��4x���.���ˍ�ȿo��)B�P���۾eܖ�q�=�n�νF���V�;�b=��C=P�V=�PG=�   �   �9X=�d2=P� = �<@@�;D��ڤ���弖~�j����ټ\)����{�ȱG<l��<RWB=��=4=�=�!�=�|�=� �=���=tHX=<�<�$��$�K�W��8��!�����*�4�\�����T���/���&ǿ}�ѿŎտ�ѿ��ƿ�ӵ�T��"���t9]���+�[����j��� c�6u��}d��Ҿ����<�A=�)g=$l=�   �   �{=�j= �K=\_'=�E=��<Ԕ�<(�B<�$<@0:<(��<���<�\=��==�Yt=�Q�=���=Z��=`?�=���=��=B۟=��P=hK<R�I��%���r�$��>%
��k;� =q�S<�������ƿ)oؿ ,�*迢�jFؿƿٮ������|r�	 =�8T�؞ľ)����j��8�o�d�<(<=J7p=�݁=�   �   ��=���=��v=�]=B D=��,=6	=H�=�7=6�=hs%=(�@=��d=�Z�=f��=���=�#�=@��= ��=<��=d_�=	��=H#K=0w�;`&g�&���灾�B˾S��E��P~��������%-п�v㿭�￤������{�[п�������r
��4,H�4��2�Ѿh����a#���������TD�<b�7=�t=�_�=�   �   t`=�)\=P�T=اL=&�F=\�C=�D=�J=ZV=�
h=N�=�K�={%�=y�=�*�=���=n�=i��=l\�=���=H��=ts�=y��=4Y
=��J|���;0�It���J׾0��@��n����$��È��qf���ʽ��f��r����I���ݍ�%�o��aB��{���ݾvę��F����,�N�p����F�<L9=��H=p�[=�   �   �<\=:�U=�)K=�4@=��6=�1=}/=�q3=��==.oN=.�e=n��=���=j�=jκ=���=�U�=*��=�,�=3��=K��=�ο=��=<U=��l������+�1N��� ӾUc�8=��j�����]��B���O@��͓���:��v����{��Z��x�k�V�>�i���ؾK���@�I8ܽFCD� k�����<�2"=�uI=<6Z=�   �   �P=�eA=�!.=�=.7=<;�<���<��<$��<,��<��=�v8= p`=���=�S�=rR�=���=��=nv�=��=h,�=Z��=���=>�=xA�vk��P��4-��Ŏƾ'B	�*	3��=^��`���ڤ�I���;��A��V���\T����� �^��!4���
���˾�6��{2�P�ƽ�#%������<�e*=�BK=$NU=�   �   H�9=�6=���<܉�<�2O< ��;��5�p���`���@���q�;h�W<���<�=��Z=nq�=|�=��=��=��=�J�=:q�=�U�=�V*=�5��t�s�J�?�m��+���$��#��K�N�q�ԉ�p6��9�����������񖿘����;q��K�u�#��@���ƶ�9y����$ܤ��@� 5�;��<N�5=2)L=0K=�   �   &�=L��<��7<`NY�����+��$K+��TJ��X��ZR��?8���
�<%�� ^�D?�<�h=�>i=�l�=P��=�S�=wq�=N�='�=�==(�<�'1�;�-J������پ4��Č2�lU���s��Å�o^���䏿:���W��Q�r��T���1���Zpپ u��J5Q�y���r�s�0`]�p��<��=$YA=HII=��8=�   �   � �<@��;��v�
��Qt��(����ɽd�%��"U��0��gɽ]F�_�t���ܲ��K�<��>=��=:��=��=y`�=�=�.P=��<��ϼyT��C?"���~������/���U�4��O�7�c�R�p��?u�Tp�)�b���M��%3�p�S��:_���}�_[$�f���$� �S;��<�@4=��I=�s?=J�=�   �   ��;@K����L�BE��wl�7��M�1���F�hCS��U�RM�*�:��) �>X���t���SV��g��JX<d�=
o=��=��=���=0�^= �<�>���Ng����pF��ޏ����FR��M��A)��K:��6E�f�H��vD���8�� '����8������틾>@��v�\Af�(@:��C�<dL%=��K=tWL=x�+=�i�<�   �   �/��jqZ�[���j��s=�>�j�@��������l���ǖ��I���(���(X�J�'�d�뽈[���M�0��;�r=VH]=NU�="�=��f=L=h�<|u������(��"�X��œ��μ������?��.x�6*�����-���޾�Y��R��>K��k��U��W���}M<$�=��N=�D]=�F= �=��C<�   �   HA>��^����HU�N��1먾�ľ"5پ�c澤:�nI�վf���|��������B�M��`;��8��;��=>\S=�p=��f=�5=���<@�컰6>��W����BU��J��E稾Tľs0پ�^��5��D侵վ����y������0�B�����5�� �� 9�;��=>^S=��p=x�f=�5=���<����   �   $���>��]�X�ɓ��Ҽ� �侓������z��,�-����R����޾�\���
���AK��n�Z��Dc��mM<��=�N=FE]=�F=�=XD<���eZ�|S���e�En=���j�o<��������T~��Ԓ����������"X�n�'�|��GU��l:����;�w=�K]=V�=�!�=��f=��= �<8����   �   ���ruF��᏾z ��V������)��N:�f9E�<�H��yD�*�8��"'����m�ﾮ����A@�@{뽀Gf��P:��>�<6K%=��K=�XL=��+=�s�<�!�;d8����L��=��`c���l�1���F��<S�i�U��KM�+�:�_$ ��N���l��dFV��R��xjX<V�=$o=��=U�=4��=��^=�< v���Xg��   �   �B"�I�~�����T3����ȭ4��O�
�c�.�p��Bu��Vp���b�٬M��'3��q����a���}�c]$��h���(�@�S;���<�@4=��I=v?=�=l�<pڹ;@�v�X���Bt�� ����ɽ������J��1�彠]ɽ�栽Lx_����@����\�<P�>=g��=Τ�=��=�`�=y�=�+P=4��<��ϼ�Y���   �   �0J������پ���؎2��	U�=�s�CŅ��_��揿s ���X��D�r�� T��1�����qپOv���6Q�������s��g]�t��<��=�YA=�JI=.�8=�=��<��7<@�X�tP���=+�FJ��X�FKR��08���
���� A[��R�<�p= Ei=%o�=��=�T�=�q�=�M�=4&�=��==��<\/1�x��   �   ��m�.��Q'���#��	K�\�q�(Չ��7��X������������`����<q��K�A�#��A���Ƕ�Xy�?��ݤ��B��0�;��<��5=\*L=K=�9=t:=��<l��<�PO<0��; �3��T��@j�����pƂ;h�W<���<��=��Z=Mt�=��=��=2��=< �=K�=�p�=U�=�S*=@ա���s����   �   �.����ƾFC	�}
3�R?^����`���ۤ���f<�����𾤿�T��K����^�)"4��
��˾�6���2�w�ƽ�#%����t�<(f*=�CK=�OU=�P=thA=P%.=2�=<=lF�<D��<`��<��<��<l�=�|8=�u`=K��=�U�=<T�=���=��=w�=8��=R,�=ઽ=���=,�=�S��n��u���   �   KO���Ӿ&d�9=�рj�+��C^��ǌ���@��7����:������
|��%Z����k�P�>�U����ؾ�J����@��7ܽ�AD�b�����<�3"=�vI=p7Z=>>\=�U=�+K=L7@=�7=�1=j�/=�t3= �==�rN=r�e=���=��=��=^Ϻ=���=V�=���=-�=!��=���=1ο=��=~R=��l�6�����+��   �   �t���K׾�0�p�@���n�O���X��爰��f���ʽ��f��O����I��Kݍ���o�paB�\{�(�ݾ�Ù��F���n�N�P���XJ�<�:=ԨH=l�[=L`=v*\=�T=��L=�F=��C=��D=~�J=�V=h=V�=�K�=X%�=�x�=P*�=���=�=��= \�=(��=���=�r�=���=�V
=���,~���<0��   �   uN��� Ӿnc�!8=��j�����]������?��g���:��􍭿V{���Y��p�k�d�>������ؾ�I��;�@��5ܽ�>D��O��l��<V5"=�wI=�8Z=p?\= �U=�,K=88@=j7=�1=�/=vu3=��==�rN=��e=��=��=��=sϺ=���=3V�=���=<-�=P��=C��=�ο=Y�=.T=�l�x�����+��   �   	-��u�ƾ�A	��3�E=^��񃿉_��Hڤ�����:��n ��|����S������^�g 4���
���˾95��"2���ƽ8%��}��&�<.i*=TFK=RU=�
P=�jA=<'.=��=�== I�<d��<0��<p��<8��<��=H}8=v`=j��=�U�=XT�=��=��=Vw�=���=�,�=���=ऐ=r�=�@�Mk��"���   �   $�m�&+���#��P#��K��q�NӉ��5��=���w�������{𖿀����9q��
K�ғ#��=���Ķ���x�����פ��2��b�;� �<�5=".L=|K=6�9=Z==`��<(��<YO<��; "3��J��pb������ʂ; �W<���<J�=��Z=xt�=��=��=���=� �=�K�=�q�=�V�=LX*=@��R�s����   �   f+J�y���Cپ(��o�2��U�͏s���:]���㏿���DV��ʓr��T���1����Nmپ�r��f1Q�g�����s�`A]�|ē<��=�^A=\OI=B�8=��=��<@�7<@�X�x鐼���;+��DJ�~X�lJR�b08�8�
��
�� +[�xS�<,q=�Ei=vo�=���=FU�=�r�=NO�=!(�=J�==P�<4$1����   �    ="���~�����3-���z�4��O���c���p�=u�BQp�Z�b���M�]#3��m����\���}�_W$��_�����wT;(��<HG4=:�I= {?=^�=��<0��;p�v�<��D@t�i����ɽ��Q��hJ�����b]ɽ�栽�w_��� }���]�<��>=���=}��=��=b�=��=�1P=���<p�ϼJQ���   �   Z���mF��܏�R��O��_��)�eI:��3E���H��sD���8��'�Y����l����ꋾ9@�o��4f�X:�XT�<�S%=��K=�^L=��+=�|�<�B�;�0��0�L�'<��b�`���1�0�F��<S�1�U��KM��:�E$ ��N��pl���EV��Q��@mX<J�=~o=��=��=c��=�^=�"�<����Gg��   �   �����X�LÓ��˼����������u��'�ߒ�x������޾�U�����Y8K�Dg�lN���?���M<T�=:�N=L]=� F=��=�D< ��bZ��Q��;e��m=�'�j�8<���������>~��Œ����������"X�Z�'�I��U��(9� ��;�x=pM]=�W�=$�=��f== �<`f���   �   *->��Q����!>U��G���㨾f ľ,پIZ��0��?��վ���u��(���'�B�����-�����@��;��=fS=�p=��f=,�5=ē�<|�3>�V����FBU�uJ��稾&ľR0پ�^��5꾾D侭վ���y�������B�����5����B�;Z�=�`S=t�p=�f=�5=���<�`��   �   X���ZZ��L���a�.i=���j�9��������2z�������������X�m�'�.�뽥L���@*�;$�=�S]=�Y�=�%�=B�f=�=X�<xn��j���t����X��œ��μ�|����2��&x�0*�����+���޾�Y��J���=K��k�cU���T����M<|�=2�N=�I]=�F=��=p'D<�   �   �`�;�$��ƩL�~6���Z����̀1�f�F�B6S���U��DM���:�B ��C���b��t5V�6��X�X<J�=�o=��=��=���=�^=�!�<�#���Kg����]pF��ޏ����R��>��6)��K:��6E�b�H��vD���8�� '����3������틾�=@��v뽀@f�;:��G�<JO%=��K=f]L=ƻ+=l��<�   �   ��<p�;��v����5t������ɽ�彞��E@�����sSɽEݠ��f_�����ٯ��s�<�>=�Ą=Z��=��=�c�=��=�2P=���<t�ϼES���>"��~������/���H�4��O�3�c�O�p��?u�Tp�+�b���M��%3�p�O��3_����}�A[$��e���#��T;���<D4=n�I=�z?=`�=�   �   \�=��<��7<`/X�ِ� ��� 0+�P7J��W�Z;R�!8�X�
����W��j�<6{=Ni=�r�=_��=�W�=�t�=�P�=�(�=�== �<�%1�P
佸,J�}����پ'����2�dU���s��Å�o^���䏿<���W��S�r��T���1�~��Vpپu��45Q�9�����s��[]����<D�=�\A=~NI=��8=�   �   ��9=4?=`�<���<`oO< =�;�1� ��0�� E�` �; �W<���<|�=L[=x�=�=l�=���=u"�=(M�=s�=ZW�=8Y*=�����s�����m��+���$��#��K�L�q�ԉ�o6��:�����������񖿚����;q��K�s�#��@���ƶ�*y�n���ۤ��>�?�;��< �5=�,L=@K=�   �   �
P=^kA=�(.=b�=�@=tQ�<`��<���<���<� =��=�8=||`=l��=�X�=�V�=9��=��=�x�=���=�-�=���=���=��=�<��j����-����ƾ!B	�%	3��=^��`���ڤ�J���;��B��W���_T�������^��!4���
���˾�6��j2�)�ƽr#%� v�� �<6g*=
EK=tQU=�   �   ?\=��U=J-K=
9@=�7=@1=�/=�w3=l�==vN=�f=���=���=.�=�к=���=jW�=���=..�=*��=��=\Ͽ=)�=�U=@�l�`�����+�'N��� ӾPc�8=��j�����]��B���P@��Г���:��v����{��Z��w�k�V�>�h���ؾK�� �@�78ܽCD� h��ȫ�<�3"=�vI=�7Z=�   �   L��<��<��<�o�<�&=dE=�x-=V#G=ھc=�k�=)�=Eѣ=P)�=*��=�,�=2�=�Q�=�G >�>? >�?�=$ �=�X�=�5q=̣<�/�ʽz�:�Rz����;};���*�|pL�yOj���z������z��������j��M�l�+��
�?oӾ6ř�9�R��n��f���O�С��Q:<�}�<Xu�<,K�<�   �   ���<t��<t��<�s�<���<J�
=&�=�|6=F�Q=V�o=E��=�t�=�G�=\\�=��=���=���=G%�=a >���=��=4R�=�t�=J{s=�q�< ��;�ý�m6�:^��$�ɾ�����'�ͺH�$f��M}�������F��mO}��Kf��6I�צ(��G���ξ�J��=;M��Z�C'��p*��`0m�@]S<pS�< n�<8�<�   �   ���<p	�<P��<���<`�<�"�<TY�<\T=$=��5=ރV=̺{=#5�=�w�=l��=(j�=���=���=�8�=�=�X�=+��=[��=��y=���<tUżOⱽCl)��a�� ٽ��)��_�r�=��Y�`p��~��v����}��o�>�Y�2>�r�g���5#¾�2��@�=��L�{����� 1�:Ж�<��<d��<(��<�   �   ���<�|�<��<p�L< T <��<h[
<�7(<ءe<�%�<�E�<=r@G=��y=_��={�=0��=��=�Q�=��=�2�=���=�=$.�= ��<�<|�ZJ���[�H�n��g��[�侣,��!-���F�!9[��/h��l���g��Z�,qF�2�,��+�_��o����x��t%��ŽhC��O��X*<�L�<�$�<0� =X7�<�   �   ��<��m<"�;@,&� �$�X脼4����㵼�&����������:(�{<,��<>?=n�=���=w�=���=2*�="��=(��=|��=ԃ�=� =���./h�����&L��=���$Ǿ�!�������.���@��BL�#P�t�K��@���-����:����Nƾ6����	Q�����������@r�:�ݬ<v�=*=�=�+�<�   �   ��<0[�;X���Ƽ�&��<O��&x�yd�� ׍��L����p��=�P~�)��L-<<=��Q=x<�=�;�=0��=z��=��=��=}��=�M)= p�;,�������%���t��'��_�Ӿ�����u�6�"��,���/��,���!����v"����Ͼw⢾�Bp�$���ǽ�B����,�<�
=zx'=��+=��=���<�   �   H�<�&�V� ��\�[��qlŽ����T�����*�N����߽�M�������w�P�����<z�+=�z=ƙ=�j�=�ӭ=r�=��=��==�^�< է��O���N����@�p���쩾1FξƔ��h��l���ha�#���Ⱦ�У�NV|�2�4��5�/}�P
��X�:<=48=n�I=p�?=�C= o�<�   �    �i�����|w�SǼ�M���Ũ�-�9�R<N�� Z�\�[���R���?���$�H-����d��\���  <T�=R#c=O��=�$�=��=��=��K=��< %���.�����ŭH�����ڞ�|P���0̾F�ؾ�ܾ�U־��Ǿ���H���r�J�4������D���	ۼ�/�;&�=:�E=�$f=8�g=t�L=�=�<�   �   1��:g���Ž/��<�4h��#��]敾�֞����������A����}�(�R�2j#�@U潢����:⼰��;D�=�R=��=\��=��}=�Q=T�=(Y<H#��r0g���Ž$+��<��h�� ���╾Ӟ�����v���k>��Ի}�&�R��e#�]N�&����)⼰�;�=��R=�=���=��}=�Q=��=pF<�   �   �.������d�H����-ޞ�T��v4̾G�ؾ�ܾeY־�Ǿ����Lr��4�����\I���ۼ��;`�=��E=F#f=��g=�L=�
=�< Ji����@�v�����N������9��6N��Y�Z�[�ҹR�(�?���$��(�缽��d�8I���> <�=�'c=ʇ�=�%�=�=��=��K=���<@S���   �   �T��&U����@��r���奄�Iξ�������9n��!�Ic�~꾾�ȾJӣ�&Z|�6�4�p:� 6}����8�:<Z=D28=��I=r�?=�D=t�<h�<��%�P� �n\��T���dŽL��;P����&������߽�E���ـ��k�0���4�<�+=�!z=�Ǚ=(l�=,ԭ=|�=P�=6�==�U�<X⧼�   �   ����i�%��u�F*����Ӿ+����w�Q�"���,���/��,�f�!�K��F%���ϾN䢾zEp�-$�Íǽ@B�(���'�<�=Tw'=|�+=Z�=���<|"�<�}�;xl�H�ż��p1O��x�_]���ύ�E��"�p�t=��d��(�(t-<@D=*�Q=?�=�=�=���=V��=��=j�=���=�J)=�G�;p���   �   	����)L��?��K'Ǿ�$��r����.���@��DL�P�O�K�y@�A�-����F���ePƾo����Q�ئ�찖�Ԫ���.�:�ڬ<Z�=�=�=�-�<4��< n<�D�;@�%�p�$�Hׄ��y���ε�L���ꇼ`b��1 ;(�{<���<�?=��=8��=y�=.��=2+�=���=<��=��=Ղ�=$=�H���6h��   �   0^�j�n��i�����.�#-�|�F��:[�r1h���l�u�g�o�Z�[rF�,�,�],����R����x��u%�C�ŽDC�x�O��T*<|K�<�#�<.� =d8�<X��<���<��<`�L<8h < 	<�v
<�U(<��e<6�<pU�<�=hGG=��y=��=N}�=���=
�=�R�=���=�2�=]��=~�=-�=��<`Q|��M���   �   \n)�@c���ڽ�|+��~����=�]�Y��p�1!~��w����}���o��Y��>�������#¾23����=�{���{�T����%�:X��<d�<���< ��<,��<8�<X��<��<��<�*�<Lb�<JY=B=��5=��V=��{=\7�=�y�=��=�k�=՛�=P��=$9�=\�=�X�=ֲ�=���=|�y=��<�^żt屽�   �   \o6�=_��\�ɾB��\�'���H��f�}N}�8��]�������O}��Kf��6I��(��G���ξ]J���:M��Z��&���(���&m�8_S<DT�<�n�<l�<���<h��<�<�v�<���<� =��=�6=�Q=��o=���=�u�=�H�=@]�=���=(��=\��=�%�=a >���=���=�Q�=�s�=4ys=�k�<�����ý�   �   ��:��z����;�;�,�*��pL��Oj���z������z��������j�DM��+��
��nӾ�ę�5�R��m��e���M�����@V:<��< w�<�L�<���<�<p��<(q�<�'=�E=y-=�#G=,�c=�k�=1�=<ѣ=<)�=��=�,�=��=�Q�=�G >r>�> >�?�=��=X�=�3q=�ǣ<�2��ʽ�   �   n6�h^��H�ɾ�����'���H��f�TM}������������N}��Jf��5I��(��F���ξzI���9M�}Y�%��d#���m�PgS<X�<�r�<��<<��<� �<��<�y�< ��<z=p�=>�6=z�Q=l�o=���=�u�=�H�=Y]�=���=:��=r��=�%�= a >���=܎�=R�=Wt�=�zs=�o�<�����ý�   �   �k)��a���ؽ��(���~���=�V�Y�yp��~�_v����}���o���Y��>�Q�f����!¾�1����=�l��x�{��~��@��:��<��<l��<���<���<P�<���<��<���<�.�<�e�<�Z=d=��5=��V=0�{=�7�=�y�=F��=�k�=���=���=d9�=��=dY�=���=���=�y=L��<�Tż�ᱽ�   �   �Z��n��f��,���+�� -���F��7[�7.h�D�l�9�g�Z�Z��oF���,�+*����[��J�x�r%���Žb�B�`�O�0m*<XV�<�-�<�� =�A�<��<��<��<��L<�t <	<�
<�](<��e<x8�<HW�<N=�GG=t�y=D��=�}�=3��=L�=ES�=���=�3�=D��=��=�.�=H��<�4|�I���   �   ����$L��<��#Ǿ���u��F�.���@��@L�.P�s�K��@���-�������Lƾ굔�Q����)���L����F�:��<��=�=�=�8�<č�<n< j�; �%�H�$��Є�Tt��4ʵ����0臼@^��> ;��{<���<:	?=0�=z��=_y�=���=�+�=p��=N��=���=��=J#= ���*h��   �   ������%���t��%���Ӿ����/t�[�"�{�,���/�w,�j�!�������r�Ͼ�ߢ��=p�(�#�S�ǽnB�����:�<0=�~'=&�+=� =��<.�<p��;X��ż���-O��x�%\���΍�ZD�� �p� s=�Pc���(�@v-<�D=��Q=l?�=^>�=*��=&��=�=�=��=rQ)=В�;����   �   �K���I��_�@�n��9ꩾACξb���[���i�^�J_�$�3�Ⱦ�ͣ��P|���4�?.��"}�<����;<V=�:8=�I=V�?=`K=\��<س<��%�&� ��\��R��4cŽ��轢O�f���%�M���n߽�E��Tـ�4k����<�<��+=�"z=cș=�l�=dխ=8�=��="�==i�<<ȧ��   �   &	.���������H�Q��؞�7M���,̾]�ؾ�
ܾxQ־��Ǿ��� ��� r�$�4�9����=��\�ڼ�|�;J�=v�E=�+f=�g=��L=
=���< �h�����L�v�����`���C��6�9�6N���Y��[���R���?���$��(�A缽�d�(H���A <��=�(c=���=�&�=��=�=��K=0��<��   �   p��(&g�]�ŽW'���<�Mh�����ߕ��Ϟ�M����:��2�}��R��`#�)E�c����� e�;�=>�R=�=B�=��}=2Q=&�=o<����+g�p�Ž&*�:�<��h�e ���╾�Ҟ�����]���Z>����}��R��e#�&N�꓊�l(⼰�;$�=�R=B�=}�=�}=�Q=�=�t<�   �   ��h�������v�幼�;���t����9��0N���Y��[���R��?�
�$��#�O޼��zd�H.�� l <� =�/c=S��=�(�=H�=��=��K=P��<p���.���� ��H�a���ڞ�?P��e0̾!�ؾ�ܾ{U־s�Ǿ���?���r�4�4������D��Xۼ�6�;n�= �E=�'f=�g=��L=`=d��<�   �   ��<@�%�� �n�[��M��]Ž���|K����� ������߽�<��р��\��D���+�<��+=�)z=R˙=Po�=!׭=}�=��=��==�g�<�̧�N��M��ә@��o��h쩾�Eξ���t��\��l���da����Ⱦ�У�:V|��4��5꽀.}������:<�=d68=��I=�?=:J=\��<�   �   T/�<P��;�I�4�ż|��$O��x��U���Ǎ��<���p�Vd=�,G�ذ(�Ф-<�N=f�Q=	C�=XA�=���=��=��=&�=���=�Q)=p��;ޗ����\�%���t�X'��*�Ӿ`����u�,�"�w�,���/��,���!����q"����Ͼm⢾�Bp��$�P�ǽ�B����</�<�={'=��+=�=�
�<�   �   ���< n<`|�;�Q%�`�$�XÄ�d��l������� ҇�1��� ;P|<X��< ?=�=���=7|�=���=�-�=���=~��=x��=���=�#=����,h�ǩ��&L��=���$Ǿ�!�������.�}�@��BL�!P�t�K��@���-����5����Nƾ0����	Q�l������У��@��:��<t�=
=�=�6�<�   �   0��<���<��<�L<p� <�*	<x�
<xw(<��e<�G�< g�<,=�OG=��y=���=]��=���=e�=U�=l��=�4�=@��=��=a/�=���<�4|�rI��c[���n��g��<�侖,��!-���F�9[��/h��l���g��Z�,qF�2�,��+�[��j����x��t%���Ž�C�8�O��\*<�O�<�(�<� = ?�<�   �   0��<��<���<���<h��<�3�<Hl�<�^=�=��5=��V=.�{=:�=L|�=h��=�m�=���=���=�:�=��=TZ�=E��=L��=P�y=t��<�Rż�ᱽl)��a��	ٽ�s)��X�m�=��Y�_p��~��v����}��o�?�Y�2>�r�d���3#¾�2��8�=����{����� D�:���<(�<��< ��<�   �   ���<���<��<(z�<0 �<x=��=�6=|�Q=��o=匈=7w�=&J�=�^�=���=F��=n��=|&�=�a >���=���=�R�=u�=|s=�r�<�����ý�m6�.^���ɾ�����'�˺H�$f��M}�������F��mO}��Kf��6I�֦(��G���ξ�J��5;M��Z�''��*��@+m� _S<�T�<�o�<��<�   �   l�����P�|��Y	��g�: wG<���<�=8zK=��}=3?�=Hc�=n)�=":�=N%�=1b�=$�>Ȯ>�8>��>�@>�a�={��=X�=��I=�&<"���ν��2�l�����������!���2���=���A���=�H�2�!�!��{����ι�=���EkK�z��e����Z��{ ��I��`p��mq��+��HM���   �   �W��4]�� x���� �%9D/<��<�Q=*�?=�p=v��=��=��=��=���=Nv�=J� >@�>��>R�>�k >
N�=��=�K�=�5L=@�9<�F��ɽ�.��(��}K��)n��%	�ވ��w/��T:�N>��L:��x/�����	�����̵������-F����𡬽�LO�|v�t���p8O��uR��{����   �   x_���e���^n�p��`3� ��;|��<�r�<<�=&I= �w=�=���=뀿=���=��=�?�=���=�\>�>���=&��=��=��=�]R=��m<z6��J��^�"��t�̦�xoվ�m�	����%�s0��3��/�̜%�Ҡ����;�־9,��X7��z�6��j��!��~.�D�����2�`>��}�H8+�X�d��   �    �@��g� �k��)K��j	� �-� �;h�Q<Ȩ�<��=( 0=6�^=y��=r��=��=�+�=Xw�=d��=��=�,�=���=��=5x�==B�Z=��<`CƼU����g��[�X���xT�����]��� ��:#����Y=�Fz��꾽B�����O�b��8��VϽt�x���(�6�� ���4; �W:��H��#���   �   �d���F�ࠁ�H���L	�� ���H&X���@}ʺ���; +�<�U�<�,+=��b=*K�=��=9�=v��=F(�=���=L�=��=���=�0�=l_b=��<Ho�BT�����%<��h��v&����̾E�������%���c���U ��/ʾ�ѥ�m���_=���eÞ�� %���c� \4; [8<�[<8O3<p̼; ���   �    I���E�Ȳ��<"߼�}�h`���P��D����d���`i����<�p�<+=T|n=ߕ=ӯ=B��=B��=���=���=e�=
4�=6�f=T>�<�\��Z~=���½4W��^X��F��`���Ǿ��ܾSl�6��y��p�پ��¾�]��&󆾡zN�������N� ������;`*�<�F�<��<ظ�<�Vs<���;�   �   @zɺX�x�����,�_���n��*����v��_������rP���	�h�`����;�9�<��C=�_�=B��=x9�=�&�=p��=.U�=���=>/e=��=�F�;�z���H��@��1�+�)`��U��V���>���ӻ��ž��������&B���P��H�M�B���ͽ�Rk����0;�;���<~�=��!=Fw=�k=���<��;<�   �   �U�p��B�/�`���׫���ѽ���tn�|�����?;۽bx��b�{����?���<t =�9i=L�=⍞=p�=�= &�=�$[==B+<�Z��H�Q�.���H��.+��;R�Bkt��T��](���ː�������b�?�:�Z��9hȽhQm�к����;���<Ģ0=�+R=/Z=��K=�*=�3�<p�i<�   �   �C����F������2�����a1�G�C���M��FN�WE�v�2��{�������M��╼�X < M=��L=~�z=�ʇ=�q�=J6t=�qG=��=pUe<�6����C���������>��X]1���C���M��AN�wE��2��w�З��z����M��ѕ��s <�R=��L= �z=(̇=�r�=�7t=rG=v�=�Ne<�   �   d���Q��2���K�H2+�f@R�8pt�{W��/+��~ΐ��������xb�>�:�����mȽdZm�l޺��^�;H��<�0=�(R=�,Z=��K=�*=�2�<0�i<��U�ph����/�\���ҫ�e�ѽ��{�Rj��w�a���m3۽Eq����{���p���<z =�>i=8�=g��=��=��=�&�=f$[=�= 7+<�   �   (����L������+�<-`�[X�����/���ֻ��Ⱦ����L����D���R����M�����ͽ�Yk����p�;���<@�=��!=�t=�i=��< �;< [ɺ��x�����,�>	_�2��fh��簞�p������[��fP���	�HY`����;�H�<&�C=ob�=O��=;�=(�=J��=�U�= ��=h.e=��=@)�;�   �   ��=�A�½Z�qbX��H���b���
Ǿ��ܾjo�H��d���پ7�¾�_����V}N�. �}���h�N�����d�;4$�<A�<,��<̴�<�Ps<���;�I���E�����߼x�:Y����������|�H���@���<l��<~�+=��n=��=2կ=��=���=��=���=Le�=�3�=��f=�8�<����   �   �Z�+���(<��j���(��N�̾���]��9�����Je�Q��}"뾳1ʾOӥ�����a=���Ş�h%���c�@14;0Q8<X�Z<�F3<о�;�>��h��F�𝁼�z��\���w���X�(�� �ɺ��;;�<he�<�3+=^�b=N�=���=;�=��=�)�=���=��=8��=���=_0�=�]b=P��<("o��   �   �����i�b[�����lV��/�꾎�#��K �<#����Z>�#{�#��C�������b��9�*XϽ�t�������6��<�� ;�:W:@�H��,����@���g�(�k��"K��`	� �-��9�;p�Q<���<*�=�0=��^=��=ì�=��=�-�=�x�=���=���=H-�=��=���=�w�=V��=�Z=0�<�LƼ�   �   �M��9�"��t�~ͦ�qվ�n������%�b0��3���/�z�%�a��o����־�,���7����6�Fk�����.���� �2��F�P�� <+�P�d��`���e���\n� �� �2����;(��<$y�<��=�)I=��w=��=N��=n��=ز�=2��=r@�=M �=�\>>���=���=���=f��=Z[R=�m<�:��   �   #ɽa�.��)���L��Ho�&	�z��dx/��U:��>�:M:��x/�4����	�����̵������-F�c�������LO��u�d����8O�pvR�(�{�T���W���\��x���� �&9�I/<��<DS=�?=��p=a��=⢧=ʡ�={�='��=�v�=r� >Y�>��>O�>�k >�M�=f��=�J�=�3L=(�9<J��   �   S�ν��2�����~﴾!��E����!���2���=���A���=�#�2���!�H{�]��yι�����ljK����d���Z�:z �tG���p��jq�0*���K��H��д����|�W	��y�:xyG<���<��=�zK=�}=<?�=Jc�=a)�=:�=+%�=b�=�>��>�8>m�>^@>a�=���=��=�I=8�&<�"��   �   Hɽ,�.��(���K��n��%	�����w/��T:��>�TL:� x/�j���	�����˵�ǰ��J,F�N��ٟ���IO��p�T���(/O��lR�h�{�t���S��(X��xx���� `(9�O/<���<ZT=�?=��p=���=��=���=��=@��=�v�={� >f�>�>b�>�k >�M�=Ʉ�=bK�=5L=H�9<dG��   �   J����"��t��˦��nվym�|��B�%��0�1�3�*�/�כ%�ߟ�����־�*��6��e�6�$g��B혽z.�ȝ����2��!�Pa�h)+���d�TW���\��0Ln�����2����;0��<L}�<p�=+I=��w=K�=���=���=��=Y��=�@�=| �=�\>(>��=���=^��=`��=^R=X�m<�5��   �   ����~f�F[�o���RS��������� ��9#����<�y�o꾱@����D�b�I6�nRϽ

t������6��e�� �; �X: XH�����p@�@�g���k�hK��M	��-��U�; �Q<<��<�=:0=��^=t��=��=�=�-�=�x�=ƺ�=2��=�-�=���=���=�x�=���=��Z=���<8>Ƽ�   �   LO�����#<��g���$����̾����i�����wb������L-ʾ�ϥ�k��[\=�� ������$�ȷc� �4;�q8<�[<(f3<���; L�@+�p�F�܏��n�� ����m����W�`���/ɺ %�;T>�<�g�<�4+= �b=TN�=δ�=`;�=b��=�)�=c��=��=��=��=2�=4bb=<�<�n��   �   �w=���½�T��[X��D���]��HǾ˾ܾ\i���O��T�پ��¾7[������tvN����<{��H�N�\s��`��;p7�<�R�<��<�Ų<�rs< �; �H�H�E�\���߼�q��S�����������伬���@��@<$��<.�+=@�n=��=�կ=J��=
��=���=���=�f�=�5�=��f= G�<3���   �   <l���D������+�@%`��S��ͨ��p���л�v¾�񆹾����:?���M����M�)��%�ͽGk��鴼 ~�;4��<8�="�!=�}=�r=��<�<<@JȺ��x�����,�_���$f������n��`���y ���dP�̆	��U`�`��;@J�<��C=�b�=���=�;�=�(�=C��=W�=�=�3e=�=pw�;�   �   K���Q��(��IE��*+��7R�Pft�R��z%���Ȑ��)��mb�B�:����`ȽJDm�𹺼 ��;���<��0=T2R=�5Z=j�K=$*=�C�<�j< 	U��X�� �/��X���ϫ�װѽ���z��i�Rw������2۽�p�� �{�F����<�z =z?i=��=��=��=&�=f(�=�)[=�=�\+<�   �   H�F{��=��;������'���X1���C�k�M�<N�
E���2��r�ڎ��r��ܯM����h� <<[=|�L=Ԫz=bχ=�u�=v>t=pyG=��=xte<P�r}��?������4����d\1�ˍC��M�
AN� E���2�iw�~��z��4�M��Е�Pv <BS=��L=<�z=͇=�s�=;t=�vG=��=(qe<�   �   �U�PV��,�/�2V���˫��ѽ�
�^w��e�2s����u*۽�h��Rt{����� ��)�<� =zFi=��=���=��=��=�)�=�+[==X]+<�M��
�Q�+��=G�i-+�;R�sjt�uT��(��zː������
���b��:�:���gȽ�Pm�Ϻ����; ��<ܣ0=$-R=D1Z=��K=*=�>�<�
j<�   �    kȺ�x��켖�,���^����va������ih����������"WP��y	��%`��Q�;p]�<�C=Pf�=���=(>�=�*�=
��=�X�=ĕ=X5e=��= u�;�o��YF��܌��+�#(`��U����� ���ӻ�vž��������B���P��-�M�(���ͽJRk������@�;T��<��=x�!=�y=0o=4��<h
<<�   �   �H���E�8����߼>n��N���������@��\���`���0@<D��<�+=��n=H�=lد=�=&��=Z��=���=�g�=�6�=*�f= H�<@7���y=���½>V��]X�XF���_��~ǾY�ܾ2l���j��e�پ��¾�]��󆾋zN����瀽���N�Ԃ�����;h,�<tI�<��<���<`fs<0��;�   �   ;�0�F�8���l��l񒼬f��P�W�����RȺ�a�;8N�<�w�<�<+=x�b=�Q�=ҷ�=>�=���=�+�=��=��=I��=��=�2�=Ncb=$	�<� o��P���<%<��h��4&����̾����������c���O ��/ʾ�ѥ�e���_=���=Þ�n %���c�`h4;h_8<�
[<�W3<@�; ���   �   x@���g�8�k��K��H	��]-��n�;�Q<���<@�=�0=r�^=9��=���=~�=�/�=�z�=|��=���=�.�=���=���=�y�=h��=�Z=@��<,>Ƽ���g�,[�#���MT�����P�۵� ��:#����X=�Ez��꾺B�����D�b��8�|VϽ�t�������6��畺�F; 	X:��H�����   �   �Z���_��`On����@�2� ��;���<��<H�=@.I=&�w=�=g��=c��=���=ڋ�=�A�=��=c]>�>��=H��= ��=��=X_R=��m<�4��I��	�"�Yt��˦�`oվ�m�����%�q0��3��/�̜%�Ѡ����9�־5,��T7��q�6��j��𘽤~.�������2� 9�0v��2+� �d��   �   xU��8Z��hx���� <(9�P/<���<BU=�?=�p=u��=�=ڢ�=��=��=�w�=�� >��>^�>��> l >�N�=p��=L�=�6L=��9<�E�zɽʿ.��(��oK��n��%	�܈��w/��T:�N>��L:��x/�����	�����̵������-F����硬��LO� v�䯌��6O��sR���{�0���   �   ���������J��Y'����Q�� �� $��}A<�B=�R=�Z�=�٫=p}�=c>�=��=�p>8E>��
>h@>��
>,o>l��=8��=Z��=�y�=Z-=�տ;���t㹽,�7�\�(������$?Ѿ�A�)����������k龘�Ѿ�紾�/��8{k��%2�,��G���d�� wZ���K�̗[�����j���«�c���   �   �G������]���[��B�N����XD%��k0<�K�<T�J=1!�=mb�=���=$��=���=r)�=$�>�y	>m >#�	>'�>��=q��=`,�=�C�=8�.=`=�;Fw������E;X��6���h��~;���2��^���߲�ɩ��;�����ʑ���e�.S-������`��L���)O�v�@��zP�hQt��w�������%���   �   P{��>M���L��ͧ����F����xB��;�;���<�23=\.v=���=aB�=8��=\��=���=Ř >�>)3>�>O�>hV�=r��=��=g^�=`1=�f<�I��n��ҹ�`�J�ݽ��;��)&���Y׾�徳Z��@�q�־L������񇾾U�VR��j�DL���a��9.�|� ��#0�f�R�`�~�sR���+���   �   դ������)3��`p��=�6��(*����:��<��	=�hH=h�=S��=�=:��=���=M3�=�D�=ް >�� >n��=:��=+��=¡�=��=��3=8�B<��ڼg�������6�w~q�^E��ﳮ�Z�¾��Ͼ�Ӿ/�ξ�l��2�������/q��:�.o	�w���0��L3)�������ܼ����� �aI��Ss��X���   �   �n�2Ow���p��[��d9�~[�\���`��`�;$E�<H�=�R==4�u=��=v��=(;�=���=��=���=n6�= ��=�:�=�D�=0x�=-�=�S3=�`q<�<���Xv���׽o���pQ�ƙ������
��h峾�+�� }��!Y�����I2{��IJ����!۽������.��ü��_��7��s�঺�4�� U1���U��   �   J�2�n�G�p�P�,�M��g@��U*�(��|gѼ]{���y�8<\h�<��=��R=8�=\��=Zs�=o�=^��=&+�=�j�=���=j<�=#8�=r��=ZD,=� �<��c�z�F��y�����e�.��,X�̯|�ׂ��&-��e��[ߒ�
���
p�D�H��q����z՛�b6�t$��`�w�@��;0P�; GB;`����t� �Ҽ���   �   ��������<;�$�N��Y�\\�N�U�n=F�"�,�r0�|粼 �����;���<�%=/e=#�=��="v�=���=ơ�=��=cM�=��=>gh=j�=�߀<�;#�(�hE��E�Խy���[-���I��I_�K�k�]�m���d���Q��,6�z��g���{��@�2��݉���s;p2�<�9�<��<o�<�O_<`oS;Xc�@���   �   ���d���{6�6Ac� �zE���c��l��^���������x�R1?�����P(���<H�<�<=<Tw=6X�=��=RƢ=�5�=B�=�Dy=�CB=�,�<H,E<��Ҹ�R�i�����j_ܽ
��=���(�0�0�
�/���&�j������Ľ3������<�x�.<d��<��=�4=�5=�R"=�> =�< ��; Ļ�   �   �DJ�t"����E��}���7���ɽ5��Q��Q�����Dݽ�h�����̕N�~׼ 91����<�Z=�M=zq=�`�=�|=x�f= �A=�3=���<06�;(FJ�8 ��ƸE�n{��m4��$ɽ���G��J��:��E>ݽHb����x�N�l׼�0����<6`=��M=X~q=�b�=��|=�f=8�A=x6=0��<�A�;�   �   ��Z����i�����cܽ���@�9�(��0���/���&����������Ľ���T���<�x.<H��<�=��4=�5=�N"=�: =�<���;�)Ļ������bz6�>c�|���B��X_���������|����x��&?��q��,(�@�<��<��<=6Yw=\Z�=�=Ȣ=Y7�=zC�=Gy=�EB=�/�<�-E<�   �   0D#��+�JH��<�Խ���^-��I��M_�b�k�{�m���d���Q�T06�j��j��)���:�2��鉼 ~s;X)�<�0�<���<�f�<�>_< .S;hr��F������J���<;���N��~Y�v\���U��5F��x,��'�`ղ��x��;�;Ī�<�%=�4e=��=:��=�w�=<��=3��=U��=tN�=��=^hh=Ī=�ހ<�   �   ��c�0G�?}���(�.��/X���|�ڄ��>/��g��]ᒾ����p�!�H�t�����؛��6��-����w����;�/�;�B;�8���u�,�ҼL�j�2���G�f�P�ܤM�4f@��R*����L\Ѽ�C{��4y�x;<@v�<~�=��R=�:�=���=bu�=�p�=ܞ�=n,�=�k�=w��=%=�=�8�=���=�C,=���<�   �   �C���]v��׽���}sQ�h����������g糾�-���~���Z��N���4{��KJ�����$۽򣐽��.�@#ü��_�X�7��s�Ȯ��"���X1�6�U��n��Qw�<�p��[��c9��Y�d������0D�;PO�<��=6X==:�u=P�=���=�<�=��=\��=���=e7�=���=p;�=4E�=ax�=�,�=�R3=�Wq<�   �   @�ڼ�����7�6�	�q��F�������¾M�Ͼ��Ӿ��ξ4n��h�������1q�R�:�:p	�'���"���5)�l�����ܼ������jdI�Ws��Z��C��������3��$p���=���L&�� u�:l��<*�	=�lH=K�= ��=��=���=8��=b4�=�E�=>� >� >��=���=M��=���=��=�3=0�B<�   �   M�Bq��S��5�J�ﾅ�l��q'���Z׾h���[��A�g�־�������)�|U��R��k�M��Fa�
;.�(� ��%0���R���~��S���,��c|��N��LM�������F������B�`I�;���<53=�0v=���=�C�=H��=N��=���=� >�>_3>�>h�>vV�=R��=ɖ�=�]�=F^1=�\<�   �   Pz����͖��<X��7���i��S;ǧ�������i��0��H�;�����ʑ���e�&S-������`��
L���)O��@�P{P�<Rt�Hx��@���!&��iH�����1^���[���N�p�� A%��o0<�M�<��J=�!�=
c�=F��=���=��=�)�=F�>�y	>s >(�	>�>k�=!��=�+�=�B�=l�.=�*�;�   �   ���乽�� �\�l(��Y���v?Ѿ B�I�����������j�O�Ѿ�紾z/���zk��$2�� ��F���c���uZ���K��[�>��lj���«�%��n���E����J��'���Q������!��A<�B=&R=�Z�=ګ=p}�=X>�=��=�p>"E>��
>I@>��
>o>
��=���=���=�x�=ZX-=pƿ;�   �   �w�7�����D;X��6���h��<;��侮�����"�����*�;�����ɑ��e��Q-�����_��hJ���&O��@�HxP� Ot��v��|���Y$���F�����\��tZ��P�N����@9%�@v0<�P�<��J=9"�=Zc�=���=���=8��=�)�=T�>�y	>� >:�	>2�>��=o��=P,�=lC�=�.=�:�;�   �   H��m��:����J�[������\%���X׾ ��xY꾈?��־�������������U��P��g佚I��0a�H5.�|� ��0���R�X�~�LP��})���x���J��!J��0���v�F������
B�Pb�;���<�63=D2v=T��=�C�=���=���=���=5� >�>w3>&�>��>�V�=���=���=�^�=a1=�k<�   �   (�ڼp	��O�����6��|q�MD��������¾��Ͼ+�Ӿj�ξk��z�����-q�o�:��l	��������l-)�H�����ܼ����~���[I��Ms��U����������/��"	p���=������� ��:T��<�	=�nH=�=���=C�=��=���=�4�=(F�=c� >H� >V��=��=��=���=�	�=�3=��B<�   �   �2���Rv�!�׽j��PnQ�`������=��u㳾�)���z��W������.{�cFJ�4���۽N���<�.��ü��_��7��s�X�������M1�܌U�z n��Fw���p�`[�b[9�"R�䑹� o�@e�;�U�<�=Z==��u=��=���=T=�=t��=���=��=�7�=m �="<�=$F�=�y�=�.�=xW3=�qq<�   �   Цc�\�F��u������.�v)X�(�|�Հ�� +���b��ݒ����Pp�f�H�#n����5Л�>	6�|���w���;0��;��B;0ߝ� �t��Ҽ��|2���G�vP�t�M��\@��J*���QѼ�1{�`�x�`F<lz�<�=��R=4;�="��=�u�=/q�=:��=�,�=Xl�=8��=0>�=	:�=���=I,=��<�   �   �#����@��ߊԽj��,X-���I��E_���k���m�n�d��Q��(6��������u����2��ˉ� Pt; A�<LG�<���<�|�<�l_< �S;0A�t-��������B1;�}N�NuY�R
\�$�U�:0F�0t,��#��ϲ�hp��H�;4��<�%=�5e=��=���=Zx�=���=£�= ��=�O�=:�=\lh=(�=��<�   �   ���ί�2�i�&�$Yܽ���9���(���0���/���&�9��=x����Ľ������x�<�Ȳ.< ��<̫=��4=j!5=�Y"= F =+�<@)�;@�û������\o6�4c�섽2>��\��������Rz��*�x��$?��n�@((��<h�<v�<=�Yw=�Z�=e��=�Ȣ=8�=�D�=�Iy=�IB=�9�<HIE<�   �   �#J�`��v�E��u��@.��mɽ��Ὢ��B��:|�Y6ݽ�Z������@~N�@T׼ 0�$��<fh=B�M=&�q="f�=�|=��f=f�A=P>=�Ī<0��;J��
��ʮE��v��f0���ɽ������H����� =ݽna��p��p�N�lj׼�0�З�<�`=��M=(q=hc�=�|=ҡf=ēA=�9=���< t�;�   �   ����&��0p6�.3c��ꄽ�;���X��������t����x�2?�`X��'�(�<�#�<�<=�`w=�]�=��=ˢ=[:�=�F�=�My=`MB=T@�<�SE<��������i����[ܽ��]<���(�a�0�j�/���&��������Ľם��x���<�ȑ.<���<R�=�4=�5=~T"=�@ =H!�<0�; �û�   �   ����6��3;�n}N��sY�R\�Z�U��)F��l,�h�Ľ��@K�@��;p��<x#%=�<e=.��=o �=�z�=���=��=��=VQ�=��=^oh=��=���<`#�< ��A����Խ��aZ-���I�)I_���k���m���d���Q��,6�P���ή{����2��܉���s;�3�<;�< ��<�q�<W_< �S;�U��6���   �   p�2�8�G��xP���M��\@��H*�ҵ�<HѼX{�`�x�Pb<Ȉ�<4�=��R=h>�=��=[x�=�s�=T��=�.�=n�=���=�?�=p;�=ĝ�=K,=t�<p�c�@�F� w��?��B�.��+X��|������,���d��:ߒ��	��]
p�%�H�~q�t��D՛��6��#�� �w�0��;pV�; XB;�
����t�l�Ҽ���   �   �n�|Jw���p�T[�\9��Q������c���;�^�<"�=p_==�u=u�=t �=�?�=���=���=�=R9�=��=o=�=ZG�=�z�=�/�=Y3=�uq<�2���Sv�W�׽v���oQ�l���k������<峾�+���|��Y�����12{��IJ�	���!۽w���t�.�$ü��_�x�7��s���������R1���U��   �   ����ڵ��1��8p���=���L���3�:,��<�	=rH=��=���= ��=��=*��=26�=�G�=� >�� >l��=��=��=���=�
�=n�3=8�B<��ڼ�	��*���d�6��}q�"E������3�¾y�ϾίӾ"�ξ�l��*�������/q���:� o	�W�������2)�l����ܼ�������`I� Rs��W���   �   xz��2L��YK�������F�Ƞ�� 
B�Ph�;8��<�83=`4v=z��=2E�=ا�=���=���=�� >v>�3>��>��>�W�=���=N��=�_�=zb1=Xp<8G��m��U����J�������&���Y׾�徨Z��@�k�־F���棥��񇾸U�NR��j�1L���a�H9.�$� �0#0���R���~��Q��$+���   �   �G�����P]��[��R�N�
��P:%�pv0<TQ�<H�J=�"�=�c�= �=n��=���=�*�=��>Bz	>� >}�	>w�>0�=��=�,�=D�=l�.=�F�;&v����i��;X��6���h��p;��*��Z���ܲ�ũ���;�����ʑ���e�)S-������`��L���)O�R�@�lzP�,Qt��w��z���Y%���   �   �O�^�J�s�;� 7$��T��Cɽ�$��4��� �e:l/�<�[]=�@�=�¾=��=�9�=�>|:	>��>�>g�>�	><>m�=��=ᤱ=G;�=^"= �;�����1K�p�#�p�P��+y�'���߾���@���!͌�Fz{�+�V�%
0�8�4ؽ.u���֐��K��Л�g��N齜0��U'��<���J��   �   �K�V?F�l�7�� �D��`ŽxȀ���� pH:x^�<�yY=�ϗ=��=���= c�=X�>��>��>�>��>U�>�#>�K�=��=���=5	�=\$=�q�; :�e���n�Ml �U�L�5t�/���q����떾Fm��������u� ~Q��G+���ոн�Σ�镊�� ���j��ς��U��J
��"�R�7���E��   �   Z=��9�i�+���������x����t���� �=9�9�<�$M=.6�=���=s�=��=V�=�>B�>q	>�Y>��>|��=���=��=���=�,�=2z=�\ <�׼L����׽d��iT@�01e�d���R���P��i҉��\���Sd���A��v�=����L��0s��2�p�Qh��ɂ�/w��`�˽^��������)�D�7��   �   M�'�|�$��
�E�����bͪ�f�c�x�� �̺��<ts6=���=��=���=���=���=P��=�>a>�t>v�=��=���=�c�=>N�=��q=�=�<�$��hn��Dý�m���-���N��>h��Ex�l�|���u�Pd���I��)����g�Ͻ����"d��7���/�K��
���[��Y3ֽ�T��m���!��   �   U�HN��[��R�HCƽ�ҙ�$XT�P��"��܍�<~^=F�[=��=�̫=\^�=2O�=�F�=���=�1�=���=���=�9�=���=�U�=���=|Y=�� =0&�;T���T�� ��������2��'H��U�(�W�%�P���?���'�(�
���ؽ�q����]�C�D�ܼ��μ� ���3��"{��k��&IϽ0󽓍��   �   8�Rx���ڽ�ǽc���q���"�M�.���TU�@��;�N�<^H!=��`=���=bR�=�޼=B��=���=2��=��=���=#��=@"�=�=�k{=0�4=L/�<��2;\o���m?����̽������L%�PW.�M/��L'����Z���hн�皽Z�P�����Ht���лp���C)��������p?a�xە��G��Zѽ�   �   ߲��iů�0���$��Sa������:XW�Z!��%ϼ A,��Y�;��<r=�UM=�T�=�?�=?�=~`�=��=b��=���=��=�=v�}=��B=�� =�d<�۝�x�ȼ�u7�xz��̭��oҽj��<�����P�� q���ܽ┵������V4�п���L��8 <�}<��<��A< p ;X�@�(��x�5�b�t������   �   �d��߁��\���ӎ�aߌ�>��*v���W�
G1����T�� ԑ��c4<���<��*=��`=!��=�K�=}��=C�=i|�=��=�Ih=��4=���<�9o< b��<L�������A��1{�ֶ���׭��\��q�ǽ�ǽ�2��.����㍽ԇT� l��ZU��Ħ;<��<�# =�
=Bd=��
=<��<��U<����)��p���8��   �   ��
��9��5a�W���Nl��w���g���^����(���
t��lF���Õ�����H	�<�F =B�4=PDZ=|�n=x�p=Z�`=�A=�#=�y�<�.<�ֻ�����
�"�9��7a�g���wk����׌������$���t�@dF���������ҍ�P�<hL =��4=.IZ= �n=�p= �`=�A=�(=���<0E<��ֻ�����   �   �F���l�A�D3{�����ڭ�Q`����ǽ��ǽn7������0荽|�T��s��vU�0��;�<� =�=V_=��
=H��<`�U< ̶��6�����8�Td��ၽ�^��^Ԏ�Tߌ�P����u���W� A1�>��F�� ���8~4<$��<v�*=� a=}��=�M�=���=Q�=�~�=��=BNh=��4=���<Ko<@铺�   �   `Н���ȼ�v7��{��~έ��rҽv����8�����Rv���ܽh��������]4�p̺�py���<l}<���<��A<  ;H�@���㼊�5��u�=���&���8ȯ�gï������a��P���RVW��V!�ϼ�,,����;��<�"= [M=$W�=�A�=!A�=ab�=���=$��=h��=ο�=���=�}=2�B=� =�d<�   �   ��2;Tq��p?����̽k������N%��Y.��/��O'������xlн_뚽\�P����P\t�`�л�7��pX)�ܛ�����2Fa�ߕ��K��

ѽ�;�l{�n�ڽ��ǽ����ٔ��~�M�<�� IU��Ҫ;W�<�L!=��`=���=ZT�=��=��=@��=���=��=2��=���=�#�=[�=�m{=�4=�1�<�   �     �;�W��T�5��!����T�2�S*H�\U���W���P�6�?��'���
���ؽ^t���]�DG�x�ܼ(�μ ���3��({��n���LϽ�	�W����O�H]��T콦DƽRә�VXT�l�p��蒂<la=� \=r�=vΫ=�_�=�P�=7H�=���=3�=���=Ć�=�:�=���=lV�=O��=�|Y="� =�   �   ��<�)���kn�Gýto�d�-���N��@h��Gx���|�
�u�4d�I�I�Z�)����d�ϽԶ���%d�"�7���/��K����'^���5ֽV�o�h�!���'���$���-����$Ϊ��c�����j̺L�<zu6=ʯ�=�=���=���=���=5��=n�>ha>�t>�v�=��=��=,d�=�N�=��q=N=�   �   �U <�#׼����;�׽����U@��2e�?���S��RQ��'Ӊ��]���Td�j�A��w�c����M��t��
�p�
Sh��ʂ��x��
�˽;��������)�X�7�k=��9�=�+�J�������y����t���� �>9�;�<R&M=�6�=P��=0�=���=��=>��>6q	>!Z>��>ɚ�=$��=��=���=�,�=>y=�   �   d�;�>�Θ���o�Dm �a�L�Ht������i얾�m��>����u�^~Q��G+����н�Σ����� ��ak��k������
��"���7�\�E�_K��?F�Ȭ7�J� �m��D`ŽzȀ�\��� �H:�_�<�zY=�ϗ=<�=$��=Pc�=x�>��>��>$�>��>X�>�#>wK�=��=P��=��= #=�   �   ���;x��Ï�FL���#���P�,y�O��������@��ῖ�͌��y{���V��	0��7�^ؽwt���Ր�KK���ϛ��f���M齇0��U'���<���J���O�>�J�Q�;��6$��T�DCɽ5$�������e:$0�<�[]=�@�=�¾=��=�9�=�>j:	>��>�>N�>�	>�;>�l�=D�=`��=�:�=� =�   �    s�;�9�I����m�#l ��L��t�蓉�����떾�l��k�����u��|Q�F+��
��н�̣�w���J���i������!�Ὠ
���"���7��E�K�y>F���7�%� �l���^Žǀ������
I:�b�<�{Y=XЗ=��=b��=~c�=��>��>��>2�>��>l�>�#>�K�= �=���=G	�=�$=�   �   d <�׼�����׽���dS@��/e�����Q���O���щ��[���Qd���A�&u�F���J���p����p��Lh��ǂ�"u��4�˽���g����)�̵7��=�e9���+���·��3v��t�t�h�� VB9�A�<~(M=�7�=젳=��=��=:�=#>��>Pq	><Z>Ҋ>��=���=d�=H��=�-�=�{=�   �   ��<����cn�Býyl��-���N��<h�NCx��|�y�u��d�?�I���)������Ͻ±���d�n�7�R�/��K����X��!0ֽ�R��k���!�6�'�V�$�\�*����ཀɪ�(�c����@�˺@�<xx6=�=��=���=d��=��=���=��>�a>u> w�=	�=���=�d�=�O�=��q==�   �   P�;XH��r�S�N��� ����2�@%H���T�:�W�1�P��?�3�'���
���ؽm��؀]�"<�\|ܼ@�μ8 ���3��{��g���DϽ��#�����K�^Y��M�D>ƽ�͙�OT�0�� 䴻d��<e=>\=|�=<ϫ=r`�=Q�=�H�=��=R3�=2��=.��=3;�=r��=\W�=���=f�Y=�� =�   �    �2;�`���e?��	���̽x�����	I%�(T.�/��I'�g��`���bн�⚽P�P�� ��8+t��л ۡ�`()�X�������6a��֕��B��� ѽZ2�~r���ڽ"�ǽ����ގ��n�M�����.U� ��;�^�<�O!=�`=p��=�T�=)�=R��=���=��=Z�=���=��=f$�=b�=�p{=��4=�;�<�   �    �����ȼNl7�tu���ƭ��iҽ\����i������j����ܽ܎������L4�����p
���><`�}<��< �A<�� ;(�@����ξ5���t������3���޺���x��[��K���.LW��N!��ϼ�,� ��;$�<@%=�\M=�W�=XB�=�A�=�b�=8��=���=܄�=l��=���=6�}=�B=�� =!d<�   �   �9���v�>�A��&{�����ѭ��V��
�ǽ��ǽ,��Ȋ��eݍ�J|T�ja�p3U�p�;H�< + =�=*k=�= ��<�V<�괺X����P8��d�Rف�nV���̎��،�����u�ĔW��:1�<��>�������4<|��<��*=�a=⣆=/N�=�=��=�~�=_�=�Oh=��4=���<�Yo<�L���   �   ��
���9��,a�����e���퓽�����}�������s�FXF�,���������`(�<�T =�4=PZ=��n=��p=��`=�%A=l0=`��<�i<@pֻ�����
���9��(a��~��te���q���z���"��H�s��`F��������@�����<LM =H�4=�IZ=֫n=гp=��`=�A=:*=X��<@O<�ֻ�����   �   �d�k܁��X���Ύ��ٌ�����u�"�W��51��1���J����4<Ȥ�<��*=a=ܦ�=�P�=���=N�=���=�=FUh=T�4=��<�po< ���H0��"s�ƏA�&{�����ӭ�!Y��Y�ǽ��ǽ�0������i⍽$�T��j�xVU�@˦;���<j$ =p=�d=��
=��<��U<@ϵ�(%��|���8��   �   ǰ���¯�ڽ��{��v\�������KW�dL!��ϼp,��К;��<2+=�bM=�Z�=E�=D�=(e�=~��=γ�=��=�«=��=�}=��B=�� =H2d<�}����ȼ�j7��u���ǭ��kҽG������������o��&�ܽ-�������U4����� H��h"<�}<��<`�A<`} ;@�@���㼴�5���t�!����   �   `6�9v�8�ڽ��ǽ���������M�8��@&U���;�f�<T!=�a=ß�=AW�=R�=d��=���=���=8�=���=��=X&�=`�=�t{=��4=�B�<@ 3;]���d?�
��Q̽�����
K%��V.��/�xL'�4����hн�皽��P� ��Gt�0�л����A)�t������l>a��ڕ�G��ѽ�   �   ��~M��Z�fP�V@ƽ;ϙ�~PT�����۴�<��<�g=Z\=.��=�Ы=,b�=�R�=5J�=���=�4�=���=���=�<�=��=�X�=%��=f�Y=H� =p`�;�E��N�S�����a����,�2�%'H�3U���W�ѦP���?�˶'��
�y�ؽ�q��$�]��B���ܼ�μ �
�3�F"{�2k���HϽ~����   �   ߥ'���$��	�f������ʪ��c�l�� �˺<�<z6=���="�=� �=���=P��=���=$�>b>�u>Hx�=3�=��=2f�=�P�=�q=$=�<���`cn��Bým�̦-� �N� >h�6Ex�"�|���u�(d���I�ڟ)����:�Ͻ����D"d���7�p�/��K��
���[��3ֽtT�Mm���!��   �   =��9���+���\���mw���t�(�� "B9lB�<Z)M=S8�=���=p�=���=�=�> �>�q	>�Z>9�>���=|��=T�=>��=�.�=�}=j <�׼Ƚ����׽����S@��0e�?���R��kP��[҉��\���Sd�v�A��v�'����L��s���p��Ph��ɂ�w��=�˽6��������)��7��   �   �K�0?F�2�7��� ���]_Ž�ǀ�4��� �H:�b�<�{Y=�З=��=���=�c�=ç>�>�>p�>�>��>	$>QL�=� �=q��=
�=&=��;�6鼦���_m�l ��L� t����b����떾?m�����u�~Q��G+���ŸнtΣ�ݕ��� ���j��Â��B��@
�p�"�@�7���E��   �   ������1��ҕ��I}��fI�j���{���}B��"λ��<Οo=�ڨ=ӝ�=~-�=N>Ju>nz>��>�|>��>$�>��=���=�=�ߡ=N�u=$b=`#V<�i��T1������ν�� �x��Y�!�}�%�y�!�H��xs�Ƨ� ^���v��>���������>½�����@'�[T�O:���Ж�0n�������   �   32���D������CÒ�Zx��CE�B���$���=��C��\��<Xnn=9��=�=n_�=�T >�o>Df>_�>75>�v>nS>�{�=XB�=0ÿ=�Ǟ=;p=�L=��L<Vj�,�.��i��M�ʽbR��W��B����!��~������ ��Qٽ�����"��A���p�4���6������H�"�p�N��Z|��l��Ť�%,���   �   ������˚�����Di�Me9����ٯ��+.�P큻���< Lj=��=~5�=���=��=�I>A>3�>vR>�7>q�=*��=b�=���=�8�=�p_=�3
=��,<��p��)�J��MN��6�콢�1��5#��g�:���9꽈Ľڞ������]�t�[�(��\¦�H��T*��3?��j�t���$)��'���   �   �������V~����x�h�R��b'��&��~ǝ�2)� ����<��a=���=H��=p!�=bQ�=���=�M>+�>�� >���=L��=
��=��=��=�i�=�MA=��<�*�;����$#�����]ڮ���սB��y��0�������T�ƽǢ�j����G�Zv&��>$���E������!��� ���&�O���t�﬉����   �   �V���H����p��W���6����_�ս8L��������d�<XpQ=��=�I�=���=H�=���=���=���=)�=��=~�=���=��=� �=�AV=8�=���<�r	��ƣ�v�"��eq�pל�z@��Pѽ��ܽF<ܽ��Ͻݕ��r6���Qq��B1��m��4���l���P\���<;�ʔ����ʽh*��2,���M�D�i���|��   �   ��T���R�^VG�G^3�@������ϵ���l��>缀���־<�7=�"�=e��=F��=S�=yJ�=[��=�G�=X��=�l�=,�=��=z�=Z�L=��=���< �};�C�T��.��(h�8Y��@R��%��e7��B����:��������P����@���%��
^��y4�������� 1��ꍽ��ʽ���\�"��v;�7�L��   �   ��$�T%�����������)u˽yK��^�P���޼`=��p��<�n=�ET=m��=a�=���=�^�=г�=eݾ=�	�=���=�Վ=�h=".=�`�<HdH<���������\p$�&�L�L�n��I��dO��v���׉�F�{���U�7$��RּLB����:xX=<@��<$�<��V<�7�:�v���e��=���j��U��[�����   �   m��#����"B߽2ǽ�٨�伆��?E��_��P�J����;�]�<=R�P=��=��=��=��=�=JC�=�uv=��A=�=���< }V��j��Ě���E/���U���q�󒁽�}���ф��Q�>�k���N�>�(�X�򼸐�� ���9<X��<�2=�d=h"=f=�T�<��7<p�����PsR�	�������F�ڽ�   �   5���ب�39��Y橽���7���X#{���M��p���ȼ�t(�p��;@�<�=>5=�Y=�p=(Bu=Vh=�>H=�=/�<�a;�w���]�$iS�@����	���ܨ��<���詽f
������$#{���M��m���ȼXb(�൐;(�<x=�5=��Y=dp=�Fu=Ph=XDH=�==�<��a;�f���T��_S������   �   �>/���U���q�@���#}���ф��S�n�k�6�N�X�(�X������3�@�8<��<�-=`="c"=�=,I�<��7<P���P���|R�:���򌼽ÓڽWr��(��O�E߽�ǽrۨ����P?E�\���{J���;�e�<4=x�P=��=��=��=!��=L�=�E�=l{v=��A=�=P��< �T�,[��P����   �   T��� �:m$�x�L�B�n�JJ���P��<x���ډ�0�{���U�<=$��^ּ�bB� �:pD=<l��<���<��V<�u�:�����m��B��p�����L�����$�%�F�������Jw˽�L���P���޼p/�����<�q=�HT="��=�=���=^`�=���=P߾=��=�=؎=��h=.=�l�< }H<����   �    ,~;H�B�Q���.�2*h��Z��:T���'��N:��d����=��!�����P����'����%� V^�@�4�H��L����1��W�ʽv��-�"��y;�G�L���T�j�R��XG�n`3���-����ѵ�$�l�D?� Ƌ�Pپ<7=�#�=���=���=vT�=�K�=ґ�=I�=��=�n�=-�=��=X|�=�L= �=��<�   �   ���< 	�(ƣ�`�"�hq�#ٜ��B���Rѽ��ܽR?ܽ��ϽΘ��"9���Vq�(G1�Pv����������e��B;�ޗ����ʽ�,�N5,�f�M��i�l�|�EX��*J���p��W���6�Ң��ս4M��j���z��e�<�qQ=���=�J�=��=Z�=���=���=��=Z*�=W�=��=���=4�=#"�=�DV=��=�   �   ���<,�;�����#�歁�"ܮ���ս���Vz�2������潍�ƽ�Ȣ����:�G��y&�FB$��F�!���H$��F! �F�&�O�ݖt� ������Lᗾ����_��|�x�ڕR��c'�;(��nȝ�*������<��a=���=���=*"�="R�=C��=8N>��>� >���=Q��="��=��=��=�j�=:OA=�   �   �3
=��,<��p��)�]K���O���콤�8 �8$��h���/;��Ľ$۞������]���[�R)���æ���j+�05?���j�F���*��	�����쇥�k̚������Ei�f9�;���ٯ�.,.� ���<�Lj=f�=�5�=p��=���= J>~>p�>�R>�7>�q�=���=��=��=9�=q_=�   �   .L=�L<�[j���.��j����ʽ�S���������!����E� �?Rٽ蔲��"������&������6��d���֟"��N��[|��l���Ť��,���2��,E�������Ò��x�3DE�v��	%���=��B�����<�nn=r��=H�=�_�=�T >�o>Xf>r�>R5>�v>�S>�{�=|B�=7ÿ=�Ǟ=�:p=�   �   �`=�V<ثi�V1����b�νB� ����|�!���%�j�!�#��<s�9��n]��Wv��±������p���=½�����@'�XT�O:���Ж�/n��������������0���ѕ�VI}�NfI�:��U{��F}B� λ���<�o=�ڨ=ݝ�=|-�= N><u>`z>��>�|>g�>�>���=���=��=(ߡ=D�u=�   �   ~M=x�L<PSj�f�.�;i����ʽ�Q���������!��}�̴�8� �NPٽ���2!���������4��M�����"���N�+Z|�l���Ĥ��+���1��1D��
�����Kx��BE�c��N#��=��1��4��<�on=㮧=��=�_�=�T >�o>hf>��>[5>w>�S>*|�=�B�=�ÿ=VȞ=�;p=�   �   J6
=x�,<��p�� )�pH���L��C�콎����!��f����,7�Ľ�מ�����]���[�)&��W�����")��2?���j�����6(��'��������ʚ�􉾮Bi��c9�2��m֯��&.��́����<Oj=?�=�6�=���=߱�="J>�>��>�R>�7>�q�=��=c�=���=�9�=�r_=�   �   Ę�<�O�;̵���#�ߩ��z׮���ս���Rw�/�����*����ƽ�â�j��Z�G�q&��9$���E�E������ ���&��O�G�t������񓾩ޗ�����|�� �x��R�G`'��"���Ý��"��=����<��a=���=׎�=�"�=�R�=���=cN>��>8� >��=���=���=���=b�=�k�=�QA=�   �   H�< ��丣�N�"�^^q��Ӝ�r<���Kѽs�ܽ�7ܽT�Ͻ����q2��DJq��;1��`��𒾼l�(P��D6;�:����ʽ&(�^0,���M�,�i�;�|�!U��G��5�p���W���6�Ğ�Z�ս�G��������8p�<�uQ=p��=�K�=ˣ�=��=��=��=l��=�*�=��=i�=��=��=#�=>GV=4�=�   �   �t~;8�B��B�$z.��h��T��rM��/ ���2��f����5��n���H�P�v��4����%� �]��4��o�\��R1�I捽�ʽ��E�"�}s;���L�$�T���R��RG��Z3���o���;ʵ�>yl�\,缀ي���<\7=w%�=☠=���=U�=\L�=@��=�I�=^��=�n�=��=o�=}�=�L=Ī=��<�   �    ���L��e$���L���n�5D��J���p���҉��{���U��-$��@ּ�*B� ��:Xu=< ʐ<��< W<�!�:�f���\��8��8e��������e��&~$�m%� ���������|n˽ME��
�P�@�޼P��< v=LT=T=��=C��=�`�=
��=�߾='�=S��=�؎=��h=�.=�p�<��H< g��   �   v:/��U���q����x���˄��F�,�k�8�N��z(�����}���N�`$9<l��<�9=�k=�n"=0
=lc�<X�7<�m��4��$hR�ۜ�������ڽ�e�;��j�:߽�ǽӨ�r����3E��I�� _J�P٤;�m�<V"=ƿP=��=p�=�=���=��=F�=,|v=��A=�=D��<�T�V�������   �   8��S֨�6���⩽)���ڐ�~{���M�c�X�ȼ0<(����;�8�< !=5=T�Y=�p=Mu=�!h=:KH=4"=�M�<�b;�Q��
I��RS���������Ѩ��1��ߩ����_ِ�J{�H�M�>e�X�ȼN(�0Ԑ;�-�<�=�5=��Y=Dp=�Gu=h=
EH=p=�>�< �a;d���R�F]S� ����   �   Sk�!��a���>߽?ǽZը������4E��G���UJ���;�u�<�&=p�P=�=��=��= ��=B�=�H�=>�v=@�A= =0ˁ<��Q�LD���r���1/�8�U���q�k���^v���ʄ��F��k���N��(���� ������ 9<��<�3=�e=�h"==(V�<P�7<����D��4rR�O���������ڽ�   �   N�$�r%����\������_q˽.G���P�Я޼�ꙻT�<y=�OT=5ć=��=H��=�b�=%��=��=��=�¤=hێ=��h=b&.=H�<0�H<���P�������`$���L���n�D���J��Cr���ԉ���{���U�T4$��Nּ(FB� Ӣ:�[=<���<L�<��V< H�:�u��Xe��=��j������������   �   Z�T���R��UG�4]3��������̵�|l��.��Պ��<R
7=�&�=T��=��=�V�=N�=���=XK�=b��=q�=�=��=��=�M=��=���< �~;`�B�,;ἶw.��h��T���N��"���4��]���:9��򣅽X�P�l�����(�%� ^�@r4���������1�^ꍽ��ʽ���$�"��v;���L��   �   �V���H����p�#�W���6�j��͓ս\I��������q�<�vQ=F=�L�=���=,�=e��=~��=���=D,�=g �=E�="��=�=V%�=�KV=��=��<���������"�^q�Ԝ��=���Mѽ��ܽ�:ܽ��Ͻ����5���Pq��A1��l��x��������[��f<;�����ήʽM*��2,���M��i�@�|��   �   �ߗ�a���~��(�x���R��a'��$��nŝ��$��[��p�<~�a=?��=���=�#�=~S�=���=�N>D�>Ϯ >f��=��=��=T��= �=�m�=BUA=��<�d�;䱄��#�Щ���׮���ս���bx�C0�]�������ƽ�Ƣ������G�v&��>$���E�ܮ���!��� �l�&��O���t�ݬ�����   �   �� ����˚���Di��d9����ׯ��(.��Ձ���<2Oj=��=�6�=h��=n��=rJ>�>��>8S>m8>�r�=/��=� �=۪�=;�=du_=�8
=��,<@�p���(�IH���L����� �����"��g���z9�SĽ�ٞ�����^�]�<�[�(��I¦�3��J*��3?��j�m���)�����   �   +2���D������/Ò�&x��CE����3$��^=�8��\��<�on=���=��=$`�=U >�o>�f>��>�5>Jw>�S>�|�=qC�=MĿ=.ɞ=|=p=2O=�L<hMj�2�.��h����ʽ�Q������b�!�s~�v��� ��Qٽ�����"��2���\�$���6��u���B�"�i�N��Z|�l��Ť�,���   �   �D��A�7������qѾM������P�;���b�j����D�=��=��=B��=��=��>6�	>[&>��	>>n0 >c��=:��=��=�?�=a�=�se=��!=��<��v;�@i�0���
K;��qi���>���-���n��!P��2��"���(��P�y���:=ӽ*.���P���������"Ӿ�l��.���A��   �   i�Kw����ﾯR;���������7�a�罰�b� �ٻjG=h2�=nt�=���=j?�=8!>P�>�	>^4>:6>�H�=]�=9 �=�|�=�=�ߌ=�,\=��= �<@&4;HKp��L���8�X�c�*�~��N���|���d�\�E� �(�6��� �<�E��e����˽��yK�l݆�UǪ���ξ@w�:��fo��   �    ��a����Qᾪm���Ý�<Cr���+�o�ֽ\eL�@�]���=4��=j�=���=���=�l>[[>��>H�>���=.��=��=V�=̲=`$�=@�z=*y?=�� = �~<�R�����.��4�/�0�T�j�ʡm���`��hG��	(���<���x~���%��qr�ַ����<�N{�7���W���
�6,���?��   �   B{��`��	㾫̾F��؎���4Z����CC��>�*�@˩:�=i��=W��=Z/�=�W�=V�=�E�=�/�=:�=��=���=s�=B}�=̗= 0{=�D=j�=�F�< W�;P�� ���M��f�%���?��K��[H��6�V���Q��8ﹼ�ȗ�����"伴Q9��o��6>�,�#�	�]��r��H󭾤�ʾ���Q��   �   ��վ�ҾFyž텱��+���]w�X�<����6���	�0c�;2�=���=�۬=@A�=c��=~D�=�=l��=�B�=|��=f��=�=aW�=B�`=r�)=���<j�<�t|;��� ���?ؼ�
���ο*���)�Ɨ�N�|lǼ���`F����������pB� 4�n�U�h��".��
9�X2q�׵���d���'þ�о�   �   *���"ٮ����������}�<N��~�U^ؽ̒}�,���P:0<j�=��}=���=>[�=���=cF�=HX�=��=��=���=$M�=
�o=��2=0{�<��l< �:��&��̢�0�⼜�	�rk�<Q#�:$��(�j� �� ڝ��"� ��Г�;`�G<(�J<�_�; d�L��:o���Ľ�X�w�?���p���������٬��   �   _���,ߊ�/��b�l� =K�%�:�������C�(�y�P�Y<��=��k=�ݕ=��=+�=�(�=h�=t1�=�<�=���=�DC=(&�<P6M<���x���7�d&7���T�T�d�x�h���a� �Q�<o9�<z�T�����pg�p��;�rr< ��<�j�<���<��<��q<��Y�K�L�w��ǽ&����5��[���z��߇��   �   T�Q�:Q��	G���4�t�%���(½�-�����*�p[V<
h	=X�O=QQ�=]ǖ=l��=��=+��=}x�=�^=>�=���<�ku�|jҼ�|>����6㡽򩵽���c��ˬ��B���yԌ�r�d�>�*���ܼHE�@50;X�<0Y�<�h=�l:=��C=�P8=�=4ֱ<�mx:`ϼ8�d�?������X^�h6���H��   �   >��@��R���P��.潣����N�O�p��P���<��<FQ(=�W=��w=䐃=Ca�=�Qi=fL:=,��<��;�9��fZ3������Ľ؆��x�������~���S��2����R!����O� �H���<���<T(=�W=�w=Ԓ�=rc�=�Vi=<R:=��< Z�;�&��FO3�����Ľ}�.u��   �   ң��a���^��~���凣�Ҍ���d��*� �ܼ E��0;��<�R�<e=�h:=��C=2L8=L=�ɱ<��v:rϼ��d�k�����:b�@l6��H���Q�&>Q�NG��4��B���½�/��
�p�*�0^V<�i	=n�O=�R�=�Ȗ=��=��=c��={�=�!^=p�=@��<��t��TҼ�p>��|���ܡ��   �   �7���T���d�$�h���a�"�Q��m9�hz���꼌����~�0i�;Hdr<H��<pb�<���<��<��q<�ZZ��Z꼤�w���ǽl�� 6�(�[���z�M⇾����`ኾ"1���l��?K�l%�}=��_����C�X�y� �Y<��=�k=�ޕ=��=��=f*�=�i�=�3�=?�=���=�KC=6�<�YM<�ӟ�� ��~-��   �   �&�쿢�<��\�	��h��O#�2$��)�����Ἰ���h"� �� u�;P�G<p�J<p:�;�������o��Ľ�[�� @���p�����ֿ��[۬�����^ۮ���������}��N�����`ؽ6�}�ح���70<��=��}=X��=0\�=��=�G�=�Y�=���=�	�=%��=�O�=X�o=��2=��<h�l< �:�   �   4t�<�|;@ �����<ؼ�
�����*� �)�̚���|sǼ���hT�`Ɔ��Ɨ���B��=�*�U��k��G0�49�m5q������f��*þ@�о(־Ҿ6{ž����2-��D`w�$�<�ܦ�򑞽��[�;*�=׮�=Vܬ=�A�=>��=zE�=��=ɛ�=�D�=^��=���=m�=�Y�=��`=*=���<�   �   ��=`L�< g�;���x���8N��ȫ%���?���K��^H��6�X���W������TΗ����x)伢U9�r��#A���#�@�]��s������O�ʾ���,�}��&��@�̾~��Տ��O6Z�ͳ��D���*����:أ=���=���=�/�=zX�=�V�=�F�=�0�=c �=�=T��=�=�=�͗=�3{=��D=�   �   �z?=� = �~< D���� 1����/��T�4j� �m���`�kG��(������l���
%�ftr�����&��<��{�/���r���Dᾅ-��o@�� ��b�E���Rᾇn���ĝ�KDr���+�w�ֽ�fL� �]�p�=H��=��=!��=>��="m>�[>��>��>^��=��=��=k�= Ͳ=t%�=L�z=�   �   -\=��=��< 4;�Np� O��28���c���~��O��:�|���d�0�E���(�����!�2�E�]f��b�˽����yK��݆��Ǫ�3�ξ�wﾔ���o�oi��w�X��d	�S;�������7�7�����b���ٻ�G=�2�=�t�=���=�?�=P!>h�>0�	>�4>c6>%I�=q]�=� �=$}�=u�=��=�   �   �re=��!=졳<@�v;�Di�D����K;�^ri�X��R���-����n�2!P�t�2�
"��(���P�U���,=ӽ*.���P���������"Ӿ�l��1���A��D��A�,��|��qѾ+�������;������j������=��=��=G��=��=��>2�	>P&>r�	>	>V0 >3��= ��=Ǡ�=C?�=�=�   �   �-\=��=`�<�94;pFp�hJ���8���c�~�~��M���|���d�@�E�̻(�����>�E��d��~�˽t��dxK�݆��ƪ��ξ�v����o��h��v����&��Q;���6�����7�����b� oٻ(I=3�= u�=���=�?�=h!>{�>>�	>�4>q6><I�=�]�=� �=\}�=��=^��=�   �   �|?=>� =�~< s�����(����/���T�bj� �m�ҽ`�.eG��(�h�D����w��n%�*nr����N<��{�T���L������*��?�Z�<a������O�ql����ZAr�P�+���ֽ�`L��e]���=o��=v�=���=���=Im>�[>��>��>���=L��=+��=��=�Ͳ=�%�=��z=�   �   �=dR�<��;p�⻸����A����%�B�?���K�~VH���6�2��H���幼T���������L9�m��(;�`�#���]�bq�����ʾ��d�Dy��b����̾���^���:2Z�����?��*�*��k�:>�=*��=د�=�0�=Y�=(W�=�F�=�0�=� �=L�=���=p�=|�=zΗ=H5{=Z�D=�   �   �y�< �|;`�����0ؼ<
����|�*�x�)�������_Ǽ����/��}���}��H[B��(�
�U�Xd���+�
9�X/q�����b���%þ��о��վ�Ҿ�vžƃ���)��iZw�I�<���̋�������;z�=̰�=�ݬ=�B�=���=F�=X��="��=�D�=���=߇�=��=Z�=�`=�*=��<�   �   Л&�4���|��r�	��a��G#�$����D��˝���!� $�`��;H�G<��J<0��;P1�0��o��Ľ,V�+�?��p�f���>����֬������֮�!���l����}�cN�M{�yXؽڈ}�@��� W0<��=�}=䉣=P]�=���=HH�=LZ�=��=
�=z��=JP�=2�o=��2=Ќ�<��l< R�:�   �   �7���T���d�.�h���a���Q��d9�Vp���꼴����&�P��;��r<(��<w�<Ե�<$�<(r<�~Y�D:�z�w�)�ǽ�����5���[�Ȝz�w݇�ǃ���܊��,����l��8K�%��2��ғ��P�C�Xfy� �Y<��=��k=.��=��=h�=�*�=fj�=4�=v?�==�LC=�7�<^M<pȟ�����"+��   �   ^������9\����������8Ό�ҋd���*���ܼ�D�@�0;��<0g�<:o=�r:=��C=W8=,%=��< z:�Lϼ�d����9���2Z��c6���H�\�Q�5Q��G��4�"�?���½�'�����*��|V<^o	=��O=+T�=�ɖ=鉡=.	�=���=r{�=p"^=�=���<��t��RҼ�o>�|���ۡ��   �   ���p��K���O��+� ��!����O����Х��.<|��<�Z(=\�W=x=���=`f�=�\i=Y:=���<��;���LC3�� ��h�Ľ(w��p�������Σ��L�v&����7����O�t��8���)<$��<�W(=�W=x=���=�c�=nWi=�R:=<��<�^�;d%���N3���x�Ľ�~�t��   �   ��Q�l9Q��G���4�'�����
½**�������*��}V<�p	=��O=�U�=�˖=ˋ�=M�=;��=2~�=�(^=��=�ɑ<�&t��<Ҽfc>��u��ա�����-��kV������i���ˌ���d�<�*���ܼ��D���0;��<`�<&k=rn:=&�C=�Q8=d=|ױ< �x:_ϼ��d����F���^��g6�S�H��   �   +����ފ��.����l��;K��%�*7��ږ��:�C��ny�p�Y<0�=�k=9�=g��=��=�,�=pl�=d6�=6B�=��= TC=|H�<X�M<`w��p穼  ��7�|�T�h�d�H�h�~�a�x�Q�b9�bo����X����=컀��;�~r< ��<�m�<���<D
�<p�q<@�Y�0J�Ԩw���ǽ����5�ҷ[�J�z��߇��   �   ����خ�Z���p���}�DN��}��[ؽj�}������Q0<n�=��}=���=R^�="��=�I�=�[�=���=R�=��=KS�=�o=R�2=(��<��l< h�:�y&�(���4�⼂�	�
]��D#��$���f��ἴѝ�p"��9�0��;�G<��J<�d�;�_�x���o���Ľ�X�[�?���p�x��������ج��   �   ��վ�Ҿyž����q+��6]w���<����*��������;ڄ=갃=2ެ=�C�=���=&G�=���=���=�F�=���=<��=~�=t]�=Z�`=T*=l��<솁<`V};���H���)ؼP
����*�2�)���� ��gǼD
��PA���������oB�03��U��g��.��
9�G2q�͵���d���'þ��о�   �   1{��I��	㾂̾������24Z����A���*��3�:j�=#��=��=1�=�Y�=�W�=�G�=�1�=�!�=��=`��=s�=���=�З=0:{=F�D=��=L[�<��;p��8���D?����%��?�8�K��XH�̴6�����O����4Ǘ����"�jQ9��o��>� �#���]��r��A󭾝�ʾ���G��   �    ��a�	����Pᾌm���Ý��Br���+���ֽ`cL��~]���=N��=��=���=	��=�m>\>P�>,�>���=���=���=7�='ϲ=�'�=��z=�?=X� = �~<�������&��l�/��T��j��m�(�`��gG��(�p�P����}���%�tqr�ķ����<�H{�3���S����0,���?��   �   i�Hw����ﾟR;����������7���罺�b��wٻ|H=�2�=�t�=��=�?�=�!>��>t�	>�4>�6>�I�=Y^�=��=M~�=��=a�=0\=��=�<`S4;HAp��H��8���c���~�sN��f�|�4�d� �E���(����� ��E��e��|�˽��yK�i݆�QǪ���ξ>w�:��eo��   �   ��[���W��HK�J8��������Ѿ�O���9U�
��=l��P/��.%=�i�=�P�=�K�=z��=��>i>��>f� >���=��=r��=)��=�1�=�'�=2��=�EX=�-= �=47�<�;^<�n�; ��:���`b+���� E4�� *� �z� }O��=���Pm���˽	 ���j��T��j]վn���^ �gP8�dZK���W��   �   ��W�ˬS��G�^�4�޾�����̾<���hP��6��~�b�@���ZT(=.��=��=�S�=�L�=f�>��>��>X��=C��=�k�=��=�L�=j��=7��=:�t=BWJ=~� =���<��<H�G<�;�; ��:�k�� +󺀀F��=:�ʀ:`���(.�����a�U�ĽO���d�c���@�о'�0C���4�ƐG�t�S��   �   �%L��:H��<���*�5��:������xŎ���B��y罀iH�`5;�	1=�U�=��=�4�=,�=���=93 >��=X��=P1�=���=׃�=��=%s�=�1p=��F=v�=��<��<(�e<�(�;@�H; T(9 �B� T9@�;0�;���;�"T;@�������@.@��ů��^�h1T�f4����þ'����=��*��<�hH��   �   ��9�1\6�B�+��b�j���n޾�v��9i��*/-��Eɽ�, �x+<�d==�ɘ=���=�h�=�%�=5��=��={�=���=�u�=�%�=�B�=$z=��J==���<�V�<�[<��;�s9; ������ � @���3=;���;x�-<ВO<�o9<��; "��s��)�����$:��Ճ�Qů�hf޾�-�}���h+��6��   �   J�"���x�����뾓����S��p]�
��X����޼�<�<�J=nP�=��=�O�=���=`��=W��=kP�=��=���=��~=8D=D�
=�B�<��< �9��׻p39�(~c���m���Z�0$.��Ի����01�;�I?<�<ȡ�<t �<x��<�ty;�� K�_@��.�J)^�8��ÿ�ɽ�.��ҥ�RD��   �   ����?������X��ž�jp{���5����x��lo���<�U=�ȗ=聶= S�=�S�=��=�f�=�	�=� �=�L=�/=�i< �;�@����b��ZZ ��V5�Jy;��4� K!��{��Ƽ@gp��{����;H߀<�T�<�L�<H�=���<$��<��:Xؼ~����'罌P/�=�r��K�����'�ྵN�����   �   A�۾��׾Ŕ˾ϫ��8������ƣG����V���*� �8���<~�[=`%�=IM�=<��=iö=!C�=]Z�=T�l=�#=hU�<����<��|�M��R��nĨ��h��Ў��_����ά���d�s��4��b㼘�=��~;�%�<4��<�:=t21= �.=v�=��< ���s
�Ø�?
��T&7�0s��;�����թǾ�վ�   �   iŧ����R9������}r�4�E�`����ҽX|��ʼ��;�6=�AZ=3��=U �=P%�= �=�=�ZO=���<���;�&����V����<-߽²��R�7 ��� �����������½.^��V&?������fغPt�<�E	=6�:=��Y=��b=>XR=��%=T{�< �j�$��m������+�-��^������������   �   �iq�y�o�S�b�M�O0��"��Lؽ���(�#��+7��@c<&�=j_O=
�{=���=���=��p=��8=��<@QǺҮ�>�l�۽#m��7�P;T��h�
oq�Ԍo�D�b�lM��R0��%��Qؽ�����#��67�X<c<B�=f`O=�{=P��=���=H�p=r�8=x�<@4ƺأ��퍽��۽�h��{7��5T�dh��   �   m2 �r� ������vy��½yZ��,!?� ���@2غu�<�D	=��:=B�Y=�b=TTR=��%=�n�< Hk����s��������-��$^�d������6����ȧ����"<�������r���E�����ҽ |�&ʼ���;>6=�AZ=⠊=r�=�&�=�=v��=aO=
�<�س;���^wV�ߧ���$߽@��N��   �   a������ߑ��?ɬ�[���s��4��[�p�=��~;$%�<���<�8=�/1=Ό.=X�=x�<`\ �&{
�7Ș����6*7��4s�<>������Ǿk�վ��۾� ؾЗ˾����n:������ͦG��%Z���*��"9�Ȕ�<~�[=�%�=*N�=z��=Ŷ=?E�=]�=�l=�+=dh�<�4��@����M�|K��Ｈ��   �   �N �(L5�zo;�:4�D!��v��ƼH^p�0t����;\݀<0Q�<4H�<�=؇�<x�< G�:$ؼ���,罻S/�"�r��M������*���Q�����K��tA�����}[�8ž�s{�I�5�ު뽌x��wo���<��U=�ȗ=���=�S�=NU�=ʡ�=�h�=.�=�#�=��L=�8=P�i< ;������K���   �    4�9�Q׻H9�0fc��}m��Z�(.�0�Ի�����+�;�D?<l�<t��<@��<D��<�8y;����zK�D����D,^��9��3ſ�P�辕��U���E�޿"�s��ny������f���6U���]��������޼:�<x�J=�P�=U�=vP�=���=���=���=xR�= �=鎛=��~=�D=P�
=�S�<X�<�   �   ��<a�<��[<�.�;`�9; �������z� p���%=;���;�y-<�O<g9< ֓;p&"��w�:,��٣�&:��փ��Ư�Fh޾�.����j+�+6�4�9�y]6�r�+��c�V��Vp޾x��"j��~0-��GɽL/ �H&<hd==�ɘ=���=i�=p&�=$��=3��=�|�=���=�w�=(�=?E�=�z=��J==�   �   ��F=��=8��<��< �e<�/�; �H; ((9 �B� FS9@�;��;���;�
T;����@��� 1@�oǯ�$`��2T�Y5����þ�����>��*�ݒ<�^H�x&L��;H���<�V�*����;�����Ǝ�ڇB��z�kH� �4;Z	1=�U�=��=L5�=�,�=>��=�3 >��=s��=�2�=��=x��=~!�=�t�=�5p=�   �   ��t=dXJ=^� =���<t�<`�G<:�;@��:�|��@=� �F���<: ��:@���+.��t�a�N�Ľ�����d�����о���C�J�4�E�G���S�
�W�A�S���G���4�,��P����̾���hP�7���b�����TT(=@��=��=�S�=�L�=��>��>6�>ؐ�=؀�=Sl�=Z�=8M�=(��=�=�   �   俁=NEX=�-=`�=�5�<�8^<�i�;���: �� f+�����>4��*���z�@|O�L=���Pm���˽"	 ��j��T���]վ}���^ �pP8�jZK� �W���[���W��HK�98�t������ѾlO���9U��	�=l��H/�(/%=j�=�P�=�K�=r��=��>i>��>\� >���=҉�=J��=���=K1�=@'�=�   �   .�t=$YJ=R� =��< �<��G< H�; ΀:�;����� F� y=:���:���8".����h�a�t�Ľ̂�f�d������о���B�g�4�P�G���S��W�@�S���G�ۥ4�g�������̾����gP�5����b��T���U(=���=D�=7T�=2M�=��>��>C�>��=��=jl�=s�=cM�=V��=/��=�   �   �F=
�=Я�<X�<�f<�G�;�I; �+9 �A� HW9��; *�;0��;�OT;�o��(�0+@��ï��]�0T��3����þ����-=�Q�*�
�<�tH��$L��9H��<���*�b�r9��l���oĎ�F�B��v�@eH��85;l1=W�=��=�5�=�,�=���=�3 >��=���=�2�=0��=���=�!�=Gu�=t6p=�   �   (��<e�<��[<�F�;��9; ��� A��(� ��� ~=;P��;ؐ-<x�O<9<0	�;@
"��o�D'�����":��ԃ��ï��d޾�,�\���g+��6���9��Z6���+��a�M���l޾&u���g���,-�0Bɽ@' ��=<�h==7˘=��=�i�=�&�=���=���=�|�=���=#x�=L(�=�E�=�z=��J=@=�   �    $�9�>׻X9��Wc�hlm��Z�.��iԻ@쐺pa�;`?<P�<���<�	�<Ȝ�<��y;䏼��J��<���	�|&^�W6������e�����U���B���"�M��rv� ����D����Q��&]�`������޼@H�<��J=dR�=��=`Q�=���=,��=Z��=�R�=d�=+��=8�~=Z D=(�
=�U�< �<�   �   �L ��I5�Dl;�R4�l?!�,q�|Ƽ�Cp�<��p<�;\�<t`�<�W�<��=���<슞<���:�	ؼj����"�zM/���r�\I��k���4��{K��N��ׯ�>�R����U�ž�꡾$l{�^�5����jx��Mo��#�<^�U=�ʗ=���=U�=V�=L��=:i�=��=,$�=@�L=$9=0�i<`�:�$���pH���   �   `��t���E���PǬ�����s�t4�N���=���~;x4�<8��<�@=81=��.= �=��<@���j
�𽘽����"7��+s��8�������Ǿ��վ��۾�׾^�˾����65��&���h�G���P��v*��u8�̤�<X�[=�'�=�O�=� �=�Ŷ=�E�=q]�=��l=,=�i�<�/�����֝M��J��+����   �   �1 ��� �ڪ���Ew𽈩½�W���?�\��� L׺���<PL	=\;=Z�Y=��b=�]R=��%=L��<@Fj�	�{g��?�����-��^��������̱��§��|��6���:xr�K�E���S�ҽ"�{�l
ʼ@I�; >=�GZ=�=��=�'�=��=���=�aO=l�<�ݳ;����vV�����g$߽����M��   �   iq���o���b�:M�N0��!�OJؽ�����#��7�\c<(�=�fO=��{=��=\�=(�p=�8=$�< ź����捽��۽d��v7�c0T�vh�hcq�f�o�o�b�{M�J0�H��Dؽ�
��b�#��7��bc<b�=�eO=��{=���=� �=��p=n�8=��<@!ƺT��d퍽b�۽�h��{7��5T�h��   �   @ŧ����9�������|r�8�E�=���ҽ��{�dʼ�4�;�<=�GZ=���=�=i)�=��=��=*hO=��<)�;����~iV�럧��߽g���H�!- �(� �s�� ��tp��½1S��l?����� ׺,��<�K	=� ;=��Y=X�b=�YR=��%=�|�<��j���Rm��V����-��^�������������   �   &�۾d�׾��˾�����7��L���ۢG����T���*�@�8����< �[=N(�=xP�=��=Ƕ=�G�=!`�=:�l=*4=�|�<0׼����֏M�^C��V���3X���~��(�����������}s��4��D㼈�=���~;D4�<̕�<�>=:51=�.=Π=��<����zr
���
��<&7�0s��;�����ũǾ��վ�   �   ����?������X供ž�졾�o{�$�5���� x�p\o�D�<��U=�ʗ=���=�U�=aW�=��=nk�=<�=r'�= M="B=�j< B:�<����/���@ ��=5�.a;�|4�7!��j���ż�6p�@.���?�;��< ]�<�R�<|�=���<@��<��:8ؼC���f'�wP/�*�r��K������ �ྮN������   �   G�"����w����Y�^����S���]�`�����L�޼�C�<��J=SR�=��=R�=���=���=��=�T�=��=3��=6�~=:(D=��
=@h�<��< ��9p�ֻ��8�X:c��Sm�ДZ� �-��XԻ�А� `�;�[?<���<���<��<���< �y;�폼8 K�9@���<)^�8���¿�ƽ�,��Х�OD��   �   ��9�.\6�<�+��b�]���n޾�v��i���.-��Dɽ�* � 5<�g==˘=@��=2j�=�'�=���=ʐ�=l~�=���=Zz�=�*�=oH�=�z=.K= =��<,r�<��[<0q�;�":; ⵹�� � ���`w=;��;�-<��O<�t9<��;�"��s��)�����{$:��Ճ�Mů�ef޾�-�|���h+��6��   �   �%L��:H�ݺ<���*�.��:������XŎ���B��x�hH��5;`1=�V�=��=6�=\-�=.��="4 >��=��=J4�=���=���=�#�=|w�=�:p=��F=d�=��<|�<Pf< Z�;`I; �,9 �A� �V9@�; �;P��;@/T;����$����-@��ů��^�^1T�c4����þ%����=� �*��<�hH��   �   ��W�ˬS��G�\�4�ܾ�����̾.���hP�V6����b� }��(U(=���=;�=LT�=hM�=Œ>*�>��>���=���=Tm�=|�=�N�=���=m��=��t=�[J=�� =8��<���<p�G<pP�;@�:@6��� �@F��D=:@ڀ:����'.������a�E�ĽI���d�a���>�о&�0C���4�ƐG�t�S��   �   A��J:���������#e��"@�s����A3��
E[�K���n�D�H@<�Q=D/�=@'�=�,�=nX�=+R�=�h�=��=B��=7m�=y��=a�= ��=�M�=f}=F
c=&�L=�,:=��+=d*!=:�=�F=��=�=�a=T:=8��<h��<@���*��q]��ӻ��p�ՠ��j1�]��97A��e��%������:���   �   M`��!����o��a���	a�Z�<����
}徝���w2V�r���0;���$<��S=�w�=�i�=kr�=F��=���=���=e��=���=pt�=��=���=Yj�=I��=��g=z�N=��9=$_)=�I=��=~�=�&=�7=��=�=�=LW�<@,�<�:7�����ǥ�bX�KHj��ͪ��L�!���=���a��ˀ��q�������   �   .���^㍿�"����s��)U��s2�ۛ�4ؾI���6�G�Ehݽ�H ���e<8�[=��=���="�=�l�=h�=�O�=�4�=���=x;�=Gn�=��=b�g=f�D=8W'=�=	 =�q�<�3�<+�<��<���<"�	=*=�w=t�=.j=q�<�*;X��������YY�����aܾ����3�iXU���s����э��   �   �<��&Ձ�
eu��_�+�B�*�"������þL�����0�w⽽���t�<Gg=�@�=�N�=0��=N\�=�V�=���=�5�=&9�=ˉ=Zs]=ċ)=� �<��< ]<�P<@��;�#�;(�<�H<*�<T�<���<0�	=>~=|{ =��=���<h>3<0���[i�]罛�>��k��� ƾ��%�"��BB���^�U�t���   �   �"i�n�d�;X��GD���*��i�-
�J�����l��Y�k����χ��(�<N�s=6#�=©�=<��=��=���=�ج=&�=�a=�G=�k�<P �;�b�����>ݼ�T��X����ּ�����4��P���p<0q�<���<J�=jv(=��(=�n=��<`!��������d�qq���zR�:���*�K\C�zW��}d��   �   �E�'B��57��&��F�ӊ�0�������@����N�V��J��=@�}=α�=RI�=���=�T�=�A�=ƌ|=�/=p�< ʺ �ż��7��o�V���7������Δ�������\q�Ȯ2� Tܼh�!��O�;�a�<�	=H�+=f;=��0=��=8bZ<�̌�ev���A�?�{���+���G쾸���$�C6�J}A��   �   ?� �����������p龯���%��,�]���g橽t���p8%<ʰ)=ځ=��=⌧=���=�^�=�3^=�=�X�;Ь���eU����z�߽����!��F�u��
^�b��7c㽘7��\�{��Z� �C���<<W�<��'=�H=��N=J6=Լ�<0�;(H��柽tK�ԏS�c����v���}�!���j����   �   |f��|@���F���о�T�����Z�e�RA%���Խ��[� �?���<?=�X�=|k�=s�=;Ƀ=��I=8%�<�������B��Ԇ���h@B��`�kVt�`q}�J�z�s�l�c�T�s�5���O�ؽ�1��~b���޻�<�<>B=j�N=��g=@�a=�9=h�<���tn$��*������eT����]^��Y˾ce㾟A��   �   ������������ԙ�,��N=W�j8$��9�2ɉ��S�0��;��<r�K=�y=詃=�t=~�>=<��<�V���-�������@SA�C�u�o���X����o������~��������י��.���AW�<$�1?�X͉�$_����;���<�K=�y=��=t=��>=��<p��V�-�Q�����MA��u� ��������k���   �   �j}��z�|�l��T�Ў5�8��,�ؽ-���[���޻DB�<NC=&�N=v�g=��a=ث9=�<���nx$�B1������jT�����a���\˾�i��E��j���D���J�\�о�W��>����e��D%���ԽL \�`�?���<?=Y�=\l�=��=t˃=��I=�4�<���b��;���}�ˡ��:B���_��Ot��   �   ]A�U��BY����[�y1����{��S�X�C��<�Z�<^�'=B�H=��N=H6=0��<p�;4X��W럽�N�#�S�����y��s��0��m�D��� �@��������t�~���i����]����ꩽ ����,%<|�)=ځ=5�=��=���=}a�=Z:^=R= ��;�����VU������߽������   �   a/�����u�������Qq���2�tEܼЀ!�0m�;Pf�<�	=&�+=J;=��0=��=�PZ<�،�mv�Oｫ�?�8}���.��K쾒��)�$�{!6��A�g�E�kB�87��&��H����v��������@�T��D�V��HJ�=��}=<��=@J�=j��=�V�=�D�=��|=X%/=x"�<��ȺDyż��7��_�%���   �   �%ݼl=������H�ռ<���8�4� ����<v�<���<��=�u(=>�(=�l=��<�P!�N�����gg��q����TᾹ��?*�7^C� |W��d��$i���d�=X��ID�P�*��j�F�鋩� �l�V[�����DՇ��%�<Ԓs=|#�=l��=R��=���=���=f۬=Y�=P"a=vP= ��< Y�;�3�$����   �   �,]< q<���;�X�;��< �H<�0�<�#�<���<��	=0~=�z =\=���<43<��j`i�=`罻�>��l��Aƾ��m�"�)DB�D�^��t�Բ���=��ց��fu�j_�r�B�<�"�{���þH����0�`佽�����<�Fg=�@�=O�=���=i]�=X�=���=*8�=�;�=4Ή=�z]=��)=D�<Ĩ<�   �   Z\'=
�=� =hy�<P:�<<0�<���<���<Ԡ	=X=�w=ֆ=4i=@n�<��);t��٥�� ��N[Y������ܾ���	3�YU��s�����ҍ�ԇ���㍿e#����s��*U�lt2�s���4ؾ����(�G��iݽrJ �p�e<��[=��=I��=�"�=�m�=i�=3Q�=t6�=`��=�=�=�p�=6�=��g=��D=�   �   ��g=��N=~�9=�`)=�J=��=&�="'=�7=��=j=��=DV�<�*�<�K7�����ȥ�Y�<Ij�<Ϊ��M꾘����=�'�a�̀�r������`��r����o������sa���<�, �l}�䷣��2V����`1;���$<��S=�w�=�i�=�r�=���=j��=.��=��=x��=bu�=$��=¤�=�k�=z��=�   �   �}=�	c=��L=�+:=��+=�)!=��=hF=J�=�=�a=H:=,��<���<Х��T���]������p������1�t��N7A�#�e��%��!����:��@��F:���������#e�g"@�X����3���D[�������D�XB<8Q=f/�=V'�=�,�=uX�=&R�=�h�=ܧ�=4��=m�=d��=a�=ٹ�=zM�=�   �   :�g=�N=$�9=�a)=�K=��=V�=f(=L9=<�=�=@�=�Y�<�.�<�&7�4��@ǥ��W��Gj�Cͪ�zL�Տ���=��a�wˀ�cq��d����_��Ɣ��*o�����ja�̠<�l��:|�����n1V����z.;�P�$<J�S=Mx�=[j�=�r�=У�=���=F��=0��=���=tu�=0��=ۤ�=�k�=���=�   �   ]'=��=� =@|�<�=�<$4�<p��<t��<p�	=$=|z=�=�l=�u�<�)*;��ἅ������xXY�����Vܾ���3�yWU���s����Hэ������⍿."��{�s��(U��r2����2ؾ6�����G��eݽ�D �H�e<��[=��=���=�"�=�m�=<i�=dQ�=�6�=���=�=�=�p�=e�=��g=H�D=�   �   �0]< v<���;�h�; �< I<7�<�*�<��<��	=F�=& =��=h��<pL3<d��Wi�9Z���>�oj����ž�
��"�\AB�!�^���t�����;��>ԁ�Icu�O _���B�ݍ"�����þ����Y�0��޽������<�Jg=B�=�O�=���=�]�=XX�=��=^8�=<�=dΉ=�z]=
�)=|�<�Ũ<�   �   �#ݼ`:��������ռ�~��0�4�@6����<�~�<���<��={(=��(=s=�(�<�� ��������b��q�/���1P�٭��*�xZC�xW��{d�l i�E�d�
9X��ED��*�h���)���0�l��V�O�����P3�<��s= %�=���=��=$��= ��=�۬=��=�"a=�P=��<`]�;�0�D����   �   �.��F���j���َ���Nq��2�\=ܼ(o!� ��;�p�<	=�,=x;=��0=��=�wZ<4���F]v����?�y��l)���D�����$�6��zA���E��B��37��&��D����f
��u���r�@�ԧ�6�V�@�I�|=0�}=��=�K�=D��="W�=�D�=4�|=�%/=l#�<��ȺLxż0�7�@_�����   �   A�����X�w��RZ㽶/����{�O� �C���<�e�<4�'=��H=�N=�6=\��<�K�;�7������5H���S�ݖ��ys��6z����h��	�ڟ ����S������l�[���V����]�X��k੽t����V%<�)=�܁=�=d��=g��=b�=6;^=�= ��;����PVU�I�����߽e��w��   �   �j}���z��l�s�T��5�`��E�ؽ�*��$W�Џ޻�L�<�H=T�N=v�g=��a=Ƶ9=�#�< ��zd$��$������`T����Z��5U˾7a�2=��a���;���B羻�о+Q��t����e��<%���Խ��[� �?�� �<|?=�[�=6n�=4�=Ĩ=��I=�6�<�������:���}꽰��x:B�p�_��Ot��   �   ��������Ƥ��jԙ��+���<W��7$��7�ǉ��J��ڢ;t��<.�K=��y=���=�t=�>=P��<�Ù���-�$������HA��u�����ࢥ��g�����������љ��(���7W�z3$�@1�`�p=�`��;8�<��K=ޑy=���=bt="�>=4��<���Ɯ-�������MA��u�󋒾�����k���   �   jf��`@���F羍�о�T��P����e�}@%�,�Խ��[��?���<?=�[�=�n�=� �=e΃=��I=�E�<@a�´�|3���t꽐���4B�)�_�It��c}���z�Ȋl�¶T� �5�.��t�ؽ�%��bO�0e޻HS�<�J=p�N=6�g=2�a=�9=�< ����m$��*������eT����T^���X˾We㾏A��   �   8� ����������}p�q�������]�Z���䩽L���H%<$�)=�܁=��=}��=(��=�d�=�A^=(=��;�y���GU���O�߽E����;�����S�޷�HR��(��Ė{��F��nC���<<j�<��'=$�H=`�N=�6=,��<��;�F���埽\K���S�Y���}v���}����j����   �   �E�"B��57��&��F�������������@�T��l�V���I�:=h�}=J��=JL�=���=Y�=�G�=ޚ|=&./=T7�<@Ǻl]żB�7�O�<���5&��遬���������0Bq�~�2��,ܼ�U!�`��;,v�<z	=,=�
;=��0=��=pgZ<4ˌ��dv����.�?�{���+���G쾷���$�B6�H}A��   �   �"i�n�d�;X��GD���*��i�
����#�l� Y�Q����ʇ��.�<��s=(%�=��= ��=���=%��=Pެ=��=h*a=�Y=���<`��;����l���	ݼ@!��0���$�ռ�k�� �4�@n����<0��<���<:�=�z(=��(=q=�"�<�� ���ҩ���d�fq�� ��vR�8���*�K\C�zW��}d��   �   �<��'Ձ�	eu��_�%�B� �"������þ%���A�0��ώ<��|�<lIg=B�=OP�=R��=�^�=�Y�=���=�:�=�>�=�щ=T�]=>�)=$�<�ר<�U]<��<@"�;���;��< I<�?�<L1�<\��<��	=��=�~ =܂=���<�B3<�	��8[i��\罏�>��k��} ƾ��$�"��BB���^�T�t�𱁿�   �   /���_㍿�"����s��)U��s2�ӛ��3ؾ2�����G��gݽ�G ��e<��[=w�=��=f#�=�n�=7j�=�R�=&8�=^��=�?�=s�=�=��g=4�D=(c'=،=P =d��<�F�<�;�<,��<���<Ԥ	=�=~z=p�=�k=s�<�*;l��򣒽���YY�����`ܾ����3�iXU���s����э��   �   O`��"����o��a���	a�X�<����}徔���Z2V�7��^0;�`�$<��S=#x�=\j�=s�=#��=��=��=���=y��=�v�=s��=:��= m�=+��=b�g=8�N=�9=4d)="N=ʋ=��=�)=:=��= = �=�X�<@-�<�57�N���ǥ�ZX�GHj��ͪ��L�!���=���a��ˀ��q�������   �   �nп��̿�¿"G��w���;탿7�U�p&%�ۏ�g
����L�^ӽ���\��<�'�=>ٶ=>�=	��=�]�=��=l+�=�+�=)��=a�=0ŕ=��=,Wn=�DY=,AK=(*D=p|C=NLH=fWQ=�]=��i=r�t=�y=�t=��\=��+=왭<�4;� �s��G�4�_�m����r��k'��~W�&����f���|���¿ÿ̿�   �   {�̿Sɿ�Ⱦ�M��~W��������Q�1"����ΐ��#�G�Z�̽,j���<��=�>�=xZ�=�i�=d��=L��=���=�}�=R��=t��={8�=>Po=�R=�H==��/=�r*=,=f�3=.�?=��N=��^=:�l=l�t=�q=��\=X.=P��<��4�h�-���kZ��ר��k�.2$���S�.������q���̾�?Mɿ�   �   $�¿�`���Y������(���/�u���F��*��$߾e{���h9�󴹽 |��x�<]�=8�=v��=*��=c�=89�=���=��=�Ӓ=8@t=��E=j8=̏�<���<<��<(�<X�<���<�
=n2#=��<=�QT=^�d=��i=\=|5=h��<@5����G�ۄ�nUJ��۝������V�G���v�7���P����:���H���   �   b岿ʯ�ʋ��[���x����`�6f5��:���ɾ�Ň�lJ#����0S���=KG�=`%�=|L�=�N�=�N�=�"�=�{�=T�{=�	<=|_�<�/�<�p;�/���j6�H~T��$7�0�ɻ@��:@2<���<��=TA)=��H=z�Z=@�Y=.>=h��<I�;�-��z���@1������;�?���5��a��M������@��򙯿�   �   a����ۛ�����f���,�k�":F��5������C�g� g���m����>�=_��=�&�=8�=�5�=V�=7��=jJ=L�<p5<��O��T��LC�<�q�����븆�2	z��S�����PGӻ��%<���<��=� B=�R=�ZF=nE=Up<�l��Ɠ�*s�F)n�hX��^������E���j��
���"��Z����   �   �|��t%��L�{��^e���H�U�'�%��G˾^���u;�E�н���(<�6=E��=�H�=�{�=���=��n=�X=ld<�_���.�ؑ�I�ƽ�����,� ��d\꽸���(��&�6�$䡼 {T;�1�<z#=65B=��J=��/=Z�<`�\��@��,۽Jc=�>���1�ɾ&
�T�&�q�F�-�c�X�z��τ��   �   ]v^��Z��N�t�;�#��Q��Zؾ�6��*Tb����<�������pq�<��H=3I�=:��=�s�=�`T=���< i;8a �uX��j?޽���ޜ:��W�T=k�H�s�|p�kb���I��}*����[X½$fr�@o׼��;��<�A'=�IH=J�D=��=(m<x���L�����
�1�\�ͳ���OԾ�+�{u!��9��>M�z�Y��   �   ��.�1�+��I"���9��fӾ.���\u��j&���Ľ��(��C�:�=fU=��y=H�s=�D=g�<@�L��H*�4�����dC��.x����W���,���Z��xp��̫�7����S�� ^V��4"�?P߽7���x�ɼ@T�;\P�<xj<=�S=z1@=�� =�;���wԲ����ȣi�:���w;j������
� ��+��   �   ���%� ����ve۾Y_��h����
q�Β-�#@ཾ�k�0>t��*�<��%=f�X=Z]a=0?=�n�<@���.�LE�������`��ϓ�b�����վE�ƙ��I���� �j���i۾,c�������q���-�BFཆ�k��Ut��#�<�%=ĶX=|_a=#?=�z�<�o���.��=�����`�4̓�I����վKﾔ����   �   6V��l���ǫ������P���XV�0"�bI߽�����ɼ�z�;�U�<Lk<=�S=�.@=,� =p��;>���ڲ�+��%�i��"���{;���}��Ҧ �h+�|�.��+��L"����=���iӾ1��;au��m&���Ľ�)����:�}=.U=�y=��s=D�D=�u�<�L��;*��+�����dC��'x�+
��tS��p(���   �   �s�up���a��I�Rx*�H��FQ½[r��^׼ [;�<�C'=�IH=�D=�~=� m<𯫼S���"�
���\�����}SԾ�-��w!���9��AM���Y�ry^��Z��N�
�;�	�#��S��]ؾF9���Wb�������а��hl�<�H=�I�=���=v�=�fT=$��<�;�S �?P���5޽ ����:��W�46k��   �   J'�����7S꽯���!��6�6�ӡ���T;�:�<&=F6B=��J=��/=�S�< ]�J�@��1۽�f=�}����ɾ��t�&���F���c�B�z�oф�~���&���{�jae��H�<�'��&��I˾�_��cx;��н��0�(<�6=���=�I�=�}�=!��=��n=\a=�d<(�_���.�Hϑ�|�ƽA�H���   �   À��鰆�8�y�bsS���<���ӻ��%<��<��=z"B=hR=�YF=�C=HHp<$v��yɓ��u�,n��Z����X����E���j����T$������ƚ�� ݛ�ߙ������6�k��;F�7���������g��h�
�m� �.�=x��=O'�=~�=�7�=��=���=NrJ=�_�<�c<��O��E�,=C���q��   �   H=6��QT�8�6��yɻ ��:�52< �<��=vD)=~�H=~�Z=^�Y=b
>=��<�2�;2��}���B1�����;A�.�5�4a��N������.A������沿-˯�ٌ��P��ey��3�`�`g5��;��ɾ�Ƈ��K#����h#S���=QG�=�%�=`M�=7P�=�P�=<%�=�~�=d�{=�<=8r�<hD�<@�p;PԴ��   �   
�<Ÿ<!�<'�<Г�<
=�5#=V ==�ST=��d=�i=��\=�5=���<pF����G����VJ��ܝ�������h�G�ܔv�������;��kI����¿�a���Z��@�������+�u���F�y+��%߾|���i9�����~��`�<b�=U8�=��=��=Cd�=�:�=f��=��=i֒=(Ft=��E=R?=,��<�   �   L==� 0=�u*=�
,=��3= �?=h�N=��^=��l=Եt=�q=��\=�W.=���<��"�h�����plZ��ب�wl�2$�N�S�v.�����wq��;��Mɿ��̿�Sɿ!ɾ�rM���W��������Q�t"�P�����v�G���̽�j���<��=,?�=�Z�=�i�=���=��=���=�=���=���=�9�=zSo=V�R=�   �   NDY=�@K=�)D= |C=�KH=�VQ=�]=z�i=�t=��y=�t=X�\=d�+=���<�5;���s�-H�x�_�����*s���k'��~W�6����f���|���¿ƿ̿�nп��̿w¿G��g���)탿�U�N&%����8
��D�L��]ӽT��h��<(�=aٶ=*>�=��=�]�=��=i+�=�+�=��=�`�=ŕ=��=�Vn=�   �   ZL==� 0=>v*=(,=2�3=��?=:�N=��^=�l=�t=0�q=��\=&Y.=\��<P���h�t���kZ��ר�0k��1$�L�S��-��S����p��G̾��Lɿ	�̿�RɿPȾ��L��W��d�����Q��"���$���"�G���̽�e�h �<i�=�?�=[�=$j�=��=��=���="�=���=���=:�=�So=z�R=�   �   �<4Ƹ<�"�<�(�<(��<f 
=J7#=
==hUT=�e=F�i=�\=�5=���< "����G���FTJ�۝�z��l��|�G���v���������.:���G��N�¿!`��Y��Π��s�����u���F��)�6#߾Nz��g9�z����t��\�<��=*9�=���=l��=�d�=�:�=���=��=�֒=bFt=��E=�?=؞�<�   �   �:6��NT�(�6�poɻ�ȿ:@=2<0�<P�=�F)=D�H=��Z=��Y=v>=��<@e�;�)�#x���>1�����O;�>���5�	a��L�������>��Ϙ��7䲿�ȯ�����N���w���`��d5��9���ɾ-ć�BH#���� S���=I�=�&�=(N�=�P�=�P�=}%�=�~�=��{=<=�r�<E�<`�p;Pд��   �   k���v����y��qS�>�����P�һx�%< ��<@�=&B=�"R=�^F=�I=�fp<<b����
q�z&n��V�����/��1�E���j�X	���!����������`ڛ�@���$�����k�'8F��3���沮���g��d��m����.�=���=�(�=l�=b8�=N�=̲�=�rJ=|`�<�d<x�O��E��<C�V�q��   �   '�{���fR꽲��� ����6�(͡��U;�A�<*=�:B=��J=��/=Pd�<�h\���@��'۽/`=�4�����ɾ��]~&�%�F���c���z�m΄�{���#��^�{�#\e�7~H�/�'�K#��D˾�[��"r;���н���)<X6=˷�=^K�=�~�=к�=��n= b=�d<h�_�@�.�ϑ�L�ƽ
�%���   �   �s��tp���a���I��w*�����O½Xr�X׼ �;0 �<\H'=lOH=��D=��=X-m<<���g�����
�
�\�(����LԾ�)�%s!�d�9�<M�o�Y�?s^���Z��N���;�I�#��O�/Wؾ�3��sOb�.����������<��H=L�=��=w�=
hT=��< ;LS �P��y5޽��~�:���W�6k��   �   $V��l���ǫ�V���UP��XV�|/"��G߽|�����ɼ ��;�^�<�p<=R	S=H7@=� =���;.��Mβ� ����i����s;����i��M� ���*���.�=�+�!G"���4���aӾ�*���Vu�f&��Ľ��(� ^�:�=�U=��y=��s=D�D=hx�<�
L�;*��+��{��RC��'x�#
��jS��e(���   �   ���� �{��Qe۾(_��,���
q�)�-��>བ�k��/t�3�<��%=��X=:ea=Z)?=h��<���:�.��6��W��z`��ȓ�K�����վ[�Z������}� �~��`۾[���}��Tq���-��7བ�k�8t��;�<��%=ʼX=�ca=�%?=l~�<@\���.��=��֧��`�.̓�B����վDﾊ����   �   ��.�*�+��I"��j9���eӾ�-��\u��i&���Ľ��(����:�=�U=��y=\�s=��D=��< vK��.*��#������C�!x�Q��=O���#���Q���g���ë�v����L��3RV��*"�`@߽����8�ɼ ��;he�<r<=�S=$5@=,� =0Ŏ;��� Բ�����i�3���w;e������	� �}+��   �   [v^�
�Z��N�j�;���#��Q��Zؾ�6���Sb�G������d����x�<|�H=7L�=$��=y�=�mT=���<��;XF �H���+޽���D�:�1�W��.k���s��mp���a�a�I�Pr*����2H½�Kr��E׼� ;)�<�J'="PH=ĳD=
�=8m<����ࡐ���
��\�ǳ���OԾ�+�yu!��9��>M�z�Y��   �   �|��t%��J�{��^e���H�H�'�	%�dG˾�]��Lu;�8�н��	)<�6=÷�=L�=��=��=̫n=@j=P�d<�P_�6�.�jƑ���ƽl����h!���X��H�	��N��|�6�$�����U;L�<Z-=z<B=�J=^�/=�^�< �\��@�b,۽0c=�6���,�ɾ%
�T�&�p�F�-�c�Z�z��τ��   �   b����ۛ�����e���&�k�:F��5�o�ﴮ���g��f�ʆm��s�L�=P��=#)�=��=%:�=��=���=�zJ=�s�<�<��O��6��,C���q��w�����$�y�NcS�j���𼼠�һ&<̠�<��=j(B=�#R=�^F=FH=�\p<<j���œ�s�3)n�cX��[������E���j��
���"��[����   �   c岿ʯ�ˋ��\���x����`�/f5��:���ɾ}Ň�"J#�M��HS���=�H�=4'�=�N�=�Q�=�R�=�'�=߁�=��{=X<=���<�Y�<`xq;�q���
6�HT�X�6� ɻ ��:�\2< �<Z�=�J)=غH=�Z=X�Y=>=t��<T�;-�vz��l@1������;�?���5��a��M������@��󙯿�   �   '�¿�`���Y������(���-�u���F��*��$߾R{���h9�~����y��X�<M�=69�=��=0��=�e�=o<�=n��=)"�=4ْ=vLt=��E=�F=��<��<tո<1�<D6�<��<�%
=|;#=N==�WT=0e=0�i=^�\=V5=���<0.����G����^UJ��۝������U�G���v�8���R����:���H���   �   |�̿Sɿ�Ⱦ� M��~W��������Q�."����Đ���G�$�̽i�H�<!�=�?�=@[�=|j�=���=���=���=D��=���=l��=�;�=HWo=N�R=BP==�0=�y*=�,=H�3=`�?=z�N=��^=<�l=Ʒt=��q=�\=Y.=���<���h����vkZ��ר��k�/2$���S�.������q���̾�@Mɿ�   �   ��-M�����h�忮�ʿ̬��H����\�8>$��� 9��y�+�b���Rϻ"�*=�`�=L�=~��=t��=�.�=4��=��=
��=n�=�}k=@1I=FM/=�<=*z=��=��*=�?=��W=�r=`�=CЏ=\�=n�=�{=|5=0Hx<�������<�`����w�D'��o_�6Z��[�����˿��~��uN��   �   vm�8������⿾�ǿ�쩿Cފ��Y�51!���K���FY'��˒��Y���--=Tݖ=I�=J�=,m�=�%�=�¾=9�=o#�=H}w=fL=�q'=�=�T�<\6�<�'�<FT=��#=�y@=�+_=�s|=��=�=}�=$z=f6=ԇ�<@�߼&3���8�
������#��S[�#Ջ�0����%ȿx:��������   �   c���|�����@"׿����ŋ��,ԃ�ʜM�R�ZԾT���;������ A�� �3=��=�b�=� �=�9�=Y¸=:�=}��=tZ=Ɯ =0��<��<8y <��f;��7;P[�;ض:<d�<�F�<�u#=��L=j�o=g4�=�9�= t=��9=��<�������)�o玾7�پ"���dO���������+��F׿��꿪x���   �   @����'Pؿƿ�Ʈ�[����q�a�;��n
�ľ��zt����4DS� .�;J|<=�G�=�ϫ=D��=�|�=�(�=�k= �#=��<�{#;H�l��Y� (��E0���/�������k���e���do<� �<H�0=��Y=��n=�h=(==DN�< �H��"��b���)~�մþ�����<��r�Kb��썮���ſ�׿[���   �   Oο_�ʿ܈��V+��/9���j��R%U�`�$�_������7O�_�۽T��8�j<ҫD=�b�=�F�=J
�=1�=
>=pa�< P�8t�ռ��S�����$��,�ڽ���s��ҽ�����O���P=�\��� p]��I�<�Y=�ED=X�S=�_==��<����.�G��U��%V�M�����/%���T��������v���俿��ʿ�   �   ZN���a���c��� ���ք��`�h�4�m�
�K�ɾ3��@y%�Q8���?��8��<�6I=�e~==��^==�=<����>]�rI���6��2"���<���N�[;V��R��E��H.����]"޽����d�'���0�(�l<��=�73=:y7=�[==2<�L�m����4)������pɾ�Y
���3�Ş^���1������5�   �   EŒ�V������+gy�H�Z��u7�9���Fe����S�:x����V�@�I�P)�<�G=(@]=��B=4a�<`h8;v��!ӛ�����2���d��;������z���{��󙩾@[��Ɏ��r�=�B���X=��L4S�(�x��X<�f=�>(=X�=���<`�� <`������Q��v��b:ݾ�P�[5��<X��?w��凿�ۏ��   �   �/i��Ee��X�\CE��,�?��Om侷ǫ��
q�/�j��0ּ�+F<ԥ=��;=��/=�2�< �8���}������X����"9����ϾЈ�!����������1쾏վ⍷��7���g��M%��dҽ|W�FJ�d7�<�V=x�#=v=�<<�~Ǽut��Y���i��f����߾X��)�d�B��'W�`Qd��   �   Z�0���-��I$�����5���վ<#���x�)L(� �ǽC2� h2��A�<H� =f�%=`��< �];>H�i���3��'l��𡾆�Ͼ����`u��"�I-���0���-��L$����'8� ־�&��Q x�JP(� �ǽbK2� �2��<�<"� =��%=x��<�^;�=�4��5/��!l��졾��ϾN���kr���"��-��   �   ����h����+쾱վ����4��5�g��H%��]ҽTW�X*J��?�<RX=��#=Xs=��;<�ǼSz��]��i�dj��ه߾�	�܃)���B�A+W�Ud�L3i�HIe���X��FE�~,����/q��ʫ�.q�z2��n���ּ�F<
�=n�;=R�/=�>�< ��80���t��j��#~X�����4����Ͼ[��i����   �   kv��^����V��#Ŏ�,�r�f�B�J���5���(S�8�x��2X<�i=�?(=@�=�<p���D`�8����Q��y��>ݾ�R��]5��?X�Cw��燿�ݏ�9ǒ�X����wjy�3�Z�Rx7�C��ྐྵg���S�*}��D�V� �I��&�<�G=�B]=��B=p�<@9;���ʛ���у2�P�d��7����ؠ���   �   4V���R��	E��B.����N޽`헽��'�~0���l<��=":3=�y7=:Z=�.2<|X�箰��7)�����sɾl[
�)�3�z�^�`���{3��n����DP���c���e��""���ׄ�\ `�k�4��
���ɾ�4���{%��;��LG�� ��<"7I=h~=⽁=��^=6=x>=<����p.]��?��J1�p,"���<���N��   �   Q����=�ѽ�쳽H��XC=�,ຼ �:��V�<n^=xHD=��S=�_==���<�p���G�-Z��(V�]��v���%��T�J	������Qx���濿z�ʿ�Pο�ʿw����,��z:���k��''U���$���񾑜��wO�P�۽�����j<ҫD=Bc�=MH�=��=64�=6>=�u�< (�80|ռ
�S����������ڽ�   �   �60��|/�.������U�� :��p�o< -�<��0=��Y=��n=�h=�==�J�<��H�N%��?���,~���þ����<�cr�\c��!�����ſq�׿ө㿹��r��{Qؿ�ƿ�Ǯ��[��8�q���;��o
����Jt�,��GS��"�;.|<=6H�=�Ы=���=:�=�+�=T�k=��#=l/�<�9$;��l�`=�F��   �   @g; 38;p��;��:<$�<|R�<�z#=��L=:�o=\5�=a:�=ft=�9=���<�������]�)�s莾��پ���eO���������n,��B׿��꿻y��t����������#׿� ��b����ԃ���M��R��ZԾ������� ����3=+�=4c�=��=I;�=Aĸ=��=N��=
Z=@� =���<P�<P� <�   �   l]�<�>�<�/�<�W=�#=J|@=�-_=�u|=S�=|�=��=$z=�e6=؅�<��߼\4���8����Π羙�#��T[��Ջ�����N&ȿ;�j���@��m�|����M��ǿ�쩿}ފ�Y�s1!�g�ᾂ����Y'��˒��[���--=�ݖ=��=�J�=�m�=�&�=�þ=d:�=%�=ހw=bL=,v'=8#=�   �   H<=�y=<�=��*=.?=d�W=ƨr=7�=Џ=:�=�m�=��{=05=�Fx<�������<�����.x�e'��o_�LZ��p����˿�濊��xN���)M�����U�忛�ʿ̬�jH����\�>$�|��8��/�+��a��Mϻ��*=(a�=^�=���=~��=�.�=8��=��= ��=j�=�}k=1I="M/=�   �   �]�<4?�<40�<.X=r�#=�|@=�._=*v|=��=��=$��=Dz=g6=���<@�߼�2���8���������#��S[��ԋ�㨪�p%ȿ:�]�����.m�������Z�?�ǿ쩿�݊�Y��0!�9�ᾨ���UX'�$ʒ��H��r/-=ޖ=��=�J�=n�=�&�=ľ=j:�=%�=�w=nL=Jv'=V#=�   �   �g; 98;P��;H�:<��<8T�<�{#=��L=��o= 6�=K;�=�t=ص9=L�<����{���)��掾?�پz�dO�t���x����*��j׿��꿡w��R���j�����G!׿�������Ӄ���M�7Q��XԾM������n��� ����3=)�=�c�=g�=�;�=lĸ=��=g��=*Z=^� =��<��<� <�   �   ~60��{/����T���S�� ��@�o<P0�<��0=�Y=4�n=�h=�==$U�<�H�s ��ڠ��'~�f�þ���[�<�r�\a��Ռ��q�ſ��׿����翐�㿽Nؿ.ƿ�Ů��Y����q��;�vm
�󼿾�t����&>S� T�;N�<=�I�=�ѫ=���=��=5,�=��k=�#=�/�<`<$; �l��<����   �   �潼���ѽ`쳽oG���A=��ܺ� �2�[�<�`=|KD=\�S=|d==��<@c��P�G�R�/#V��	��_��%���T����<���Bu��Y㿿�ʿWMο��ʿ.����)���7��_i��4#U���$����ۘ���N���۽*��(�j<̰D=�d�=nI�=G�=�4�=�>=�v�< ��8�{ռ��S��������p�ڽ�   �   4V���R��	E��B.�N���޽y엽��'��t0���l<�=.>3=�~7=a=�S2<,?�����1)�����nɾ�W
���3�E�^�b탿$0��ԙ��V쭿nL�� `��$b�����Մ�5`��4���
�X�ɾ�0���u%�93���/�� �<�<I=�k~=��=8�^=:=�@=<����$.]��?��=1�d,"���<���N��   �   av��K����V��Ŏ���r��B�����4���&S�(�x��?X<n=E(=>�=� �<����2`��|��ĦQ�Yt��7ݾkN��X5��9X�C<w�䇿�ُ�PÒ�-T������cy�#}Z�s7�����߾Tb���S�Zq��^�V��I�P7�<RG=�F]=��B=Ls�< 9;`��gʛ����2�D�d��7����Р���   �   ����[����+쾔վx����3��ɏg�gH%��\ҽ�W��J��G�<l]=��#=�|=#<<�lǼ�n��6U���i��c���߾��~)�2�B�8$W��Md��+i��Ae�z�X�@E��,�����h�)ī��q��*�uc����ռMF<
�=��;=��/=�C�<  �8>���t��R��~X�����4����ϾX��e����   �   Z�0���-��I$�����5���վ#��mx��K(���ǽP@2��.2��J�<�� =��%=���< �^;�2�5���*��l�b顾��Ͼ5����o��}"���,���0�8�-�jF$�����2��վL��ux�G(�3�ǽ�62���1��Q�<�� =��%= ��<�2^;X<����/�}!l��졾��ϾL���jr���"��-��   �   �/i��Ee��X�RCE��,�.��'m來ǫ�#
q��.��h���ּX<F<d�=��;=��/=xN�< d�8֡�m��g���wX�&��G0�� �Ͼ�}辱��� �������#&쾆վ����0��r�g�]C%��TҽHW���I��Q�<�_=��#=�z=�<<{Ǽ�s���X�n�i��f����߾X��)�b�B��'W�_Qd��   �   EŒ�V������&gy�>�Z��u7�*�c�e��$�S�3w��:�V��cI��2�<^G=�H]=X�B=���<��9;�w�H������}2�1�d��3���z��.����q������bR��������r�;B�����,���S�(�x�XYX<�q=�F(=�=��<����:`�z�����Q��v��]:ݾ�P�[5��<X��?w��凿�ۏ��   �   ZN���a���c��� ���ք��`�]�4�`�
�)�ɾ�2���x%�C7��:�����< <I=0m~=���=��^=�!=xi=<$坼B]�6���+�(&"���<�S�N��,V���R��E�Q<.�����޽u䗽ʘ'�8M0���l<�=A3=�7=B`=�H2<�H�ݩ��`4)������pɾ�Y
���3�Ğ^���1������6�   �   Oοa�ʿވ��U+��.9���j��M%U�V�$�F��՚���O���۽$��`�j<��D=^e�=�J�=P�=�7�=�>=X��< ��8_ռ6�S�Cx��l���vڽ:�� u㽠�ѽ�⳽?��v3=��ĺ� 8� j�<jf=OD=^�S=�d== ��<����ƈG��Uｨ%V�D�����-%���T��������v���俿��ʿ�   �   B����(Pؿ�ƿ�Ʈ� [����q�X�;��n
�����@t�����BS��?�;\<=�I�=hҫ==���=�.�=��k=��#=<D�<��$;�vl�� �
�H'0��l/�6�����H<���˂�h�o<>�<
�0=��Y=��n=h=�==0S�<��H�J"��=���)~�ϴþ�����<��r�Jb��썮���ſ�׿\���   �   e��������?"׿����ċ��)ԃ�ƜM�R��YԾA���	��.��� ����3=)�=Pd�=H�=�<�=<Ƹ=��=0=�Z=� =���<��<�� < �g; �8;��;P�:<���<|a�<�#=&�L= �o=^7�=<�=pt=�9=��<��������)�h玾4�پ!���dO���������+��G׿��꿫x���   �   wm�:������⿿�ǿ�쩿Cފ��Y�11!���A���0Y'�I˒�`T���.-=ޖ=+�=<K�=�n�=�'�=+ž=�;�=�&�=��w=�L=�z'= (=Pg�<�H�<d9�<l\=D�#=�@=f1_=~x|=��=��=���=�z=8g6=T��<X�߼ 3���8�������#��S[�$Ջ�0����%ȿx:��������   �   �)�� &�3����|;�� .ٿv�����oT��_���ɾswu�����Xd$���< ?j=ť=���=R{�=Q��=��=N�=<̀=2@P=�#=L��<��<��<x̫<$h�<(��<h�=�A=�ji='�=���=/E�=��=$z=NZ=�Ƹ:��b�I�1R��)$о}�#�W�h���).��Raڿ���
��I�]&��   �   :+&��/#�i���n�'����տ�ϯ�������P�����žn�o�:���F&����<�Ti=�_�=JY�=:4�=��=���=�}�=:pc=��-=���<�.�<x�a<()<x�+<��f<�֩<m�<~c$=ĴP=��y=}ь=f��=�x�=j�v=�=�);�9Y��	�'�|�x�˾�y��S�2����I�ֿ���������\)#��   �   z������|���J�)|˿y;�������E�R<�:Ṿ��_���ὖ�����<�f=��=�-�=h�=P!�=�S�=(�J=d=!�<�k�:�)�����Ը�0#�����������;�)�<��= �<=J]j=䌃=�g�=$*l=��= �;*I=�b���%k��)�����m�G�DĄ�f��]̿��Q��S������   �   f�~���k��A���ۿ�m��C���]Pq�<Q4�o����Z��R�F�����D;¼��<��^=���=�g�=z1�=��b=^�=�ˆ<P�ǻ���>�E����'���YZ����xՐ��gk��\$���� ��9DZ�<t�=ҘK=j�c=��X=�I=��-<J��:�׽[P�o���H�O�5���r�����x��5bۿJ������u��   �   �2��7��2~�Sqݿ��ÿ~Ħ��N��^U��7�W�ݾgޏ�?�&�.�����X� b�<B\P=�Pu=�i=Z`6=��< �� ��^󂽡�½�+���4��$�V+���'��t��1���ٽ�V�� �@�\H��`��;�0�<v`)=r#9=��=���<�h���%��Z�-�m���V�߾q��}GU�'��E��	ÿ7sܿՒ𿦨���   �   ��޿�;ۿZGп�྿C���~��Q�h�8�4��(�PU��6�j�$R��#\�@���	�<�E8=�<=\=xR<,e����d���ɽH��t�?�czh�E����K��5���Z萾֩���~q��1K��������b������\��<N�
=��=���<�� �Bt�����m�������$4���g�� ���Y��{���g1Ͽ�ڿ�   �   J~��|����O��ȑ��C�����k���>���2+־�Ƒ��{4�������"<��<��=���<�I�;X��6B��S� �7�=���}��?���x���Ѿ��߾���8��`Ծ����ϣ�l���J����Qx��06"�p���Д�<��<$,�< DE;pC��X��F�4�-���Ծ���<���i�7��j2���/�� 굿�   �   m���25��������|��]��Z:�Ň�����X� ��Eq�@3J�p߃<H��<��<�H�;�J������Z�5�Y������¾��Js	����ʶ"��{&���#��}����eN��ȾT{��DCe�x�����nz��`3���<��<P�e<(�Q�j�l�H�����T�ŝ��%��/�l�7��Z��Az�劉�Q����   �   ��c��1`��%T���@��A(�5W��޾\��a_j�#��>����� �; ߰<l}�<�-�;@�ɼ䕽��22b������پ�z	��f%��Z>��3R��&_��c��5`��)T���@��D(��Y�|�޾�_���dj�����������0Й;�ݰ<��<�W�;��ɼ�ݕ�q�A,b�����]�پ�w	��c%��V>��/R��"_��   �   x&�k�#�9z�����H�\Ⱦ�w��Y=e�������hq��3���<l��<�e<��Q�N�l�}�����T� ���d)�q2���7���Z��Ez������������q7��۟����|���]��]:�9�����䋣�`Y� ��Mq�XDJ��܃<D��<�<`��;(5��﷠�
U���Y������¾d��%p	�O��7�"��   �   ��r�ᾎZԾ���Iˣ�����J�����p���+"�@h��\��<,��<,*�<�E;JJ��]��(�4������ԾN����<��i� 9���4��82��\쵿����Џ��,R��Γ������k�s�>�$��M.־:ɑ�
4�)������<|��<��=\��<0��;����9��� ���=���}�F;��us��0Ѿ��߾�   �   �����㐾����wq�&+K�L��f	潐����� ���|��<j�
=R�=h�<`� �$It������m�I	�����&4���g��"���[�������3Ͽh�ڿ�޿�=ۿ�Iп�⾿��������h�4�4�Q*��W��Z�j�4T��(\�@�
�<4H8=��<=c=��R<8K��^�d�f�ɽ4��f�?�zrh����]G���   �   ��*� �'��n�$,���ٽSN����@��1��0��;�<�<~d)=z%9=�=��<�p��)����-�N�����߾'���IU�X(���F���
ÿ%uܿ��Ϫ���3��9��)��sݿ��ÿ�Ŧ��O��*U�A9�_�ݾ�ߏ�!�&�u����X��a�<�]P=DTu=b�i=�g6=t�<�����Tꂽ/�½K ��5.�o�$��   �   Q���頽�̐��Wk��N$����� ��9j�<z�=0�K=�c=��X=|I=P�-<��D�׽�P����h���5�n�r�����y���cۿ������v�R�a���l�C��]�ۿ�n��+����Qq�[R4�����[��בF������>¼X�<��^=���=�i�=+4�=��b=H�=8�<�>ǻp�� �E�$���x���   �   �������@�`~��p(�;x8�<=�<=aj=4��=�h�=�*l=f�=0�;4L=�����'k�&+��c����G��Ą�< ��X̿����������+��|�S����K��|˿<��~�����E��<��Ṿ��_�"�ὸ�����<bf=��=/�=*�=�#�=�V�=�J=|"=x3�<���:��(�����   �    4)<��+<��f<�ߩ<$u�<�f$=��P=�y=OҌ=���=y�=��v=��=`);�;Y��	�D�|�A�˾Qz���S����~��ٸֿ����ؘ�O���)#��+&��/#�����n��'��ܮտ Я�ʳ���P����'�ž��o������&�8��<`Ui=``�=�Y�=5�=8��=(��=w�="tc=l�-=���<L9�<`�a<�   �   \�<̫<�g�<���<�=��A=�ji=�=|��=E�=e�=�z=�Y=���:� c���`R��f$о�}�N�W�����C.��laڿ�����I�`&��)�� &�3����c;���-ٿ]�������nT�j_���ɾwu�l����c$���<r?j="ť=Ʀ�=d{�=`��=��=$N�=?̀=:@P=�#=8��<X�<�   �   X4)<�+<��f<�<�u�<Fg$=��P=��y=�Ҍ=J��=y�=��v=�= &);�8Y��	���|�$�˾�y���S��������ֿx���=�����)#��*&�!/#���\n�~&����տ@ϯ�.�����P�5���žD�o������#����<�Vi=�`�=4Z�=F5�=X��=;��=��=0tc=z�-=���<X9�<��a<�   �   X���8������`{��@,�;�9�<�=ȟ<=bj=׎�=^i�=�,l=T�=�'�;jF=�����$k�)������G��Ä�����̿��ȟ����V�����(�����I�9{˿�:��R����E�y;��߹���_�9��h�����<�f=r�=�/�=z�=�#�=�V�=:�J=�"=�3�< ��:h�(�蓘��   �   �P���頽�̐�`Wk��M$� ��� S�9|l�<��=�K=T�c=��X=�M=У-<
����׽�P�(���g� �5��r����ew���`ۿ˭����u�y�����j��?����ۿIl��*����Nq��O4�2����X���F�"���$0¼<'�<ޛ^=���=tj�=�4�=$�b=��=��<P=ǻ,����E����x���   �   ��*���'�yn��+���ٽ�M����@�/�����;A�<g)=)9=��=���<�]��1"���-�ص��*�߾����EU��%���C��lÿhqِܿ𿈦���1��5��!|�goݿ7�ÿ�¦��M��9�T�,6���ݾy܏�h�&������X��m�<�aP=�Vu=�i=�h6=��<`�����?ꂽ#�½? ��/.�f�$��   �   �����㐾�����vq��*K�
����ȸ�����T��D��<D�
=��=@��<`� �6:t�z��/�m�)��/�}"4�1�g�c���W������>/Ͽ̖ڿ\�޿P9ۿEп�޾�a����
����h��4��&��R���j�O�`\� |� �<�L8=|�<=�d=@�R<�I����d�C�ɽ(��`�?�trh����ZG���   �   ��g�ᾀZԾ���.ˣ������J�T��p��@)"�Q��4��<��<H9�<�E;$;�JS����4������Ծ��v�<�p�i�F5��b0���-���絿�{������M������V�����k��>�����'־.đ��w4���F��PC<��<p�=��<П�;<�伤9���� ���=���}�E;��ss��.Ѿ��߾�   �   x&�h�#�3z�����H�>Ⱦmw���<e����f����n�`�2�@��<��<h�e<��Q�Կl�E�����T�����!�J-�l�7���Z��=z�Ĉ���������2��������|�]�]��W:�����㾁�����X�$ ��9q��J���<@�<��< ��;�1��n����T���Y������¾d��$p	�O��7�"��   �   ��c��1`��%T���@��A(�'W���޾�[��_j�������P����;x�<���<���;�ɼ@ו�0��&b�#�����پ@u	�y`%�FS>��+R��_���c�a-`��!T�?�@�5>(�LT�4�޾X��0Yj�\��철�H�鼰6�;��<荷<�v�;��ɼ�ܕ�8�#,b�����Y�پ�w	��c%��V>��/R��"_��   �   l���25��������|��]��Z:�������Ȉ����X�� �Cq��"J�X�<4�<D�<�˂;4�����6P���Y�����S¾���m	�����"�mt&�П#��v�b��@C�cȾhs���6e����z��bd�`b2�h��<x��<0�e<��Q�N�l�����{�T�����%��/�k�7��Z��Az�抉�Q����   �   K~��}����O��ő��?�����k���>���+־�Ƒ�p{4�����p� 7<h��<ƌ=8��<�߾;l���1���� �j�=�k�}��6��tn���Ѿ�߾"�律���TԾ����ƣ����2�J���h��^"�������<��<P9�< �E;�@��W���4����Ծ����<���i�7��j2���/��굿�   �   ��޿�;ۿZGп�྿B���z��I�h�,�4��(�0U����j��Q�� \����|�<N8=R�<=*k=`�R<�1��@�d���ɽF����?��jh��{���B�����Mߐ�:����nq��#K������彪�������)��<¯<>�
=F=,��<� ��?t������m�������$4���g�� ���Y��|���h1Ͽ�ڿ�   �   �2��7��3~�Tqݿ��ÿ|Ħ��N��VU��7�<�ݾFޏ���&����8�X�@k�<�bP=�Yu=��i=�o6=<.�< $����tႽ�½����'�Ǘ$���*�9�'�h�&��ٽ�D����@����� <0O�<�k)=�+9=��=�<Hc���$�� �-�^���N�߾p��|GU�'��E��	ÿ9sܿ֒𿧨���   �   f����k��A���ۿ�m��@���WPq�5Q4�\���kZ���F������6¼�$�< �^=�=l�=7�=��b=�=���<�ƻ�n���E�X���o���G��n࠽�Ð��Fk�4?$��ڥ� ��9�}�<��=�K=��c=��X=N=��-<`����׽5P�e���F�N�5���r�����x��6bۿN������u��   �   }������}���J�+|˿w;��������E�M<�+Ṿi�_�v�� ����<�f=��=�0�=	�=�%�=�Y�=ַJ=�*=�E�<���:X�(��|����������0ڈ��'�� w�;�I�<�=j�<=�fj={��=~j�= .l=��= #�;�G=����%k��)�����l�G�DĄ�e��]̿��R��T������   �   :+&��/#�h���n�'����տ�ϯ�������P����׾žY�o������%���<RVi=�`�=�Z�=6�=R��=���=��=xc=��-=���<D�< �a<�K)<(�+<��f<h�<�~�<\k$=~�P=x�y=�ӌ=*��=z�=j�v=r�=�%);D9Y��	��|�u�˾�y��S�2����I�ֿ���������])#��   �   �HP��-L��@�#5/��S�����ٿ�����y����=��� �z��h4����Pû �#=Ɋ="˧=���=�8�=��=��y= �A=��	=D��<0�6<C�;@�:��; p�;� t<���<�=��L=��z=ノ=1��=��=�hc=�V�<t���<����<?���������A��G��>ݮ��yۿt�������/�"�@�\2L��   �   �fL�KpH��%=�>?,�$��ا�ֿ<���5��\X:�����������/�諕�0���f�"=��=Qڢ=]x�=v|�=픉=��[=�4=H��<H�%<�O^�p��؋=��+�P�����x;��~<L?�<� /=��b=��=v��=�Y�=&�^=���<_��[���)|:�-⣾�@�=v=��䂿Sګ���׿^��P�},�t0=��gH��   �   �eA���=�(p3�l�#�T��y����˿ɡ�%8u�DQ0��I�l���D#�[(���z	�R�=�d=6��=�F�=�Ā=z�G=4��<�C<��(ż�����@�d�P���I�P�,�D����v��&;��<�e=�dP=��r=�v="�P=��<��H��Ӛ���,��\���=�%�2�|�w�����Ϳ�������#�y@3���=��   �   ��0���-�t�$����{R���㿕컿Q����s`�[� �u�׾�$��t���Sb��.�: =�ra=��r= �W=�=�Q�<@���V�
x�F���ҽ�2������4�۽�4��靌�:4� Ֆ� V�;(��<��)=D�E=��6=8��< ���[�����,
��g|۾�{"�8b��f��Wd���4�8O�8E$��-��   �   ����`�j��Ih�l��t˿�G��BŃ���E�I����Yc�:�>-��R�;��=��3=%=LC�<���:4T��)�iԽ7*�RQ2���M�Z�_�8�f��Tb��R��89�ܭ��罈˛��Y&���8u<��<��=�_�<��غII������i�`~��ͦ�q�F��<����ʿ� ����������   �   �(�>�����3/�w�ͿO��9�����`��'���~�����7�F��DV�Ȇ<��<���<��i<@�C��$H�������YL�a>��
��������xܾ�%`���ԯ��]��+���-DV��_��ս2�o�h��@N�;4ؤ<��< �H;�S
���~c;�u꛾�r��u'�1`��׎��*���̿��#������   �   ���6޿tBӿ����f5���p����l��8����+���,�r��\�8#��H���p%<���<���;���<�v����Zb6�D���ۦ���̾ �������HQ�L�������Ѿ���vA���"@�����춋� Nۼ ��9��><�ɽ;�H��놽-����r����� �6��j���G��������ѿa`ݿ�   �   %ܵ��	�������������~g��;����Ѿ`���a2�˽��x�������<`);�㫼"�~�=���'�G����o�þ#U��D����,��>?�8K���O�R=L�J#A��f/�f�����ʻȾ����ښO��)������м �i��=�;�E߻�J!��<���e0�oS��:KϾ�8�ڪ8�{d��P��������L���   �   ���Km���8���_o�,�Q���/�����;־b.��~�J��ｎ�j��D����:��;4Q��*�_�N�	oE��̕���ѾU
�l-�8�N��~l�(���Љ������o��6;��Cdo���Q���/�����?־�1��8�J����أj�4M�����:`�;�D��֬_��轫iE�ɕ��Ѿ�R
���,�B�N�=zl����HΉ��   �   O�O�9L�<A� c/�������0�Ⱦ���T�O��%�����@�м��h�=�;�a߻R!��B��2j0�xV��JOϾ";��8��~d�S�����������N���޵�2��@��坛�) ����g��";�S���Ѿ��qe2��������@���<�Y);�ҫ�2�~�(����G������þFO�������,��:?��3K��   �   �M��������󾄲Ѿ����=���@�����X���<ۼ h�9��><@½;tQ��#`��q�r�[����6�K�j�������e��M�ѿ0cݿ��Έ9޿Eӿ�����7���r����l�/8�i��񯼾�r�4_�+&����ps%< ��< +�;���z�v����[6�P��*צ�3�̾���j�/���   �   �־��Z���ϯ�DY�����=V�Z���ս"�o��S�����;�<��< tH;�X
�O���f;��웾"v�x'��3`��َ��,��̿���҄�����B*���#����1迊�Ϳ�P������"�`��'����j���n�7�I���[��<$%�<���<�j<��C�H������rRL�:��=������-��   �   �f��Lb���R�	29���������L&�h���/u< )�<D�=p`�<��غ�MI�����i�����]����F�����u�ʿ��<������	��*b����\i�M�dv˿I��Vƃ�G�E������\c��<��-��O�;��=��3=J%=�T�<�6�:�6��冽�^Խ�#�@J2��M�N�_��   �   Ғ����ű۽+��m�����3����Т�;�<N�)=��E=D�6=���< ��^��Ѷ����c~۾}"��9b��g���e�����;P�TF$�<�-�&�0���-�|�$�s��BS���㿩�.���u`�[� �ݧ׾�%�����Vb� !�:D=�ua=�r=nX=<=�f�<m�fG���w�����]�ҽ�'��   �   ~�P�<�I�`�,�����؆v�`�;�*�<�k=biP=.�r=*�v=�P=�~�<�H�n՚�A�,��]���?�/�2���w���~Ϳ���������#�QA3���=��fA���=��p3��#�ߓ�\����˿�ɡ�
9u��Q0��J�	����D#�)���	�,�=ff=���=I�=�ǀ=>�G=���<��C<��令�ļ���қ@��   �   �q=�X�+��O��@Ly;��~<�G�<@/=D�b=��=/��=VZ�=R�^=x��<�a������}:��⣾MA��v=�#傿�ګ�2�׿a^�OQ��},��0=�xhH�AgL��pH�&=��?,�h����kֿ|��!6���X:�;���ށ����/���� ����"=!�=ۢ=fy�=�}�=���=��[=�9=���<н%< �\����   �   ��: �;Pn�;h�s<��<N=��L=b�z=���=��=��=�hc=lU�<ܸ������=?�΄�����!A�H��[ݮ��yۿ�����ː/�,�@�a2L��HP��-L�׌@�5/��S������ٿ�����y��^�=�w� �B��h4����� û��#==Ɋ=H˧=���=�8�=�=��y=0�A=��	=P��<�6<�B�;�   �   Hq=�0�+� O�� Ny;8�~<0H�<�/=��b=�=x��=�Z�=t�^=���< ]�������{:��᣾�@��u=��䂿ګ�D�׿�]��P��|,�0=��gH�HfL��oH�/%=��>,��������ֿ����5���W:�����������/�l�������x�"=��=bۢ=�y�=�}�=���=�[=�9=���<�%< �\�����   �   x�P�*�I�0�,����x�v��;�+�<�l=:jP=L�r=��v=�P=Ȅ�<�H�Қ���,��[���<�p�2���w����Ϳ�������B�#��?3�§=�eA���=�So3���#����V����˿Jȡ��6u�>P0�`H�P���uB#��%��`<	��=2h=?��=^I�=�ǀ=��G=���<��C<��付�ļ���Л@��   �   Ȓ���𽩱۽�*��1����3��������;P�<ܗ)=ҴE=@�6=x��<��껀Y��p��	���z۾�z"��6b��e��8c���
�h�LN�+D$��-���0���-�]�$�����Q���I뻿=����q`�� �u�׾>#��V��JMb�@��:=xa=��r=dX=�=�g�<(l�DG�~�w�}���^�ҽ�'��   �   �f��Lb�|�R��19����:��w��J&����P7u<.�<Ի=�j�< �׺�BI�����0i�{|��~����F�x탿�����ʿ���������k��V���_�(�� g�\��r˿:F���Ã���E�����캾aVc�%5�t-����;"�=��3=(%=,W�< L�:�5���䆽�^Խ�#�AJ2��M�N�_��   �   �־��Z���ϯ�6Y��򼅾�<V��Y��ս��o��O�����;��<"�<��H;�L
����t`;�\蛾�o��s'��.`�d֎��(���̿�濎�����m'��������,�:�Ϳ&M��������`��'�������D�7��@���D꼐�<0/�<��< $j<��C�VH������kRL�:��<������-��   �   �M���������r�Ѿ����=���@�#���Y����6ۼ b�9��><�;9��Q憽��r�r�+
������6�ʺj�*��$���{����ѿ�]ݿ���3޿�?ӿ���3���n��T�l��8�T��թ��6�r� Y����������%<@��<�D�;����:�v�����[6�J��*צ�4�̾���k�/���   �   P�O�
9L�8A�c/��������Ⱦ鯕���O�?%�������м�mg��}�;߻4A!��6���a0��P���GϾ6�ާ8�|wd��N����������fI��iٵ�������������%{g��;�R���Ѿ9��]2�����P���İ�(�<@�);t̫�D�~������G������þFO�������,��:?��3K��   �   ���Km���8���_o�%�Q���/�����;־>.���J����"�j��:�����:�8;<2��:�_� �罖dE��ŕ���Ѿ�O
���,�z�N��ul�w���ˉ������j��|6���[o�'�Q��/����6־�*��ТJ�n��H�j�/��@B�:�";�;���_���oiE��ȕ���Ѿ�R
���,�E�N�Azl����JΉ��   �   &ܵ��	�������������~g��;�����Ѿ3��Ia2�R������ܰ���<`�);������~�V���N�G����þ�I�����7�,��6?��/K��O��4L�A�D_/��������,�Ⱦ�����O�� �a���H�м�Mf�`��;�߻�F!��;���e0�WS��.KϾ�8�ڪ8�{d��P��������L���   �   ���6޿rBӿ����c5���p����l��8�w�����Ür�\�b!��T����%<x��<�s�;�젼��v�����U6�����Ҧ�ں̾�������J�:��T��J�ݬѾ���9��F@�S������"ۼ ��9��>< �;�>���醽���{�r����� �6��j���I��������ѿc`ݿ�   �   �(�>�����2/�t�ͿO��6�����`��'����T���j�7��D��`M��<L2�<���<XAj<(�C��H�P���	�WKL��5������^���繾SѾ�)U��sʯ�\T�������5V��S�2�սH�o��8���ۻ;��<�&�<@�H;�O
���� c;�]꛾�r��u'�1`��׎��*���̿��&������   �   ����`�j��Hh�j��t˿�G��?Ń���E�>���hYc�9��-��z�;��=��3=�%=Lg�<���:���2܆�jTԽ��OC2�R�M�G�_���f��Db���R��*9�<��=��D���<&�����Yu< :�<|�=�m�<��׺FI������i�P~��˦�r�F��<����ʿ� ����������   �   ��0���-�v�$����{R���㿔컿O����s`�S� �_�׾�$����\Qb����:D=za=l�r=	X=�=l{�<0;��8�f�w����zҽ��t��������۽!��T�����3��������;��<
�)=&�E=Ҋ6=X��<����Z�����
��\|۾�{"�8b��f��Xd���4�:O�8E$��-��   �   �eA���=�)p3�m�#�T��x����˿ɡ� 8u�@Q0��I�X����C#��'�� V	���=Li=f��=+K�=(ʀ=ζG=|�<(
D<P,�l�ļ�����@�B�P�"�I�Ě,�����Xv�@[;`<�<Zs=�oP=Rs=|�v=ғP=��< �H��Қ���,�u\���=�%�2�}�w�����Ϳ�������#�z@3���=��   �   �fL�KpH��%=�>?,�&��ا�ֿ<���5��YX:�����������/�����Э���"=��=�ۢ=kz�=�=+��=��[=.>=L��< �%< &[�hm��U=��|+����@�y;h�~<�Q�<�/=�b=m�=���=�[�=v�^=ą�<�\��	���|:�&⣾�@�>v=��䂿Tګ���׿
^��P�},�t0=��gH��   �   G�|��w�{�g�dQ�T�6�� �6 �I̿�j��
d�]��JFɾ1�i���@�����<�5a= ��=ʚ=fL�=�E{=�B=`�=d�<� ;;0��H쀼 5��잍��9� �� ^:<���<Jn&=F�\=1��=�ڊ=�Ձ=��A=�Q}<���8��r��Pξ����g��q��ŉο?-��0��z7��Q���g�4$w��   �   iw�S r�@2c�0EM���3���������ȿd˙�� `�1��07ž�d���ܽ���|e�<�:[=�'�=���=�2�=�^=�6 =��<P!�;��#�ҵ��[��\�	�x��طμ��j� �E���<��=R�@=�o=��=��x=�?<=�|<Z�����Km� ʾ���pJc�߭��>˿I
��È�,64�-�M�xBc��r��   �   }�h�ad�ԉV��xB�̧*��_�C'�Lc��-%��HT�Rk�}r���U��~˽Zμ�H�<��H=4v=`�r=�|J=b=�W<h�������MK��p���}���梽坽������]�J��Xww��|�;x��<�+=��S=��W=��*=��v<����ڽMX]�V���B�� W�`�������(������*��gB�jJV�9�c��   �   7ES��RO���C��42�
���R�ݿ�;�������A�r��$��I>�M���i��4ե<��&=Bk:= @=\�<�]�r��"��]���d����y�8	� �$�.� ��y���B�ɽ�ύ�>@ �v/���[<�b�<��=�e= �a<��ټ�����D����������C�+�����%޿�&�r��<�1��C�=�N��   �   ��9�+�6�2"-�>\������ſ����c7m��\*��3�E��k7!�l���xy�x��<@}�<|��<`D�;|��,Ll�S˽�����>��f�}-��_���y��������>���Bl�ȟE�b��ڽC��,� ��� ��<��<`�.<��������B&�z���J���x+�:n�R㜿��ſ��c��|�PK,��86��   �   %:�·�^�������Ͽ�P��gE����I�ɰ����ԩl��?�B`���7� <<��%<00���+�3�������E��傾򘢾D��{�վ��e�a ��^ؾ�v¾;~��3����,M�2M�;㰽T</���>�@�;�I�; }��p�1����o��6����I��酿6����ͿPB�w�����E)��   �   o��l�������_��Eʿ�}���5���]���$�+��㝘�48�6h½�-"�����P�0�j���7��������l�k��I�ξ�m��$��v�!���+�6�/�N�,��#�r��k	 �ߣӾ�ԥ�,�s�Ƞ%��ɽ�aL��e��`G���-P�L&,�K"ƽ"$9�ߵ��=H��#�
�[�W��Gު�xGȿpF������6��   �   ŊֿJKӿe�ȿ<��ⵢ������`��;.�mO �����Fe�������2ݼ��>��3����;�~����Q&�V��/I��)��P�li5��?P���e�rms��x���t��g���R��58�(�?|��EY��FK���+���Ƚv�H��?���#[����K����9�x�c��m��u#��_,�5�]��p���Ѡ�tW��#Xǿ�iҿ�   �   m���*^��`������,�z�)vS��r*����ᦽ�h���W3 ��N��\6'��J��F����"��C���$�n�|�w���� �4�'�kP��w����3Ě����S���a��
��q�����z��yS�v*�=������4���67 ��S���;'��L��H@����"��=��y �#�|�>���ż ���'�gP�={w�e��t���(����   �   ґx�Ât�T�g���R��18�� ��v���T��H��G�+�O�ȽT�H��7���#[����y���d=���c�Tq��9(��b,���]��r��VԠ�=Z��"[ǿmҿ�ֿaNӿT�ȿ�>��I������`�b>.��Q �@��� Ke�r������6ݼ��>��(����;������L&�5���D��j��JM�qe5��;P��e�qhs��   �   �/�0�,�	#�޵�B �|�ӾoХ�0�s�y�%���ȽWL�Y��p2���1P�,+,��&ƽ�'9�����L羜�#�F�[�O���િJȿYI�����p8����������b�DHʿ����7��t]�Ư$�t��/���48��k½�0"�������`j���7����8��^l�af����ξ_g��~����!���+��   �   �^����Xؾq¾Ty������%M��G��ڰ�<0/�Х>� �;�U�;P}�8p������o�n9��
���I�U녿(���O�Ϳ�D������*��;�i�����]����Ͽ�R���F����I�f��6	��Ӭl��A���`�(�7��G< �%< 俻��7�������	E�SႾꓢ����U�վ����   �   ��������B:���:l���E�:��{ڽ�:��\�� ��,��<(	�<��.<���r���CE&�S�����辧z+��n��䜿ǂſ���d�"~��L,�p:6���9�ʿ6��#-��]�����w�ſӵ��V9m�n^*��5澣��9!�����y����< ��<���<0��;a���:l�XH˽1��!�>���f��(�������   �   g�$��� ���=���M�ɽ�ƍ�&2 ��H/�`�[<$o�<�=�g=��a<��ټ)����D�`�������C�3��Z��>'޿�'����{�1��C���N��FS�PTO�ԵC�62��L���ݿ�<�������A�H��%��\J>�pN���j���ץ<��&=Pp:=4G=h�< S\��������������s����   �   �ޢ�ݝ�5󋽾�]����Lw����;���<��+=��S=t�W=��*=��v<����ڽ�Y]�����*��WW�(�������S��;��d�*��hB��KV�e�c���h�}d�ЊV�yB�v�*�p`�(��c���%���HT��k�7s����U�o˽�ZμlJ�<��H=�v=
�r=ނJ=�i=��W<�V�Ի��Z?K�i���u���   �   ��	�����μ@rj� �?���<��=��@=� o=޽�=��x=�?<=��|<���s�� Mm��ʾ'��-Kc�W����˿�
��+���64���M�Cc��r��iw�� r��2c��EM��3�L��V�����ȿ�˙�`�f��r7žh�d��ܽ8���f�<�;[=m(�=̊�=4�=�_=^; =x�<S�;(�#�Xõ�,L���   �   P5��@����9�@��]:<p��<�m&=��\=��=wڊ=�Ձ=b�A= O}<�����	�r��Pξ���V�g��q���οQ-�1�{7��Q���g�;$w�G�|��w�n�g�TQ�@�6�x �$ ��H̿vj���d�2��Fɾ��i�r�⽰�����<R6a=-��=ʚ=L�=�E{=D�B=v�=��<�;;��X쀼�   �   ��	�����μ�qj� �?�l��<��=ֹ@=Z!o=)��=��x=�@<=ؒ|<@��t�콁Km��ʾ_��Jc������˿�	������54���M��Ac�Fr�ihw��r��1c��DM�J�3����O�����ȿ�ʙ� `����b6ž��d�)�ܽT�j�<�<[=�(�=���=/4�=_=t; =��< S�;@�#�dõ�8L���   �   �ޢ�ݝ�&󋽖�]�����Kw����;Ԑ�<H�+=��S= �W=<�*=@�v<���!ڽ&W]��������MW�ԣ�����D�������*�gB�hIV��c�N�h�7d�V��wB��*�=_�%&�_b��k$���FT�nj�2q��9�U��{˽8Qμ�P�<��H=�v=̟r=N�J=j=h�W<�V�Ի��b?K�i���u���   �   j�$��� ���"��� �ɽ�ƍ��1 ��E/���[<r�<,�=�j=Hb<��ټ������D�~�������C�Z����h$޿�%�}���1�=C���N��CS�^QO�$�C��32�	���ѓݿ�:������A�H��"���F>�cI���]��h�<��&=r:=NH=��< N\�Z������������s����   �   ��������=:���:l�x�E���{ڽr:����� )��D�<��<��.<���-����@&�ꌒ���Kw+�8n�✿eſ��b�j{��I,�*76�R�9���6�� -��Z�I���(�ſ���5m�&[*��0�M���4!� �����x��<Ȍ�<���<��;�_���:l�GH˽0��"�>���f��(�������   �   �^����Xؾ	q¾Gy�������%M��G�Cڰ�N./�К>��+�;���;��|�� p����4�o�-4��p�޾I�L腿v���Ϳ�?�������'�r8����������� Ͽ�N���C����I�֮�����l��<�ju`�(�7�x^<��%<�ѿ�"�ח��Ɣ��	E�QႾꓢ����Y�վ����   �   �/�.�,�#�ڵ�: �i�ӾWХ���s�%�%���ȽRTL��P��� ���P�\,��ƽ� 9�\����D���#��[����$ܪ�Eȿ�C⿷���.5�ƻ�ǹ�r����\�'CʿW{��4��W]���$�D��������7��a½<#"� t� �� Rj���7�M��
��Fl�\f����ξcg�������!���+��   �   ֑x�Ăt�P�g��R��18�� ��v���T���G��қ+��Ƚj�H��+����Z� ��ԋ��k6���c�~j����B\,���]��n��lϠ��T��:Uǿ�fҿ��ֿ)Hӿa�ȿ29��V������ي`��8.�M �s�+Ae�����8ݼ��>����H�;����8L&����D��g��KM�te5��;P���e�uhs��   �   p���*^��^��򧎿&�z�"vS��r*��������7����2 �M���0'�d:���-��,�"��6���7�|�N���=� ���'�KcP��vw����Ǿ��T�������I[�����_�����z�rS��o*����������^. �IG��0*'�\5���0����"�<�� ���|�-���¼ ���'�gP�A{w�h��w���*����   �   ǊֿKKӿc�ȿ<��޵�������`��;.�^O ���(Fe������p$ݼH�>�L��Б;�@|��hG&�w��;@�����J��a5�A7P�B�e�cs�Ìx��}t�}�g��R��-8�Z���p��;P��JD����+���Ƚ��H�T!��`�Z� ��"���R9��c��m��j#��_,�7�]��p���Ѡ�xW��&Xǿ�iҿ�   �   p��m�������_��Eʿ�}���5���]���$�
�羰���� 8�@f½�'"��v�@��h7j���7�u������G�k��a��U�ξa�������!���+���/��,�#�,��� �ØӾ�˥�r�s�^�%�_�Ƚ`HL�TA���฻P�� ,�� ƽ�#9�����,H��#�
�[�X��Iު�{GȿsF������6��   �   &:�·�^�����~��Ͽ�P��cE��~�I�������U�l��>�zz`� �7�He<`�%<������y���T���E�)݂�
�����J�վ?���W�x澕RؾRk¾0t�������M��A�BѰ�� /�Xu>��Z�;@��;��|�>p�~��U�o��6����I��酿7���	�ͿRB�y�����F)��   �    �9�-�6�2"-�=\������ſ����^7m��\*��3����6!�������x�x��<���<X��<���;|F��B*l�>˽
����>�{�f��$���؍��.����5��a2l���E����pڽ�1����� ��X�<D�<`�.<0������YB&�V���:���x+�=n�R㜿��ſ��c��|�PK,��86��   �   8ES��RO���C��42�
���P�ݿ�;�������A�i��$���H>��K���a����<��&=\v:=�N=\+�< �[�.��f��*~������gm�>��ȥ$�#� �������ʧɽ˽��x" ��/� �[<���<<�=�m=b<H�ټ`��)�D����������C�,�����%޿�&�r��=�1��C�>�N��   �   }�h�ad�ՉV��xB�̧*��_�C'�Lc��+%��HT�Mk�jr��֛U��}˽UμP�<ֆH=nv=ܣr=ވJ=Pq=(X<�+�����j1K��a���m���֢��ԝ�V닽�]����@w���;���<��+=��S=J�W=D�*=��v<H��ڽX]�I���A�� W�b�������(������*��gB�jJV�:�c��   �   iw�T r�A2c�1EM�3���������ȿd˙�� `�/��(7ž�d�~�ܽ��<i�<6=[=G)�=鋒=x5�=~_=�? =�%�<`��;�x#�д���<����	���t�μ�Uj� <9����<��=ܽ@=�$o=a��=f�x=2B<=��|<&������Km�ʾ���pJc�߭��>˿J
��È�,64�,�M�wBc��r��   �   Z���^���|���,t��!S�/�1�x��F鿸s��JÃ��7�d(�d�����:�T���;T�1=��{=V߇=��|=.+O=�=�>�<��:�Cf�`׼�t��]�d
�$��\������xff<�}�<2�;=0Ji=��{=�g=�Z=��#;�k��*�j���.��N�9�E���������V`�7 3��T�H�t�N����c���   �   ����,��О���]o�lMO���.���`�応��|��\�3����
���q���N�`��;� += +o=@e}=�0d=v�/=|��<0D�;(/@���鼞�+�:�O���]�ȦT���4�`b�`}�`q3;m�<�*=�P=ܞi=�[[=V=@�;��d�ʈ�����c��2b6�e�� t�������`�/�pP�@�o������&���   �   �1���,��{���a�iD��8&�<��:�ڿ�᧿��u��)�H�۾"Z�����w>����;�p=�8I=<7E=4_=x.�< uV���⼼�S��*���t��g�н�|ٽY5ӽ�^�������Pd�����xk<F�=@�1=t�5=�"=@<�:B�R�T�������߾c?,�idx��m���\ܿ^�	��&���D��a���z�����   �   C�v�%�q�Lc�4�M�� 4��������ɿPM����`�Z��gǾv�i�����-'��כ;p��<J�=`��<�-�;� ��(�]��S���p��^A��
5�6GE��gK���F� �7��) �x��.d��l�r��lݼ J9Š<�y�<y�< ��9H�9�p���:Do�x	ʾ�r���b��K��.�ʿ�d�����3���L��b�7qq��   �   �W��,S��bG�ߏ5�b����������\Ո��!F��Z�����r�H��rȽb����:��`< �<81�ҽ-��z��5k��v8��j�h�������9q�� ӭ��c���u��t���o��?>��+�+|���TB�0n}� ޓ;�9<�Z��#�>SнϦL�踮�x��4G�hD���ܳ�����1�16��4�8fF�4�R��   �   ,�6�7�3�fO*�b���
�/:��¿�l����i���'��������#�:��(����� �λ�ȼ�q��ܽ��+���q��ŝ������0�>��[m�#�	�m�I��X3徂6žH8���px�f�1��G置9��01�Pk"� �*�Lj�V�ܫ&�8X��#�(�6�i�/��w¿Q�꿰	�d���=)�S�2��   �   �v��#����!3�����Tſ�/��DP�d�?�~ �������a��^���o|�P�h⟼h	�������F��������~������#*��<�~�G��L�u�H�՞=��,�2��^����lľZg��L�K���
A��4��`���$��G򁽉� ���b��������>�
�}�����R�ÿӴ俌��������   �   ����q��L�'�ҿ�Q��𤞿ڒ��NAJ�b�2�Ҿp���U(��R����@�����������>���hN�lX��g1׾�r���0�I�R� q�����HN��L.��i݌�ׇ���s�vxU��63���m�ھ	$��w�R����㑽8� ��;���D��Һ�,�'��щ�MPѾ��NuH�aI��I���Y����пx�����   �   �)��p6���Ҳ��ƣ�UY��}Ot���E����{�߾eF���F�����1�r��hw���{�Fy�v�C�[n���%ݾ����sC��Qq�֯��_&��)����z��-���9���ղ�Nɣ��[���St�X�E������߾�I���F�P���7����:t���{��r�c�C��j��!ݾ����oC�QMq�>����#�����w���   �   q+���ڌ�-�����s�tU�133�֢���ھM ���R�.��lޑ��� ��;��HD��׺��'�qԉ�]TѾ����xH�~K�������[��пע�s�"����� P�1�ҿkT��F���Δ��sDJ��!�ĭҾ쁊��X(�oV��^�@�L���Ά� ��w6���bN�\T��$,׾vo���0�ǿR��q�ւ��vK���   �   L�ʜH�h�=��,����;���ugľ\c��9�K����;�����\(&����0� �>�b��������>���}����ÿʷ�3��������x��%�c���4����MWſ�1���S��?�\"�������a��b��Zs|��N�$ٟ�H_	�;���e��_
F�~������zx������*�:<���G��   �   i�	���B��-��0ž�3���hx�2�1��>��2�����U"�@�*�Jl�e�����&�hZ��P&�E(��i� ���¿���.	���n?)�T�2�6�6�/�3�6Q*����

��<���¿1n��-�i���'��㾶����#�!�����p���bλ4�Ǽ�q���ܽ�+�h�q���������*�<����i��   �   �ͭ�e^���p�������o��8>��%��r���FB�@E}���;�H<��Y�L&�^Vн��L�����y��6G��E���޳����53��7�̎4�hF�?�R��W��.S��dG�k�5����ɠ����y���vֈ�P#F�\�����^�H��tȽ�� #:��`< <��0���-�q��(e�Bo8�wj����������k���   �   X`K�f�F�#�7��# ����|Z��`{r�\Sݼ �S9dӠ<<��<�}�< ��9�9�N����Fo�Sʾ:t�b�b��L����ʿef��� �d�3�:�L�՗b�sq�3�v���q��Mc���M��4�������ɿ2N����`�O���Ǿ�i�2�콜.'���;X��<��=���< ��;l��X�]��I��0e���:��5��?E��   �   �sٽE,ӽV���Bd�������p>k<r�=��1=@�5=$=�-�:��R�������?�߾j@,��ex�yn���]ܿ	�	�Q�&���D��a��z����o2���-��C{���a��iD��9&������ڿm⧿��u���)�  ܾ�Z����� x>�P��;�r=Z<I=v<E=f=�?�< �U����>�S��"���k��9�н�   �   ��]�:�T���4��Z��E}� �3;tv�<h.=��P=Ҡi=�\[=�=�|;��d����.���N���b6�����t��&��z����/�P���o���.'��|���)-��$���-^o��MO�3�.�;��������C|����3������q���N�P��;�+=-o=�g}= 4d=ʑ/=���<Pu�; @���@�+�z�O��   �   �]��
����܅�����@ef<0}�<��;=�Ii=b�{=��g=FZ=`�#;�k�+�����~���9�c��������k`�N 3��T�^�t�V����c��Z���^���|���,t��!S��1�c��F鿔s��+Ã�k7�(�+�����X�T� $�;Ώ1=`�{=~߇= �|=f+O=.�= ?�<��:`Cf�0׼�t��   �   �]�@�T���4��Z�xE}���3;�v�<�.=�P=Z�i=�][=�=@�;ȵd�w��V������a6�7���s��'������/�P���o�5���]&������\,��l����\o��LO�r�.��������{����3��~�F
���p���N� ��;$+=�-o=dh}=n4d=�/=��<`u�; @���L�+���O��   �   �sٽH,ӽV��zBd��������@k<"�=��1=��5=n&=���:�R�_������߾�>,�}cx��l���[ܿܽ	���&���D�Ѳa�p�z����0��,���{���a�hD�8&����0�ڿ�৿S�u��)���۾Y��~���r>����;u=�=I=R=E=�f=�@�< �U�h��@�S��"���k��C�н�   �   _`K�j�F�!�7��# ����UZ���zr��Qݼ �T9P֠<���<d��< 6�98}9�n���9Bo�ʾ�q�6�b��J���ʿ.c������3�L�L�k�b�`oq�T�v�B�q�XJc���M���3���������ɿ.L����`���{ Ǿ��i�{��&''�`	�;x��<��=��<P��;���&�]��I��3e���:��5��?E��   �   �ͭ�g^���p�������o�p8>��%��r���EB�8>}�`)�;@X<��Y�
�aOнC�L�#����v�3G�FC��z۳�ʉ��0��4���4�idF�6�R�pW��*S�aG�7�5���������l���Ԉ��F�_Y�Î��8�H��mȽ"����: �`<<@�0�ܭ-��p��e�Bo8�wj����������k���   �   k�	���B���,��0žu3���hx���1��=��1���鼈D"��x*�4b�����&�<V��X �)(���i�����¿���N	�ʿ��;)�\�2�!�6�5�3��M*����3
��7���¿�j��٣i���'��㾜��	�#�������0��0Cλ@�Ǽ��q�W�ܽ�+�`�q���������!*�A����i��   �   L�̜H�g�=��,����+���_gľ>c���K����9������഼���W큽|� ��b�������>���}������ÿ���
���Ҍ��t��!����x1���NRſ�-���L��?�F�����a��W��Td|��:�`̟�L[	�������.
F�s������|x�����*�=<���G��   �   t+���ڌ�,�����s�tU�*33�̢�h�ھ( ����R����Zܑ�\� �,(���D��̺�0�'��Ή��LѾ���"rH�mG����jV���п1��s� �����lI���ҿ�N��n��������=J����ҾV|���P(��K���@�P���������O5��GbN�GT��,׾uo���0�ʿR�q�؂��yK���   �   �)��p6���Ҳ��ƣ�SY��vOt���E����[�߾5F��� F�Պ�*,����j���{�!k�j�C�lg���ݾ���-lC�Iq�ƪ��� ��|���t���&��63��yϲ��ã��V���Jt���E������߾�B����E�7��|$����k�.�{��p��C��j��!ݾ����oC�TMq�@����#�����w���   �   ����q��L�%�ҿ�Q��줞�Ւ��DAJ�U�	�Ҿ/���T(�RP��&�@�����|�_����-���\N��P��4'׾`l���0�w�R�$q�2����H���(���׌�t����s��oU�9/3����"�ھ����R�L���֑�N� ��$��bD��к�w�'�[щ�4PѾ���LuH�bI��L���Y����п|�����   �   �v��#���� 3�����Tſ�/��=P�Z�?�m �������a��\���i|��<��ş��S	�믋�����F�v������br��n���*��<�)�G�RL��H��=��,�פ�����bľ�^��U�K�3���2������״����&�� �n�b��������>��}�����U�ÿִ俍��������   �   ,�6�8�3�fO*�b���
�,:�
�¿�l����i���'��㾾����#��������P��@λh�Ǽ��q��ܽ��+���q�𻝾S����#�[���
f���	��;��w&�+žw.��[`x�Y�1��3�G*�����)"�Hl*��b��什�&�X��#�(�8�i�0��y¿S�꿱	�f���=)�T�2��   �   �W��,S��bG�ߏ5�a����������ZՈ��!F��Z�ϐ��؍H��pȽx����:ha< :<��0���-��g��\_�Fh8��nj����s���tf��'ȭ��X���k�����B�o�1>����h��L6B��}�0i�;l<�{Y���]Qн?�L�¸��x��4G�iD���ܳ�����1�26�!�4�:fF�6�R��   �   D�v�%�q�Lc�4�M�� 4��������ɿMM��|�`�Q��IǾ�i�9�콘)'�P
�;`��<��=P��<pا;볼(�]�@���Y���4���4�s8E��XK��F��7�� ����(P���ir�@6ݼ �_9��<��<0��< ��9
~9�����Co�`	ʾ�r���b��K��1�ʿ�d�����3���L��b�8qq��   �   �1���,��{���a�iD��8&�<��:�ڿ�᧿��u��)�8�۾Z������t>����;^v=�@I=�AE=�l=�P�< (U�P��@�S����>c��,�нmjٽ#ӽ/M���朽�3d���H���ck<$�=�1=��5=�(= ��:��R���������߾b?,�jdx��m���\ܿ_�	���&���D��a���z�����   �   ����,��О���]o�kMO���.���a�忛��|��X�3����
��Lq���N�`��;~+=/o=lj}=L7d=��/=���<��;��?���$�+���O��]�b�T��4��R��(}�@24;���< 3=��P=$�i=�_[=<=@�;��d��������^��2b6�f��!t�������`�/�pP�?�o������&���   �   ���
ߧ�l��d���u�m� 6F�D�!��	��ǿܒ�2sM���j���(�/����� S��2�	=4Z=�p=<�[=�,*=(��<@�;�hB��/� �)�,�L�2�Y�|P���/�<���hpj� �w; [�<r=��O=h�c=֞M=�C�<���ꗘ�
84�7x������O��g����ȿ�/��#��qG���n�f	���4������   �   ���^������͇��i�#�B�6�>���d�ÿ�Z��7�I�{O�c5����+�2w���h���w=8�L=f0\=�@=�=(hp<�H��$~ռV$5�~Sp�6v��*���P$����v�r�=��8꼐���@<���<��4=��O=�I@=�\�<8k��$��8=0���:��L�<Α�,�ſ� �U ���C�*�i�z��몘�D���   �   ���,E��7ڎ��%��
\��8�p�����O�������>�P���@���� ��N��p"ϻ���<(�#=<!=0��<Pz�;얌��N3�!K��Lc��9��|�������G ��C齕DĽ�����?�@v��`�;P4�<ȷ=<G=���<h��8|����$���\���n�@��?��ŷ�����bR�O]9��T\�d������"���   �   2X���K���t���f��H���)����*߿�i���'{�+.�eU⾶�������~n����Ę�<�3�<�HT<`��ď�Gg�����h,�L*9�rCT���e�=nl�{g��tV��<�Җ���齖���6�(�0:���!<<�<��a<p�8�^R{�=~�������-�/�L�|�/P����	��)�_H��Cf���<���   �   CHr��m�Jo_��kJ�qy1���?���$ǿ�A����]�*��5�ľ59j�07��ܲR��+Q� ��:`�|�@Bм.>v�f�ֽ� �g�X�뇾稠��c��k<��S�ž�¾�ϵ�F�������]�`�$�)�޽@��� �`Sܻ@���P|��]�/ ���dm���ƾ����^�3���<ǿ�Y��r��5�0��iI��o^���l��   �   N�K�r#H�'Q=�%�,�����|�Ф׿Hh��1L��LL<�� �U;��ĀA�3�̽�U<�4꫼�Z���s$�+���|K�m���δ�Ηܾ ��N�>�����/�8D�_�8Z߾u�������L�O���
��Ħ���/��]���/��t E���н`�C��B��� �"�<��C�������ֿ�����/�+�ZB<�.G��   �   (�'�(!%�����x���K3ڿ�γ�Z��4DV��V�8Ͼ�Â����1���H72�0���0L�Ah�����g����\۾�T
� 3&�m?���R��_��&d�c:`��T���@�P(�v�<s޾�7����k�i��ù���T����s8��B�����%���Ͼ��U�U��p������ÞؿH�����6��@�$��   �   M;��'��J�����Wο.⯿���o�a�X�(�>���ߞ���E��
�$_����9�||\�t"��F��^�p���NA�����TF�`�k�{z������.�����܈���w������F#n��H�x_!��1���+����s����۝��n�a��y=����tm�d~E��U��Mq��'�$``������\��/N̿
�濣���d���   �   ��ӿaGп��ſ�|��/?��z����]���+�����~$���Bf�H��:���jaW���V�ḷ����cd�ꫮ�������)���Z�:��������0�ĿҚϿ>�ӿ�JпP�ſ����A�������]�%�+�����(���Gf�e������bW�F�V�ȣ�J��r]d�����g����)���Z�����ο��� ��оĿM�Ͽ�   �   ���ʅ���t��똇�{n��~H�\!��,���'����s��������z�a��y=�k����r潪�E�Y���u��'��c`�����_��IQ̿z��Z���X��G=��)�,N����M ο�䯿�!����a��(�0�➾��E��潃`����9��u\�T���|���p�9찾~;�����OF�m�k��w��������   �   �!d�C5`�	T�~�@�X�'���m޾3����k�4d������T�����t8��E�����o'��#Ͼe���U��r��d�����ؿ����޿�<��f�$�X�'�E#%�����������5ڿѳ�#���FV��X�#Ͼ�ł����
����62�(��"'L��`���	���g�[���+V۾xQ
��.&��?���R��{_��   �   ���'	�c@��[�T߾/���R���r�O���
������/�R���+���E�S�нn�C�1E���� ���<�oE�������ֿn������+��D<���G���K��%H�AS=���,�E��5~��׿�i���M��SN<��� �@=��
�A�^�̽�U<�,㫼�K��(h$��"��t�<K�����ɴ�r�ܾ� �K�/���   �   @�ž�����ɵ����	���]���$��޽[8����pܻ����{���]�����gm���ƾ.��X�^������=ǿ�[��ά�ڹ0��kI�8r^�+�l��Jr�h�m�lq_��mJ��z1���+����ǿ�B����]�y����ľV;j�M9����R��"Q�@��:�|�|)м�-v���ֽ6| �\�X�t懾�����]��m6���   �   �el�Wg��lV��<���������.�(��9��"<p"�<��a<��8�@U{���L���(�侤�/�D�|�rQ��n�
�$�)��`H�vEf���c��^Y��M���u����f�^�H���)���,߿�j���({�:.��V⾖�������n����\��<@�< lT<p��Ȁ�
^����&�#9��;T�V�e��   �   ����B �$:��;Ľ���r�?�P`��P[�;�A�<��=JJ=4Ŀ<X���}����$���������@�z@��������!S�@^9�V\�������l#�����F���ڎ�3'��\���8����x��O��K��7�>�>���ҋ���� �	O��ϻ���<:�#=�&=`��<���;����@3�$C��fZ�����Z����   �   U�������v�H�=�4*꼰��H3@<���<��4=�O=8K@=�]�< n��%��>0�������L��Α���ſ� �~U �@�C���i����g������;�����j����͇�i�z�B�H6�������ÿ�Z��y�I��O��5����+�w��b��y=X�L=T3\=��@=��=�~p<����nռ�5�RJp�gq���   �   <�Y��P���/�����pqj���w;lZ�<=(�O=��c=`�M=�B�<���o���j84�xx����K�O��g����ȿ�/��#��qG���n�s	���4��������ߧ�b��W���Y�m�6F�.�!��	��ǿ�ے��rM����*���ϊ/�v����M��Ɗ	=�Z=Np=��[=�,*=���<@�;�gB�X/���)��L��   �   \��������v�<�=�*�H���3@<@��<��4=��O=L@=8`�<�e�$���<0������L�Α��ſp ��T �U�C���i�&�������
��?���������*͇��i���B��5�������ÿ<Z����I��N��4����+��u��`R��Rz=&�L=�3\=@�@=ʽ=pp<����nռ�5�^Jp�lq���   �   ����B �%:��;Ľ���<�?��_���^�;$C�<��=�K=<ɿ<Ц�z����$�Q��Y�����@�9?�����؂��Q��\9��S\�������!�����GD��cَ��$��	\�7�8����|��*N����h�>��������\� � L�� �λd��<��#=�'=t��<���;H���@3�)C��mZ�����l����   �   �el�^g��lV��<������齋���~�(�(�9��"<�&�<�b<�8��L{��|�޼������/���|�0O����D��)��]H��Af�	����W���J��{s��I�f���H�ϫ)�+��;)߿�h���%{��.�GS�3�������wn������<0D�<qT<x��\���]��ۍ�&� #9��;T�`�e��   �   I�ž�����ɵ����		���]�޹$���޽�7����� ܻ@���X�{���]������am���ƾ!��2�^�����z:ǿ�W��=����0��gI��m^�U�l��Er���m�m_��iJ��w1�v����Vǿ4@����]�y����ľ�5j��1���R��	Q���: �{��&м�,v�y�ֽ.| �^�X�w懾�����]��u6���   �   ���)	�e@��[� T߾%���C���=�O�p�
������/��H�������D��н9�C��@���� ��<�{B�����r�ֿ���R��^�+�B@<��|G��K�!H��N=�7�,����{�p�׿Sf���J���I<�B� ��8���|A�>�̽@K<��ի�@C���e$�
"��<�K�����ɴ�v�ܾ� �#K�4���   �   �!d�F5`�	T�|�@�U�'���m޾�2����k��c�����*�T����j8��=������"��mϾ����U��n��ŷ��#�ؿ8���H��B��&�$���'� %���)��0���s0ڿ~̳�\��AV�T��Ͼ�������܊���+2�<���"L�l_��-	���g�Q���&V۾yQ
��.&��?���R��{_��   �   ���̅���t��阇�wn��~H�\!�w,��f'����s�,��������a�8o=��}���f�	zE��R��6m��'��\`�����dZ��@K̿������z��U9��%��F��F��:οr߯�`����a�R�(����qܞ���E�)潴X��z�9�"o\�J���{�_�p�$찾v;�����OF�p�k��w��������   �   ��ӿcGп �ſ�|��.?��w����]��+�����O$��2Bf�P��+����WW�X�V�����?���Wd�C���}�����)���Z�g������������Ŀ֓Ͽ#�ӿ�Cп��ſ{y��T<�������]���+�P���^ ���<f���������TW��V�%ţ�f���\d�ӧ��X����)���Z�����ѿ��� ��ԾĿP�Ͽ�   �   O;��'��J�����Vο,⯿���f�a�J�(��ߞ��E�7�[��2�9�j\����w�Z�p�谾6���~��KF���k�u��!�������������q��%���{n��zH�eX!��&���"����s��������}a�bm=��~���j潤}E��U��2q��'�#``������\��1N̿�濦���f���   �   *�'�(!%�����u���H3ڿ�γ�V��+DV�qV�ϾIÂ���������,2�Ώ��L��X��L�ͯg�镤��P۾N
��*&�o?�γR��v_�Td�0`�&T��@�8�'�~��g޾C.��L�k�b^������T����fi8��?������$��dϾ��R�U��p������ĞؿJ���	��8��C�$��   �   P�K�s#H�'Q=�#�,�����|�Τ׿Fh��.L��BL<��� �;���A�z�̽JM<��ѫ�`7��J[$�x�� �M�J����JĴ�R�ܾw �UG�.������<��W��M߾���������}O���
�ȳ��:�/�P:�����$�D�K�н��C��B��� ��<��C�������ֿ����1�+�\B<�/G��   �   DHr��m�Jo_��kJ�qy1���?���"ǿ�A����]����ľ�8j�5����R�@Q����: g{�мDv�[�ֽ�u ���X��ᇾ����7X���0��5�ž����6ĵ�Ԁ��U���]�#�$���޽g/�����0�ۻ�֒� �{���]�'���dm�z�ƾy���^�6���<ǿ�Y��s��6�0��iI��o^���l��   �   2X���K���t���f��H���)����*߿�i��~'{�%.�HU����3��dzn�P��@��<�N�<`�T<0^�Tr�+U��>����9��3T�B�e��]l�!
g� eV��<������4���^{(�У9�H,"<\3�<�b<��8��M{��}�������)�/�N�|�2P����	��)�_H��Cf���<���   �   ���,E��7ڎ��%��
\��8�p�����O�������>�>���!����� �UM��`�λ4��<Д#=�,=���<@�;di���33��;���Q��,��n���h���= �n0��2Ľ����D�?�H��p��;\R�<v�=�O=Pο<����z��3�$����O���l�@��?��Ʒ�����dR�P]9��T\�f������"���   �   ���^������͇��i�#�B�	6�>���d�ÿ�Z��5�I�xO�U5��V�+�zv���W���z=r�L=�5\=R�@=��=��p< ύP`ռ�5�fAp��l��{��������v���=�x����@K@<���<�4=��O=:N@=8c�<�b��#��=0���7��L�;Α�-�ſ� �U ���C�)�i�z��몘�D���   �   :=��������9&������)kV�.��i
��տ&���;^�����ó�IE�錭�y��C�<A=nxX=8C=t�= �<@0����f���X�|�ℽn~~�к[���$����`�z�8c�<�=�<=��Q= :=TN�<�2��]t��
%H�o���*�C�_��E���׿�G�W/�ScW�����g��ɫ������   �   �������j̧��Д���}��xR��+��.�>-ҿx���AZ�;��'��T�@�1��(�{��[�<R�2=(bC=�t&=H��<@��;h8{�
���e������Υ�����ܦ�8����Zj�6��,5��@T�;p��<�n=�i<=��+= ��<� ��c̮���C����(C���[�煜��ӿz����+�vLS��l~�{���m֧����   �   O����}��鿜� f��h�n�#DG���"�����ȿ$�����N�k��Կ��)5�
������@��<l=�=���<�>ͺt��B�d��5��`/޽lU�s��0����z��D�uʮ��5l�8$�l`�d�<H%�<�c =l5�<�2��������7��q��		�pP�����|ɿ�J��J#��G�t!o��^��R����a���   �   ���Ql���V���{�m�X��o6�L���4ￃ!��c��*�<�z��������#������v���}
<x�l<pp�;�9��t�J��A��FF��*�|�N�F�k��H~�B�����m�?�P��,�Z��tĶ��aS�,��@�,;��P<p��;�բ�X핽cS%�#������4�=������ʸ�j��+�8y6�b�X�Y�z���9���   �   l���J��>�r��Z�Z�>���!����\gտW����Uo�{�%��J׾t���K!��҂����������Z�"��KF��d����4���p���u^��obžӾ��׾��Ӿ[ƾޤ��a��r�s�њ7�M\��B����� kv��Z�d�Ƽo0��h���̂�y~ؾOH&�Cp�
���ӈտt��n�!��T>�h�Y��q��
���   �   �W\�9X�7L� �9�^�#����'�� 鷿�@��݉K����4��p�W�q:콤m��> ��/��*�T�鞽����ib�l����$ƾ���_e�*���F$���'�ݤ$��,��C����Ⱦ�C��x\e������ �[�D�����lr�D��Y��Ŵ� �+�K�;��b���<P�e#���"���8��3K�H�W��   �   tW4�M1�V"(�A��Aa�~����ԯ��Mg��&�;��D����+�� ����a�l�9��~���ҽ,�*������ʹ�{�Qk�X34��N��c�(q�8�u�J�q�c�d���O��y5�����|����ꁾ'�,�0ֽe���pA>��_e�o�½�,�SY����ᾤ�%� �f��7���꿿&Q���q(��e'���0��   �   ���`�����������ܿ�u���Ú�xWs��T6�'��4��º[��B��K����h�� ���ӽ��+�u8������R��-�H�V�|~��ᐿF�������ᪿ���i��ϲ������X��c.���?oþNO��,k-��=ս�����(k�4��mc��[����+;�g�5�8r�(FX��:ۿ�m�����u5��   �   ���A߿�ӿ(j¿�֫�����n��K9�E0	��T��F+~��{�-���t����r����@����|��V��Wm��08���l���������U���ӿS�޿j���߿��ӿgm¿�٫�+���n�RO9��2	��X���0~�H�����D���"q��쿽N����|�~R��~j��,8��l���о���R���ӿ��޿�   �   rު��	���e������:��FX�3`.����jþL���f-�/8ս���Z(k����,f���[�w����=���5�<r���*[��j=ۿKq������7����u�����0�����ܿ�x���Ś�([s��W6�F��(����[��D�,M����h���9ӽ��+��4�����6	�-���V��v~��ސ����ǫ���   �   ��u�՛q�3�d��O��u5�Q��!������]灾�,�)ֽ ����=>��`e���½��,��[�����4�%�_�f��9��E�,T迣��o*�h'���0��Y4�tO1�}$(�* ��b���u�������Gg�3&�]��S��<�+��"��J�a� �9�j�}���ҽs�*������ȴ��tﾊg��.4��N���c��q��   �   W�'���$��(��?�o��+�Ǿ�>��#Ue�M�o���"w[�������nr����KY�cȴ� ���K��<��|����R��$���"���8�U6K��W��Z\��;X��	L��9��#�"��l���귿mB��	�K�4��D���W��<��m�F; ������T�������ab������ƾ���a�}�?B$��   �   1�׾9�ӾUƾ\���:\��$�s���7�|Q��������HKv�XI���Ƽ�1��8��$΂���ؾJ&��p�����Ɗտ����!�|V>���Y���q� �����)L����r��Z� �>��!�����hտ�����Wo��%�qL׾����s"�ӂ�	��@`���cZ����c=���X��w�4���p���X��Q\ž��Ҿ�   �   �{��`	�n	m���P���,����	����RS�0���N-;�Q<0��;�բ��U%����͕��è=������˸���7��z6��X�m�z�C��b:������m���W���{���X��p6�'��J6ￋ"���c��L�<���������#�]����s����
<�m<���;� ��v�J�
8��Z@��*���N��k��?~��   �   -+�0��u�v;�6®��'l��� �_���<�/�<$g =48�<�3��⒤��7�s���	��P������ɿhK��K#��G��"o��_��F����b��S����~�������f����n��DG���"�n��2ȿ������N����q����5�R��l������<dp=�=�ǝ<��˺���p�d�X-���%޽BP��m��   �   ����צ�x����Qj�r���'����;��<Fr=l<=&�+=���< "��hͮ���C�I���C���[�d�����ӿ����+�MS��m~������֧�����)��;����̧�Dє��}�AyR��+��.��-ҿGx��BZ�h�0(��x�@�����{��^�<��2=DeC=�x&=H	�<0��;�{��|���d������ɥ��   �   ℽ�~~���[�8�$�����z��b�<��=j<=.�Q=�:=M�<X4���t��p%H�����Z��_��E���׿�G�r/�qcW����h��#ɫ�����:=��쵸�����+&������kV��.��i
�ʦտ�%��Z;^����\ó��E�a��� y��D�<�A=�xX=�C=Ɠ=��<@,�0��2���X�|��   �   ����צ�y����Qj�j���'����;���<�r=�l<= �+=d��<����ˮ�A�C�K���B���[������ӿG��Q�+�LS�'l~�����է�s�����+����˧�nД���}�DxR�.+�M.��,ҿ�w��AZ���7'��2�@�t��(z{�pa�<h�2=�eC=(y&=�	�<���;�{��|���d������ɥ��   �   7+�7��u�v;�/®��'l�T��_� �<�1�<�h =d=�<�+��������7�1q���
	��P�:����ɿOJ�6J#�<�G�T o�$^��s����`��L����|������/e���n�CG�5�"�\���ȿ]���ɱN��������Y5�2��t������<�q=
�=ɝ<@�˺@��n�d�Y-���%޽JP��m��   �   �{��h	�s	m���P���,����ۺ��8RS�\�� f-;�Q<0��;tʢ�tꕽ�Q%���������=������ɸ���M�x6��X�u�z��
���7��@��k���U���
{���X�an6�F��S3�2 ��
b����<�8�������> #�񑽠h����
<Xm<0Ƒ;���J��7��V@��*���N��k�@~��   �   <�׾@�ӾUƾ\���7\���s��7�!Q��x���X��X@v�8�,�Ƽ�,��,��˂�j|ؾ�F&�F p�����*�տh���!�S>�\�Y���q�?	����iI���}r���Z���>�A�!�ǡ�neտˬ��[So���%��G׾����o��͂������>��0YZ�V���<��WX��l�4���p���X��[\ž��Ҿ�   �   [�'���$��(��?�k��$�Ǿ�>���Te��~���(t[�J�Z���cr��
Y�~ô������K��9�������M�"� �"���8��1K���W�DU\�n6X��L�ݪ9���#�9�����緿P?��G�K����j��Z�W�!4콤m�4 ������T�:�������ab������ƾ���a�
}�CB$��   �   ��u�ڛq�7�d��O��u5�N���񾪉��9灾x�,��'ֽĨ��l6>�BUe���½`�,��V�����_�%���f��5��^迿ZN�=���&��c'�@�0�U4��J1�  (�@��~_�{鿍��������g�b&�b��w����+�����va�ؿ9���}�U�ҽ�*������ȴ��tﾊg��.4�	�N���c��q��   �   tު��	���e������9��AX�-`.����jþ�K��f-��5ս}���dk�b����_�v�[�ۣ���8���5�a4r��왿�U���6ۿj�����e3�i��F���~�����4�ܿ�r��%���hSs��Q6����� ��j�[��>��D����h����ӽ��+��4������0	�-���V��v~��ސ�"���ʫ���   �   ���D߿�ӿ)j¿�֫�����n��K9�80	��T���*~��z����|���Xk��_忽����|��N���g��)8��l����𻪿iO��|ӿ�޿ؤ⿂߿y�ӿ�f¿�ӫ� ��5n�DH9�a-	��P���$~�w�v�������8l���追]��6�|�YR��vj��,8��l���Ҿ���R���ӿ��޿�   �   ���a�����������ܿ�u���Ú�oWs��T6�������[�:A�^G��x�h������ҽt�+�1������L�z-�S�V��q~��ې��������$۪�r���b���������X�O\.��
��eþTH��a-�|/սꩈ�fk�����b�N�[�Ԧ��;�b�5�8r�)HX��:ۿ�m�����v5��   �   uW4�!M1�U"(�@��@a�~����ү��Fg��&�	�������+���� xa�8�9�T�}�>�ҽى*�����ô��n��c��*4�M�N�{�c�=q��u�X�q��d�+�O�Aq5����Î񾝄��Wま±,��ֽ����$1>��Te���½͉,�Y����ᾜ�%���f��7���꿿'Q���s(��e'���0��   �   �W\�9X�7L���9�]�#����$��鷿�@��ՉK���������W��7��m� 2 �D
��~T�(���"��IZb��ƾ"���]��x��=$���'�9�$��$� <����A�Ǿ:��'Me� ������g[�~�����cr�l��.Y��Ŵ� �'�K�;��d���>P�f#���"���8��3K�K�W��   �   m���J��=�r��Z�Z�>���!����ZgտU����Uo�o�%�bJ׾"���8 �Nς�������@9Z�h���4���M����4���p� ꕾ\S��XVžH�Ҿ��׾�{Ӿ�Nƾ����1W��t�s���7��E��������8v�0!�T�Ƽ-��V��;̂�R~ؾHH&�Bp����Ԉտu��p�!��T>�i�Y��q��
���   �   ���Ql���V���{�l�X��o6�L���4ￂ!��c��$�<�^���`����#�~򑽘h��ئ
<05m<��;��
�J��.���:�s�*�K�N���k�N7~�aw��� �m���P���,����갶�BS�0ꢼ��-; 3Q<@�;PǢ��ꕽ�R%��������2�=������ʸ�l��+�:y6�c�X�Y�z���9���   �   O����}��鿜� f��g�n�#DG���"�����ȿ$�����N�c�������5����p���|��<4u=2�=lם<@�ʺ�q�Ztd�-%���޽>K�eh��%����p��1Ὗ����l�L��,_�0!�<�=�<m =�B�<t)������,�7��q��	�nP���ɿ�J��J#��G�v!o��^��S����a���   �   �������j̧��Д���}��xR��+��.�=-ҿx���AZ�8��'���@�m��}{�(b�<��2=hC=l|&=h�<��;({� u���d������ĥ�����Ҧ������Hj�&��D�����;���<�v=�o<=X�+=���<����ˮ�f�C�}��$C���[�煜��ӿz����+�vLS��l~�z���m֧����   �   �
���a��TҴ��-��P����0`��O5�����0޿����Oh���&F��M�Q������߫�`��<�+2=�ZJ=�?4=\m�<��Q<�����߼�8��r��݋��c��#B�� t�z�:�0b���� vG<�/�<l�1=b�G=�/=D��<�a������IS����S���h��6����޿�O�p�5���`��.��!L���޴�_d���   �   ʞ����8������s#��0�[�12�����ڿ2�c����;����tM�kԺ����th�<�#=~�4=8�=4̰< i�:X���0�i��T��|۴����F������t��V�2� ��� �I:hf�<p=~�1=n� =|��<�b��忼�k�N��M��ne���d�`d���%ۿ�����2��N\�(I��������������   �   �����e��@����r�� ,z���O�lA)���@пf͙���W�1u�����FA��s�����P�h<x{�<���<8�p<�߻�	������~���{���>�����~��M�K�뼽67��������(�e<;�<�#�<��]<�¸�*<���%B�-[��x��pX�[.���vпh
� �)��P�MGz��o�����Y���   �   9����/���^��:}��xb�J�=����j���m�����CE��d�L蝾�..�������ü��l;�� <���$�¼�Bg��4ýH7�y�5�4h[�y�C��%y���F��%�y�$2\��6��#�LŽ4�j�@ɼ@����<�0B;<%ɼF0��o /��}��X��9tE��L����������H����=�]b��`���<��g���   �   ���Ȇ���}�@d�%�F��5(��
���ݿ.��pcy�-���ᾎ���T�"�����(�R�����"7/�&<����X�@��2��#���|���/Ͼ.,ݾj�zeݾ7�Ͼ���뺞�n1����A��������>2�TD��8�\�x������������c�xZ-�
�y�]N���ݿ��
�U(��gF�J�c��W}��i���   �   M2f��a��T��A�z�)�����o��쾿[ߑ��2T����,���od�P���������p����p�x�νFz$�Cp�<���Gо�o�����d�!�P�+�/���+���!��L�=���Ѿ(����Rq��y%��}нXps��/��B�������e�y���6�uIT�+ݑ��Ѿ��-�Đ�r_)��@��'T��ha��   �   S�;�CJ8�~�.����DN������ǿ����[{p��Q-��W�~�����6�Êѽ��|��S��u��M��`�5�퇾lD��>��y�wX<��W�Rm�t&{����0`{��m��BX��<����(#������~����6��������j�U�bO~�);ҽI	7��Η��^�6A-�aHp��b���ǿ+l���PK�5.�+8��   �   ^���p�6� �>�俵\ÿ&�����|���=��k������#h��{����i끽�l��M�=7�c���d�˾�h���4��`�����	斿j/���R��Ä���{���x���@��V
����`�t�5�����n̾�#��Y�7�X+�l
���[��\��8��{h��h��B��=�1�|��C����¿���� ��,�����   �   �2뿫M�Z�ۿքɿ	0������bw��@�!'��]ɾǅ��r(��Cн�8��%#��1�Ͻ�+(�������Ⱦ���np@�I�v�.��ظ���ɿ�Zۿ��u6뿃Q� �ۿ.�ɿ3������Ngw���@��)��aɾ�Ʌ�lv(�QGн�9��L!��t�Ͻ�'(�w���"�Ⱦ����l@���v�J+������1
ɿ'Wۿ��   �   V����x��ou���=�����,�`���5�����i̾6 ��°7��%彥���[���^����6h�l���D�1�=�^�|�dF����¿j���� ��.�*��A`�>��#r�� ���俄_ÿ������|�|�=��m������'h�~�{��\ꁽi��_F�7�����g�˾�e���4�%�_�٩�� 㖿),���O���   �   ����Z{���m��=X���<�?�����%��� {��s�6�+��S~����U��P~�h>ҽz7�xї��b��C-��Kp��d����ǿMo����gM�Z7.��8�ݤ;��L8���.�����O����Y�ǿ����q~p�6T-�9[쾤���6�6��ѽ��|���S��p�� �q�5�釾2?���7��#u��S<���W��Lm�� {��   �   v/�J�+�|�!��H�=6���	Ѿ[���Kq��s%�~uнes�P)���l���M����e��{���8�LT��ޑ�Ծ�]0�[��[a)�&�@�*T�~ka�-5f�˥a���T��A�@�)�@��1r�������4T�k��.��Hrd�����B�����\���p�H�νt$�/p�/ ��lAо�h������!�ъ+��   �   ���^ݾ��Ͼ6���ᵞ�"-����A�>���񧽄22��3�� \����F��s�����3f�Q\-���y��O���ݿ�
��(��iF���c��Z}��j������>�����}�5Bd��F�U7(���
�t�ݿl/��yey��-�������V������鼠iR��͚�t)/��2�������@��)�p���v��J)Ͼ�%ݾ�   �   �t��mB����y�S*\�-�6�����Ľ��j�lɼ ��X <@^B;8%ɼ�1��)"/�W��x���uE��M������X���_��U�=��^b��a��&>���������'1��/`��<~���yb�z�=���l���n���	��qE��e�F靾�/.����T�ü`�l;�� <��8�¼h2g��*ý"1�U�5�3`[�[y�����   �   ���ky��H�lA�⼽�/����� >����e<�E�<p*�<�]<�ø��=��='B�X\��Z��?qX�-/���wп�؄)��P��Hz��p�����Z�������f��+����s��1-z�l�O�B)�����п�͙���W��u�H����A�t��Ы��H�h<l��<���<`q<��޻6�	����v��,���,9��   �   ����A�����Tp��^x2�(�����J:ho�<�=��1=�� =<��<ld������^�N��N���e�U�d��d��p&ۿ��%�2�9O\��I��<���������Z���������������#����[�M12�Փ�`�ڿhS�c����p����tM�LԺ�@����k�<8�#=��4=l�=|ְ<@4�:I���0�Sd���N��&ִ��   �   �c��2B��&t���:��b�Ё��tG<�.�<�1=��G=d�/=���<Hc�������S���AS� �h��6����޿�O���5�ߡ`��.��2L��ߴ�ed���
���a��HҴ��-��?����0`��O5�����0޿a���h�����E����Q� ����ݫ����<,2=@[J=�?4=n�<��Q<���p�߼��8���r�z݋��   �   ����A�����Vp��Nx2�,��� K:�o�< =f�1=�� =��<`��<���
�N��M��;e�E�d�)d���%ۿt��X�2�$N\��H��T���}���d��;���m����������#����[��02�>��v�ڿ��E�c�.��l����sM��Һ�����pn�<�#=>�4=��=�ְ<�7�:I��0�[d���N��.ִ��   �   ��uy��H�sA�⼽�/��|���:��H�e<�G�<�-�<`�]<����M:���$B�gZ�����9oX��-���uп�	�]�)��P�Fz�o����X�������d��?����q���*z�w�O��@)�w��7 п�̙���W�Jt�[���e	A��p��������h<���<��<�q<а޻�	�����
v��4�$��69��   �   �t��vB����y�X*\�+�6���h�Ľ"�j�� ɼ�٦��	<��B;�ɼT-���/��|��~��sE��K�����:���a����=��[b��_���;��������i.���]�� |��<vb���=����h���l�������D��c��松q,.������|ü� m;�� < ����¼�1g��*ý1�W�5�8`[�hy�����   �   ���^ݾ��Ͼ:���ᵞ�-����A���z��02�L.���m\������J�j����a��X-���y�M��T�ݿ��
��(�fF��c�MU}�
h������J���8�}��=d�:�F�n4(���
���ݿ|,���`y�/-� �ᾘ���Q�7���\��PXR�8Ț��'/�u2�������@��)�r���v��R)Ͼ�%ݾ�   �   }/�O�+���!��H�<6���	ѾP����Jq��s%��tнbs��$�`������M���e��v��5�+GT��ۑ��Ͼ�`+�R���])���@�%T��ea�n/f�8�a�v�T�TA���)�8��6m��꾿�ݑ��/T����)��|kd�ƍ��q�����������p�j�ν�s$�p�' ��jAо�h������!�֊+��   �   ����Z{���m��=X���<�;���������z����6�����{���U��D~�[5ҽ�7�i̗�i[��>-�HEp��`���ǿDi�[��RI��2.��8�̟;��G8�)�.����qL����H�ǿq����wp�8O-��S쾗���d�6���ѽ2�|��S�$n���}��5��臾!?���7��"u��S<���W��Lm�� {��   �   Y����x��pu���=�����*�`���5�����i̾ ���7�c#���.V��
V������
h�9e���?��=�\||�~A����¿���9� ��*�ѱ��[����n�N� ��|俷Yÿ������|�/�=�i�����h��w��
���䁽{e��#D�d7�����N�˾�e���4�&�_�ک��㖿,,���O���   �   �2뿯M�\�ۿքɿ	0������bw��@�'�x]ɾ�ƅ��q(�f@н�3��X����Ͻ4#(�s���	�Ⱦ���'i@�S�v��(�������ɿ�Sۿ<翠.��I翢�ۿ_�ɿ�,��D���Q^w�P�@�#$�Yɾ�Å��m(��;н�1��9��9�Ͻ�&(�-�����Ⱦ����l@���v�K+������4
ɿ+Wۿ��   �   
^���p�7� �>�俴\ÿ%�����|�y�=��k�d����"h�vz�����䁽�b��r>��7�,�����˾�b���4���_�<�������(��)L���}��:u��.r���:�����h�`���5�b���d̾S���7���Y ��%U���W��Ԉ��h�Mh��B�ߪ=�.�|��C����¿���� ��,�����   �   V�;�FJ8�}�.����DN������ǿ����T{p��Q-��W�)�����6��ѽb�|�^�S��i��=v你�5�A凾=:��[1��eq��O<��W�HGm�({�;���T{�5�m��8X�"�<�N��c�������v���6�f�形v����U�D~�7ҽ&7��Η��^�,A-�^Hp��b���ǿ+l���QK�5.�.8��   �   O2f��a��T��A�y�)�����o��쾿Zߑ��2T����,���nd�j�������p��6����p��νn$�zp�]����;оb������~!�`�+��/�ή+�1�!�E�%/���ѾA����Bq�Vm%�ckнDUs���������������e��x���6�oIT�*ݑ��Ѿ��-�Ő�s_)��@��'T��ha��   �   ���Ȇ���}�@d�$�F��5(��
���ݿ.��lcy�-����<���S��������hFR�����x/��)������@�j!�j��q��#Ͼ�ݾ��@Xݾ��Ͼa��������(��j�A���<觽#2�0�� V\���U�������xc�oZ-��y�_N���ݿ��
�V(��gF�L�c��W}��i���   �   :����/���^��:}��xb�J�=����j���m�����=E��d�蝾(..�����|ü�Nm;� <���ع¼t"g�� ý:+�s�5�lX[��y�6���o���=���y�T"\��6�t�$�Ľ��j���ȼ@����$< �B;`ɼ�-���/��}��K��3tE��L����������I����=�]b��`���<��g���   �   �����e��@����r�� ,z���O�mA)���?пe͙���W�(u������
A�*r��������h<d��<���<`4q<@c޻��	������m���������3�V���s�:C��7�ټ�0(�����@�����e<TT�<�6�<��]<@����:��V%B�[��q�� pX�\.���vпh
��)��P�OGz��o�����Y���   �   ˞�� ��8������s#��0�[�12�����ڿ1�c����*����tM��Ӻ�\���,o�<t�#=��4=�=�߰<��:x;���/��_��J���д�e	��L<������k���o2�0�����L:Lz�<\#=��1=� =T<8^��#���0�N��M��ke���d�_d���%ۿ�����2��N\�(I��������������   �   �v������2���r��L���a�R�6�n����߿? �� �i��%�J3��TqT��J½4����ժ<xG.=R�F=�k0=0F�< Z@<�$�؅�*�=�Xuw�I��p[���卽v�v���<����� �E<��<$�1=&H=B�/=D׭<$����H���S�ɾ�����i�x���*�߿���t6�a�a������c���,�������   �   E��$i���
��k͝��*��R�]�V}3���c+ܿ�,���e��5�-d��&P�����L��h��<�=n�0=��=.�< ٖ9|h���Z5�`��;���ER���A��������U����4����� �&:t
�<�+=�$2=�!=l{�<p������tO����"��%de�����ۿl��K3�'e]����/Ý�u��Gj���   �   �������"��>}��Y�{��IQ�nc*�T���vѿ���Y����h����C�����\w����V<�*�<d8�<x�^<����n��Ƀ��ʾ�{w�;��&��Da �����I����}��" ����������d<��<���<��\<�O�������B�(��z��CY������<ѿ|���B*��.Q�3�{���Q*�������   �   �,��%G���S��^M��Y�c�o�>�F�������������Q�F�q���{���l0�@餽�μ �";(�<@?��ͼ�m���ƽ\D��<8���]�.r{��<���}��p'��#{�-Y]�!�7�@��G�ŽR�k��ʼ�
��x?<�H9;�˼�����/��0��R��LF�X捿��������{���>���c�?\���e��#S���   �   Q����`��h!�ile���G�b)�r^���޿
5��B{��V.���Qn���N�츔�L��H�e�X��\5�������xHC�Q�������*��i�о��޾ӏ�+�޾k�о*亾Zj��Y���H�B���iǨ�`j3�D*���n`��M�8
��i��h6�����	3.��z��%��P�޿�c�<)���G���e��P��o���   �   �g��b���U���A�Td*��d�����߿�®��΃U������=�f��� ��m��������ؙv�(qҽ�&�p�r�`����EҾ���� ��"�ȹ,�T"0��,�/�"�����B���ѾZ��4Fr�21&�ϓѽ�)u�������↽�� �df�w�����DzU�#���￿��{����*�f	B��U���b��   �   ڵ<��09��B/�^@ �M������ȿ�O���q�WS.�������^�8�{aԽW���P�X��A�����[48��a��*!�����������=��gY�� o���|����D�|�K�n�$Y�}�=���F��D�������7�0F����D�W��{��J	Խr`8�AԘ�D��].�,�q�ek��f�ȿ[���@q ��m/�fJ9��   �   y,�������T��C��
ĿJ=��!~���>�e(�㳷���i�2���i���+���ꗽ�d��"9�h����;6����6���a�8�������O���e���{��eP���)���ӗ�ᄅ��za��96��e��S;׍���8����I���e���E��4���i��ɷ�.?�*	?�R~�6m��qKĿ~��B}���ћ��   �   q쿎[近�ܿa<ʿ�˲�d���Ox���A�e���gʾ}���,�)�GWҽ�#��s2���ҽ*�)�o���ɥʾ�����A���x�$W������~ʿ%�ܿ�|�u�k_�:�ܿ�?ʿ�β�����Sx�;�A����kʾ;�����)��Zҽ�$���0��K�ҽ�)�S���`�ʾ�����A��x�cT��l
��4{ʿf�ܿ	y��   �   �x��M���&���З�=���mva��56��b�UO;�Ӎ���8����y���C����G������i�vͷ��A�z?�KV~��o��tNĿ��/�� ����.������V�G��Ŀ�?���~���>��*�������i�s��5k���*���旽^罎9����}�;����6���a�w���u���GL�� b���   �   7�����|���n�Y��=�\����X������z�7��>罧���z�W�h|���Խ�c8��֘���N`.���q��m���ȿ��}��[s �p/��L9�k�<�L39��D/�aB ������\�ȿ�Q��&�q��U.���☾�8��cԽ�߀���X�\<��[��d.8�x]�����$�������=��bY�%�n�3�|��   �   �0���,��"����;��(�Ѿ3U���>r�g+&�f�ѽZu���ȸ��ㆽ˶ �qgf�#����
��|U�ಒ�.񿿰������*��B���U��c���g���b�~�U���A�f*�Cf�Z��῿D����U�b�-���֯f��� ��m��������v��gҽ��&�N�r�J����?Ҿƥ������"�@�,��   �   �㾉�޾$�оl޺�He�����.�B�r��վ���]3�����\`��K���G��8��H���4.���z��'��S�޿-e��)���G� �e�eS�bq��ۋ��Zb��$��ne��G��	)��_�R�޿d6��P{�X.��㾇o���O�h���X�󼠢e�󤼘�4�[����� AC����o����$���о��޾�   �   �x���"��g{�QQ]�0�7�T����Ž��k���ʼ���� V< v9;�˼����/�i2��,S�<NF�l獿���P����|�M�>���c�]]���f���T��m.���H��/U��dN����c���>�/������ү�������F�?���|���m0��餽�μ ;#;h�<@���ͼZ�m�l�ƽ,>��58�˹]�ni{�P8���   �   �[ �d���D�������������������d<�#�<��<`�\<�P�����S�B�R���z�
EY����=ѿ$��^C*�0Q���{����T+�������������#��~����{��JQ�d*�ϱ��wѿa򚿬�Y�����h��3�C�9���u���V<�3�< E�<�^<�|��a�������m�Ӂ�~���   �   x<��W�����ʌ���4�,��� 4(:��</=$'2=R!=@|�<�������uO���������de�L�i�ۿjl�!L3��e]�(���Ý�	���j������i��/���͝��*����]��}3�#���+ܿ�,��j�e�!6�ad��NP�����h �����<j�=��0=�=�8�< �9hY��RR5������L���   �   p[���卽��v�(�<��������E<��<��1=� H=��/=֭<Н��4I����S�[ɾ���X�i�����T�߿��0t6���a������c���,�������v������2���r��;����a�7�6�V����߿ ����i��%�3���pT�J½�����֪<�G.=��F=�k0=�F�<X[@<�#�D����=� uw�;���   �   �<��`�����͌���4���� ;(:��<d/=�'2="!=�~�<����Y����sO���������ce���|�ۿ�k�UK3��d]�n��������i������h��#
���̝�"*����]��|3�����*ܿ,��Y�e�_5�[c���P�̈́�����l��<H�=8�0=|�=9�< �9XY��NR5������L���   �   �[ �l���D�������������� ����d<�%�<�	�<�\<�H�������B�c��zy�CY�F����;ѿ���A*�.Q� �{�M~��c)��������������!��Y|����{��HQ��b*�����uѿ񚿦�Y����f���C������l����V<<7�<G�<��^<p{��a� ������m�܁�����   �   �x���"��r{�ZQ]�0�7�L��\�ŽF�k�X�ʼ�ɶ�H_< �9; ˼����/��/��1Q�oKF��卿���2����z���>�4�c�;[��Hd���Q���+���E���R��@L����c��>�.������\��������F�C�z��j0�8夽�ͼ�v#;��<���$�ͼ܈m�E�ƽ$>��58�ι]�yi{�W8���   �   �㾓�޾,�оt޺�Ke������B�P��Z���D\3�L��@K`��=�N�����4���~㾇1.���z��$����޿�b��)���G�n�e� N�gn��ƈ��^_����je�̡G��)�3]���޿n3���{��T.�V��Xl���K�����x�� �e�����4�ݩ�����@C����p����$���о��޾�   �   �0���,���"����;��&�Ѿ+U��o>r�'+&���ѽxu�j��R���݆�K� ��`f���� ��wU�����������ڎ*�?B�c�U�&�b�0�g�8�b�^�U�s�A�ib*�5c�V�ݿ�����U��������f�c� ��g����������v��fҽd�&�&�r�A����?Ҿť������"�G�,��   �   :�����|���n�Y��=�Z����H������
�7�a=�G�����W��v��xԽ�\8��ј����I[.��q�ji����ȿp����=o �xk/��G9�M�<�R.9�=@/�F> �x�����F�ȿxM����q��P.����ݘ��8��ZԽڀ�<�X��9������-8�V]������������=��bY�)�n�9�|��   �   �x��
M���&���З�>���jva��56�}b�;O;�Ӎ�8�8����掗��ꃽ?�����F�i��Ʒ��<�'?�>N~��j���HĿ;��i{�y����?*��������R�Q@��Ŀ�:���~�n�>��%����j�i�����b��
%��D㗽�[��9�}��a�;���6���a�x���v���IL��#b���   �   "q쿓[迕�ܿd<ʿ�˲�d���Ox���A�Y��hgʾ2���/�)�Tҽ����*��S{ҽ��)�I���>�ʾ���D�A���x��Q��k���wʿ��ܿ2u�/m쿬W�ؖܿ�8ʿ�Ȳ�����Jx��A�b��cʾ����)�GOҽ����+��ҽ�)����3�ʾ�����A��x�cT��l
��8{ʿj�ܿy��   �   |,������T��C��
ĿI=��~���>�T(�����$�i����3e���$��}���V�F9�%��ß;���{6�(�a�կ������I���^��u���I���#���͗�����qa��16�@_�:J;�ύ��8����'����都�@�����@�i��ɷ�?�"	?�R~�5m��rKĿ~��C}���қ��   �   ޵<��09��B/�_@ �N������ȿ�O���q�MS.����1���<�8��]Խ�ڀ���X��5����罉(8��Y�������������=��]Y���n���|�V����|�t�n�Y���=�j��z���������7�
5�򥏽h�W�)v���ԽJ_8��Ә���].�&�q�dk��d�ȿ\���@q ��m/�hJ9��   �   �g��b���U���A�Ud*��d�����߿�®��ȃU���ñ��[�f�7� �i��h��H���~v��^ҽ��&���r�o����9Ҿ�����\�"�˰,�10��,���"�!���4���ѾP��R6r��$&�N�ѽ�u�L�����ކ��� �/cf�7�����=zU�"���￿��{����*�h	B��U���b��   �   Q����`��i!�ile���G�b)�r^���޿
5��A{��V.�����m��pM�z������(e�ݤ�z�4�J������9C�}���a�������о<�޾N���޾˟о�غ�`��������B�S������N3����3`��8����P��6����� 3.��z��%��R�޿�c�=)���G���e��P��o���   �   -��$G���S��^M��Z�c�n�>�F�������������K�F�d��{{���k0��椽�ͼ �#; �<@��L�ͼ<ym���ƽ88��.8���]��`{��3��Qt��V���{�LI]�	�7�"���Ž��k�Xmʼ ���pz< �9;�˼���/��0���Q��LF�Y捿��������{���>���c�?\���e��$S���   �   �������"��>}��Y�{��IQ�nc*�T���vѿ���Y�����g���C�Y����m����V<�=�<�Q�<8_<�T�lU�����Z����c�|�����U �ȩ�@?�������񂽸��P<��p	e<,2�<��<�\<(F����p�B��� z��CY������<ѿ}���B*��.Q�4�{���Q*�������   �   F��$i���
��k͝��*��T�]�T}3���d+ܿ�,���e��5�d���P�х��������<��=��0=��=B�< ��9�K��XJ5���'�G��7���� ���
���4�0��� �):t�<�3=�*2=�!=L��<Ĭ��@����sO�������$de�����ۿl��K3�)e]����0Ý�w��Fj���   �   �g��'Լ���������ב��}N[�Z�1��p��iڿ�ԡ�־c�A���W����L�!����w��Ĳ�<�X5=�0M=�t7=�U=(�g<�~��LμJH.��-f�a˄�y���#���8,c�J6*�Ѐļ0�����}<�=��<=�R=��:=���<��'���TbJ�����ͷ��Tb�砿k:ٿǷ��1��}Z��:�����戯��ϼ��   �   ���*���:����9���Ł�7W�t�.�����ֿl���_�$��]�����H�]ܴ�Hl�����<'=|�7=�j=0�< :@;H}���/&���t��d�����@v��>&���͗�ܤp�D%!�����@c�;D��<�
 =*Y==�,=D��<�G��  ���+F��������I^��-��9�տ�p
��.��kV�������؎��=����   �   �q���(��[���U��2�s��BK���%��R�A̿L�����S����-ڪ��@<�@�������`}}<���<�#�<�<0���j���v��崽�)�$B���T�S��
S�-��Z�����p�R���t��o�<���<2� =�K�<p���覽�:��x����
�܈R��=��#e˿L��|u%���J���s�!\��F5���@���   �   P��'��������D�\�H�9��p��������C����@��D��pH����)�Ϭ��h���P#�;�	7<�2p:켳��]����GG�"-1��U�{wr�h���t��D���Fq�\T��a/�Si�;J��x�V��榼�-; �M< m�;���{��ͮ'�3%��k����$@�>ĉ��5���#A�#�9���\��	���M�������   �   `ʆ�����n�v�^�v�A�z\$�5���ؿ����4"t�M)���ܾ�����������L7ؼ�j4��d��|&�,w���K�D<��Hy�����=��SNʾ��׾L5ܾ�K׾!�ɾ^0���_��}�v�x�9��D ��㜽���<'���v�X�ͼ	���g��҄�K�۾��(�ӕs�o����ؿ����$�A4B���^��;w����   �   �{`��[��N��<���%�~j���ְ��K���a^O����{��%+^�� ���:}�����D���e��"Ƚ0& ���j�J}��1�˾�/�������M�'�<�*�'Z'��u��"������_ʾ���h� ���Ľ
L`��f�8�
���x�l���	]�S귾6d�T6O������溿4������,&�_�<���O��2\��   �   �j7��3��>*������	�\"쿮ÿњ��j�f
)�3E�B���]1�lɽ�p�\H�E:����ܽ�1�O�B3��^&��L_��8�j{S�F{h���u�3z�AZu�j�g�6}R���7��]��c��u���x���aU/�x7ڽ�����D���l�Ƚ�m0��P��X=��-)�Lk�G6��u�ÿ��~
�zl���*�D4��   �   /1����*	�m����޿��������v�69�6��Y����`��E�� ��v�gm���ܽ��1��?��OǾl���y1���[��8��$������˪����R}��
v���g��!�����Z��d0����ƾ�X����0�}Hڽo#���Et�����-�a�������3�9�~zw��H���n����߿R�����	�t���   �   H��#�A�ֿ��Ŀf��������p�ɡ;����\þ0m���!"�4�ƽ?���r��4Zǽ��"�E����8ľ�����<�Rr�>s�������{ſQ׿����K濿'�АֿD�ĿR���5���O�p�6�;�f��`þ�o��%"�ٶƽ�?���p���Uǽ޾"�=�@4ľ����<��r��p��꒮�dxſsM׿.���   �   ����z���r�� e������~Z�a0���		ƾ�U��@�0��Bڽ� ���Et�����>0��a�	���%�m�9��~w�?K���q��S�߿�����	����Z3�և�$ 	������޿z���f�����v�!9�`��\����`��G�)"��&v��i��`ܽu�1�!<��,JǾ@���u1���[�6��'������PȪ��   �   j-z��Tu�,�g�cxR�t�7�Z��]������ҙ��P/�D0ڽ���мD���l�>Ƚq0�#S��A�u0)��k�l8���ÿ�!��
��n���*�rF4�4m7�w�3�A*����3�	�6%�ÿ�Қ��j��)�iH�a����1�>nɽp��VH�5����ܽ�1�Z���".�����r[�p�8�pvS��uh�]�u��   �   ��*��U'�qq�������Yʾ_��Vh�y���Ľ�@`�H`��
���x����]��췾f��8O�a����躿Ǝ�g���.&���<��O��5\��~`���[�}�N��<�=�%��k��꿸���Ɵ���`O�@��<}���-^�'#��;}�����<��e��Ƚ  �
�j�Sx��6�˾�(���������'��   �   �.ܾLE׾{ɾ�*���Z���v���9�>? �Vۜ�������d�|�ͼ�
���i��Ԅ���۾��(�B�s��p����ؿH��-�$�6B���^�k>w�����ˆ�����v�,^�+�A��]$�F����ؿP���8$t�yN)���ܾ䮅���4���p2ؼ�S4�R��&�n��F��<�+@y�r���\7��Hʾ0�׾�   �   8p�����p>q��T��Z/��c��@��L�V�tϦ�@�;(�M<���;����|��w�'��&������J&@�Hŉ�7����.B�z�9�h�\��
���N������`Q��u���2����ν\�t�9��q�z�������D����@�zF��eI����)�O���D����C�;`$7< �r:p����t]�꼽:A�&1�(�U��nr��c���   �   �N����M�Ɵ�����}p�h:�� rs�l~�<��<�� =|N�<p��ꦽ":�z��z�
��R��>��%f˿���Kv%���J�W�s��\��=6���A���r���)��A���V��[�s��CK�D�%�7S��A̿������S�?���ڪ�dA<���������0�}<���<�/�<T��<Ū��]���v��ܴ����<�6��   �   �p��!��*ɗ��p�j!�������;��<� =~[==l�,=��<TI��%��r,F�d��:���J^�.��ӱտ1q
�4.�-lV�뀁����d���̌��|����������:���Ł��W���.���5�ֿ���V�_�U������ؐH�Jܴ��j�����<^	'=��7=*o=@:�<��@;�n��"'&�:�t��_��h����   �   |���1���`,c�|6*�<�ļ ���h�}<��=N�<=~�R=H�:=X��<��������bJ�켷����Ub�&砿�:ٿ޷��1��}Z��:��������ϼ��g��!Լ������Ǒ��_N[�A�1��p��iڿvԡ���c���NW����L�����v����<Y5=L1M=6u7=V=��g<�|���μH.��-f�R˄��   �   q��(!��2ɗ�
�p�f!�������;l��<8 = \==4�,=Ț�<E��}���$+F�h������I^�n-���տ�p
�r.�(kV�<������b�������b����������%9��BŁ��W���.�^�K�ֿ���K�_����������H��ڴ�<f�����<N
'=<�7=�o=�:�< �@;pn��'&�6�t��_��p����   �   �N����M�П�����}p��9��`ls���< ��<� =�S�<\���榽�:�*x���
��R�0=��od˿����t%���J�ڞs�e[��d4���?��|p���'��a��U����s��AK���%�R�@̿~�ĪS�ؐ��ت��><�Z}��x�����}<���<�1�<���<�����]���v��ܴ����<�>��   �   @p�����|>q��T��Z/��c��@��އV��ͦ���; �M<��;p���8x���'�$�������#@�qÉ��4����C@���9�0�\����_L��[����N��τ�����ۥ���\��9��o�j�󿁿���B����@��B���F��H�)�ب���y��a�;�-7< �r:����4t]��鼽-A�&1�*�U��nr��c���   �   �.ܾXE׾{ɾ�*���Z���v���9� ? ��ڜ�������T��ͼF���e�oф�6�۾S�(�ԓs��m��.�ؿ��\�$��2B�z�^�J9w�����Ȇ�@���͍v��^���A��Z$�����ؿh����t�/K)��ܾƫ�����޸���$ؼ8B4��L��H&��m���E��<�@y�q���^7��Hʾ7�׾�   �   ��*��U'�uq������YʾZ��5h�<���Ľ$>`��[��}
�P�x�1��w]��緾�b�4O�8����亿��r��+&�N�<�8�O�B0\�&y`�_�[���N��
<���%��h�
꿹��������[O����Gx���&^�M��x/}�Z��48��e�Ƚ� �܁j�Gx��/�˾�(���������'��   �   o-z��Tu�1�g�hxR�w�7�Z��]�����������O/��.ڽ6��n�D�P�l�hȽfj0�4N���9澑+)�?k�Y4���ÿ�}
��j�P�*��A4�Kh7���3��<*������	�N�ÿ�Κ�x�j��)�JA�h����0�Seɽx
p�(OH��2��<�ܽ`1�8���.�����o[�o�8�rvS��uh�a�u��   �   ����z���r��e������~Z�a0����ƾQU����0��@ڽ0���:t�&����)�T�`�W�����B�9��vw�pF���k����߿������	�X��/����$	��{��+�޿�|������ۅv�� 9����VU��,�`�nA����v�5f��ܽ��1��;��JǾ7���u1���[�6��(������SȪ��   �   H�$�D�ֿ �Ŀh��������p�ġ;����\þ�l��� "��ƽ:���j���Nǽ�"�G���:0ľ�����<�~r�n������uſ�I׿m��9D�5 ⿟�ֿ��ĿX��� �����p��;���DXþ�i���"�e�ƽK8���k��_Rǽ޽"���4ľ�����<��r��p��뒮�exſuM׿1���   �   11����,	�p����޿�������v�.9�'���X����`�:D�F���
v��c���ܽI�1��8���EǾE��r1�X�[�p3��D������Ū�Z����v���o��b���~��uyZ�"]0���ƾ�Q����0�":ڽ����8t�����,�0a�W�����)�9�xzw��H���n����߿T�����	�u���   �   �j7��3��>*������	�^"쿰ÿњ��j�\
)�E�򃓾B1��hɽ�p��KH�_.���ܽ1�����?)������W�%�8��qS��ph�ؽu��'z�,Ou�ڨg�usR�	�7�0V�^W������ʕ���I/��&ڽ�����D���l�vȽ�l0�IP��&=��-)�Dk�D6��t�ÿ��~
�{l���*�
D4��   �   �{`��[��N��<���%�j���װ��K���]^O�����z��I*^�����1}�T���1��e��Ƚ% �kzj��s��w�˾"���������'�S�*�gQ'�Bm� �	���Tʾk��Oh�(��Ľ�1`��S�z
���x�����]�귾$d�M6O������溿4������,&�`�<���O��2\��   �   bʆ�����n�v�^�x�A�{\$�6���ؿ����3"t��L)���ܾe������[���$#ؼ�04�h<��(�%�0e��^@��<��7y������1�� Bʾî׾(ܾ�>׾�tɾ%���U��_�v�B�9�J9 ��ќ�������<� �ͼ����f��҄��۾��(�Еs�o����ؿ����$�@4B���^��;w����   �   P��(��������D�\�I�9��p��������C����@��D��8H����)�c����y���v�;�C7< u:\����d]�H༽h;�X1���U��fr�$_���k��f�� 6q��T��S/��]��6���wV�����@b;��M<���;@󧼯x���'��$��M����$@�<ĉ��5���$A�%�9���\��	���M�������   �   �q���(��\���U��2�s��BK���%��R�A̿M�����S����ڪ�J@<��~������h�}<|��<\<�< ��<�u���Q�<�v��Դ����7��
�I�q���H�&��i�np�� ��`�r�菎<P��<t� = Y�<��9禽L:��x����
�ڈR��=��#e˿M��~u%���J���s�"\��F5���@���   �   ���*���9����9���Ł�8W�t�.�����ֿl���_�"��P���x�H��۴��g�� ��<�'=��7=�r=�C�<��@;a��V&�j�t��Z��U����k�����1ė�Ȓp�!�tr��;���<Z =*_==��,=���<8C��_���H+F��������I^��-��9�տ�p
��.��kV�����
��׎��=����   �   �w���-�����K���ǀv�B_M�1�'����Lο������U�+�h?��h�;��e�� �D�,��<�*F=��\=�(H= �=<F�< �k:�q����lk@���a�v�k�J�^�� ;�4k� 2~��cT;��<��=~�R=�Wg=h�P=��<@������l�7������\�q�S�a����̿����d&��2L�d�u�&����ܡ��'���   �   �b��|,��J���Ό��uq�o�I�-�$��f���ʿXޕ��	R�zR
�<�����7��ޞ���F��q�<&�8=�zH=h�,=p:�<@�<pA��#���N����ٖ�e����]��S���G��?��Pp��~=<T�<v
7=6�R=�C=T\�<�d��%����3�B/�������O������-ɿnl�K�#��H�6�p������>��k2���   �   �����Ȟ�dד�����Gc��>�Yp�����1���K$��G�F��i�5���Z�+�����0QP�,ϫ<��=��	=a�<�n�:X�¼d�P��͞�6=Ͻ6=�����Br
�,����ʽ����E��T�� $�;�.�<D�=z=$�<xB#�{����N(��>���� ���D�{
���y������غ��%>�yc��������"���   �   !\��
��O~��7�m��gN��y.������`��p
����4�>I�"̎��>�*܆�(0n�(C6<�\�<���;�;o���8�R�������!�m�C���^��#p���u��o�p]��HA��u�K��.����,��A��C <��<@�^<�D��A��s��쌾�	�͎3��D���3��r3� ��.o.���N�NWn�U؄��%���   �   Vz���t�3�e���O���5����� ���̿�뜿�;e��e��p;N�v�H���Ro�`���w����!�������m��+�ھe�����@�����T�Ⱦ�̾��Ǿĺ����3,����a��(�$y�oC��@��h��L�<����e��/���s�M�˾����`d�����Tx̿� ��+��}6�6|P��~f�dNu��   �   �Q��M���A���0�����K��ܿѯ���� KB���s��:�K��1ܽ�6V���ۼ�ּ�e@�$ ��fl�n�W�Rғ��ɽ�����}���u��!��uR�A���Y�� ��K������p�S�����.��x6��#ż�˼��N��qؽ��I��0��v��JB����2"��Giݿ���7���1���B�pN��   �   4|,��%)��( �[�����z�޿2����~��;\�����%־^��"� �ͯ���wI�H�#� �f���Ľ�[!�: u����t���s�^-��wF��KZ��f���j��!f�;Y�"�D�}r+����-��9���*7q�^��Ϳ���^���D��Q������ȇ�5־^(�k�\�\��5�����߿�������!���)��   �   b�
�+D��?�{ �0�ѿ�<�����g���,��V�����W�M���t%����N�*�s�!vý��!�VQ}�_T��[ ���N&�cmN���t��n��m���j㠿����k��Ɨ��b����r��iL��$�Po���L���Xz�d��Q]���3o�H�K��%��L�LN�����^����-�&�h�t(������r�ӿ��������   �   FBٿ 7տ�!ʿ,���@�����H�a�JH/� ~�H贾b�m��i��`����h�n�i�,{��Ru�}Ro��G�������0��c��΋�����f���G˿>�տ�Eٿ�:տ@%ʿH��gC������O�a��K/�����봾r�m��l�Ld��:�h�$�i��v���q��Lo��C��փ�N�0���c�#̋�%����c���D˿��տ�   �   ꋣ��h��&×��_���r��eL�q�$��i��cH��pRz�"���W���.o���K�K(��8Q�N�X���Gc����-��h��*��f�����ӿ������i�
�%F��A���2�ѿ0?��=��vg�k�,��Z��c���M�I���&����N�R�s��oý�!��J}��O��]���J&��hN���t��k��a���>࠿�   �   .�j�nf�EY���D�rn+�m��y�⾸���L0q�Y�$ǿ���^����D��T�����4ˇ��־�*���\�c������� �b������!�6�)�y~,��')��* �+��f��-�޿u���W���\�����(־] ��x� �ӱ���vI�B�#�B}f�݃ĽvV!���t����d��2p�%-�<sF��FZ���f��   �   ��UN�Y���U���nF������s�S�8��$'��~m6��żĢ˼��N�Muؽ��I�3��=���B�8��1$���kݿ(�����1���B��N���Q��M���A�|�0�V��M��ܿ�ү����=MB�D �s����K�'4ܽ$7V���ۼּ�Y@������f���W��͓�DĽ�&��z���I���   �   ի̾��ǾJ��������'����a�P(��n㽀;��4���*�@��`��z�e�~1���s���˾j��cd����,z̿� �G-��6�=~P�:�f��Pu��Xz��t�t�e���O�i�5����� �U�̿�윿�=e�3g�^r;��v�f���So����� K����!���h|���b�2�+���e����E;�����*�Ⱦ�   �   
�u�Ao���\�eAA��o�4@��%��D�,���@��c <8�<��^<��D�[C���)��D�3��E���4��5����fp.�=�N�1Yn�oل��&��[]��6��[����m�#iN��z.����\��e	��6����4��J�͎�x?��܆�8*n��R6<�i�<0��;0o�\�8���{���$y!���C���^�/p��   �   m
���Q�1�ʽ/���z�E�|>���k�;�<�<4�=�=��<0D#�����*P(��?���� ���D�:���z��,�������&>��c�U���j���������zɞ�3ؓ�D���Hc�޶>��p����������$���F�)j�΁����+������LP�Pԫ<�=��	=�p�<���:4�¼�P��Ş��3Ͻ:3������   �   g����X��ŵ���G��0���V���=<l\�<�7=j�R=�C=]�<(g��&��ة3��/������O�����.ɿ�l���#���H��p�e���?���2��c���,���J��3ό��vq�ΌI�r�$�g�.�ʿ�ޕ��	R��R
�l����7�iޞ�H�F��t�<V�8=�}H=\�,=0D�<�<P�@�|�РN��z��Ԗ��   �   t�k�^�^�� ;�fk��2~��_T;|��<H�=*�R=XWg=��P=���<h�����ʝ7�ˡ���\���S������̿ы��d&��2L���u�5����ܡ�(���w���-�����<�����v�'_M��'����Lοt�����U���$?���;�<e����D�t��<t+F=�\=)H=z�=�F�<��k:q�����0k@���a��   �   r����X��ȵ���G��0���V�(�=<�\�<�7=��R=�C=�_�< _�%����3�/��\����O�T���=-ɿ?l�
�#�ËH���p�����*>���1���a���+���I��hΌ�Buq�ًI���$��f�O�ʿ�ݕ��R��Q
�x���گ7��ܞ��F�tw�<D�8=r~H=��,=�D�<�<�@�n�ҠN��z��Ԗ��   �   
m
���]�;�ʽ2���p�E�(>��@n�;�=�<&�=0=� �<�4#������M(��=��C� ��D��	��y�� ���H��7%>�w c��������;��ɸ���Ǟ��֓�����Fc��>��o�����9����#�� �F��h������+�����=P��٫<��=��	=r�<@��:��¼ڙP�zŞ��3ϽC3������   �   �u�No���\�mAA��o�1@��%��ڄ,���@�i <d �<��^<`�D�2?�����댾\꾱�3��C���2��,2�0��"n.�Y�N��Un�Kׄ�c$���Z�����3}��N�m�0fN��x.����r����p	��W�4�G쾎ʎ�1<�]؆�n� a6<n�< ��;Xo���8�����[���y!���C���^�4p��   �   ޫ̾��ǾR���Ɔ���'����a�H(��n�;��<��@��E�����e��-�.�s�U�˾W���^d�Y����v̿� ��*�e|6�QzP��|f��Ku�dSz���t�ڇe���O�&�5�V��� �ڞ̿ꜿ�9e�d��m;��v�~���Io����� )���!�� ��{��,b��+�{�e����D;�����0�Ⱦ�   �   ��ZN�^���U���nF��~���U�S���[&���j6�ż�˼ΛN�mؽ��I�h.����-	B�:��l ��gݿa������1�e�B�
N���Q�D}M�H�A���0���SJ�v�ܿϯ�����HB������C�K��+ܽ,V�Puۼ�uּ�V@�����Pf���W��͓�8Ľ���z���L���   �   2�j�tf�JY���D�tn+�m��t�⾩���0q��X��ſ�&�^����$�C�rL��3���Ƈ�־/&���\����򯸿7�߿��٨��!�̬)��y,�f#)��& �y��&���޿����v|����[�!���!־���� �P����kI���#��xf�`�Ľ�U!�{�t����T��.p�!-�=sF��FZ���f��   �   싣��h��*×��_���r��eL�p�$��i��LH��Rz�����U���'o���K�S ��CE��N�����Z����-���h�@&������h�ӿ������[�
�-B��=�����ѿ�9�����g���,��Q��
��1�M�7�����0�N�^�s��mýU�!�J}��O��G���J&��hN���t��k��b���@࠿�   �   HBٿ7տ�!ʿ0���@�����G�a�GH/�~�"贾ޓm��h��]���h��ui�Xp��fm�)Go��?��K���0��~c��ɋ�Z���n`��A˿�տ�>ٿi3տrʿ�����=��������a��D/�^{�䴾!�m�
e�fY����h�vwi��s���p�,Lo��C��ȃ�E�0���c�!̋�$����c���D˿��տ�   �   c�
�-D��?�~ �2�ѿ�<�����g���,�jV��P����M����S!���N�T�s�{hý�!��C}�aK�����]G&��dN���t�0i��g���ݠ������e��"���]����r�)aL���$��c���C��EKz�����O��� o�~�K��!��UI�wN�ؖ���^����-��h�p(������p�ӿ��������   �   7|,��%)��( �]�����{�޿2����~��8\����g%־��� �_����lI���#�~pf��{ĽQ!���t������徵l�-��nF��AZ���f���j�*f�<Y���D�Gj+����r��֣���(q�'S�#���F�^�V��h�C�[N��|���ȇ�־P(�c�\�X��2�����߿�������!���)��   �   �Q��M���A���0�����K��ܿѯ����KB���8��e�K�/ܽP.V��qۼ�iּ^L@���`���W�!ɓ�Ѿ��Ǘ�|v�(��*�����0J�d��MR�$��@���|���S�F������^6���ļȍ˼
�N�4oؽ�I�^0��d��@B����/"��Eiݿ���6���1���B�rN��   �   Vz���t�6�e���O���5����� ���̿�뜿�;e��e�_p;��v�@��|Lo�������P�!�|���s���W꽌�+���e�.���5��1���Ⱦ��̾��Ǿy���c����"����a�r(��c㽗2�������@���	��T�e��.�]�s��˾����`d�����Sx̿� ��+��}6�7|P��~f�dNu��   �   "\����P~��:�m��gN��y.������a��q
����4�&I��ˎ��=��ن�(n�8k6<|x�< 7�;8�n�P�8��|��n����r!���C���^��p���u��o���\�:A��h��4�f��vu,���@�� < -�< 	_<�D��?�����쌾�	�Ŏ3��D���3��r3� ��/o.���N�NWn�U؄��%���   �   �����Ȟ�dד�����Gc��>�Yp�����2���L$��H�F��i������+����(?P�ܫ<��=��	=��<�٩:�¼V�P�����+Ͻ�)��j���g
���v���ʽ���N�E�L&�����;0M�<�=H=�%�<`0#�����mN(�c>���� ���D�z
���y������غ��%>�xc��������!���   �   �b��{,��J���Ό� vq�n�I�-�$��f���ʿYޕ��	R�xR
�.�����7��ݞ�ȫF�x�<z�8=��H=܈,=M�<�#<��@��n�N�Av��Hϖ�{����S������G� !��(;���=<�f�<�7=��R=�!C=�b�<�[��$��¨3�4/�������O������-ɿol�J�#��H�6�p������>��k2���   �   ]���ߙ�f���&���W]�p,:������������؊�"�A�²���&����"��
��@�Ⱥ��=Nc^=�fs=(0`=RV1=t=�<�o*<`�ڻț����	�V�'��r0��m#������� ea�f<N�=�B=�%q=�=�=�o=nJ#=�5A;&p������Pm��?�?'���o����4����8�#U\����mF���ٙ��   �   S���h���>����z��Y�W�6��_��t�VN���b���">����%敾��}�@�Ժ�0=��Q=�`=�F=�=��<���������LQL���m�.~w�fDi��?D����x�U;�!�<�`!=�W=�q=��b=��=��6;��i������������;�nˆ�ha���>��5�^�5�|>X���z�u3��o���   �   e��-���a����k�e�L�FY-���d�俬����;��U�3��$����nN��=k�`R�T;�<�*=�&=0G�<��/<`�J��+�C}�t��D�ͽ=g�D꽓ή8ɽ�ڤ���n�B���� u<$c	=��7=��;=�h=�;��X�B1�W�����澒v1�����w����T$���,�l�L���k������ʌ��   �   HN����|���l���U�8�:�����r��:ҿ�d��+l�*J#�W�Ӿ�5|�T��ZQ� x���<Lc�< `�<`p��\��腽��ν*�
�4'*�d�B�>TR�P/W��P��)@�~�&�bu��pŽ 7y��� =�9�I�<��<���< �8H�@�����<w��о�!��;j��k��9Uѿ�#�W���>;�DgV�:�m��;}��   �   ��`�q�[���N� �;�h`%��T�i
꿺˺��Ŏ�ɛO����-L��oYX�VM�L�4��/���>�; :l����Y��EĽ1Q�0JI�M�|�i��Gq���Ѳ��l��챾�ƥ�+.��T�w�s�C�<��S��R�G�(,�� ��;`�<Щ����&��"ٽ��T�DE�������N�#Z������I꿹���(&��<���O�#U\��   �   
�=�]$:���/�X� �30�D��}ɿX$��/7s�l/�a�ϗ�P1�����
w���u���l�$�	�QL������ �<�҂��5���ξq�������������� ���Y˾y������S7��>ۆ�����w8���E�PZ�bA��w.�V������n/��Ks������Xʿ��� 8��!�F 1�h�:��   �   �>�|7��"�<��.X��˿�T����`�F�G������po���	�_K���_��޼.|,����w
��'W�ڙ��;w���<�2|3���E��Q�$�T�|DP��.D�ߗ1��.������ ʾ�Ö�RR��L��<��D>!��?˼�a	��틽dQ��n��뾾!G��G�AԄ�'�����̿�|����#����   �   �������e5�Tqؿ�x���,��5�����P�͢�uV۾�!���v2�ygʽ��\�R����7������
�ۘ^������������:��P^�k�}��⊿�z��㔿�푿{剿{{�ï[�/c8�!����zb���Z�����V���x1�l%�,�Y���ɽ��2�Ǒ�{�ܾ����R�(ˆ�Qդ��l��?qڿ>�����   �   >wƿ��¿�_��ل��:j���I{���K������%V��=O������n����,�N�-�����`����Q�p���>���}8N�7>~����$�����,jÿ�zƿܬ¿�b�������l���M{���K���A��Y���AO�����r����,�H�-����������Q�����9�ʅ��4N�}9~�[���!��ӯ���fÿ�   �   ���둿�≿s {�H�[�T_8����փᾘ^��I�Z�����Q���s1�%�n�Y�;�ɽ��2�ʑ���ܾ�����R�W͆��פ��o���tڿ���F��_���H���8�stؿ�{��]/��;���Q�V��5Z۾l$��z2�SkʽL�\������7�.�����
���^�u��"�來����:�L^�/}�����w���   �   8�T��?P�]*D���1��*������ʾ޿��R�<H�v6���6!�(9˼�b	�h���T�E�n��[I��G� ք�m�����̿�￯�f%����@�o9��$����[�f ˿�V������F�@����8to���	�=M��_�T޼$s,����tr
�� W��ՙ���;���8��w3��E��Q��   �   �����������T˾�򥾙}���6�5�kԆ�h����`8��E�0\�iD���y.��������/�xNs�c����Zʿ����9���!�@1���:�4�=�r&:���/�� ��1����ɿ�%���9s��m/�&��kї��1�ҏ��fw�Шu��l��	�tD��D���#�<��͂��0���ξ���:�����   �   #g��u汾h���\)��տw�4�C�@	�TJ����G����@;(�< ����&�&ٽE�T�eG��,��̔N��[��W���K����*&���<���O�PW\�Ȋ`���[���N���;��a%��U�A�9ͺ�ǎ���O�י��M��[X�hO��4����g�;�$:�ꤼ��Y�];Ľ�J��BI�v�|�d���k���˲��   �   �'W�b�P��"@��&��o��fŽ�&y���� Y�9�X�<��<���< D�8ܢ@����G?w���о<�!��=j��l���Vѿ�$�j��@;��hV��m��=}�RO����|�]�l��U�m�:����|s��;ҿ�e���l�/K#���Ӿn7|�1��:Q� x���<o�<�p�<����M��߅�y�ν�
�e *��B��LR��   �   ��.���/ɽ�Ҥ�tn������/u<�i	="�7=n�;=*j= �;��X�j2�M���t�澙w1���}x�����$���,�t�L�@�k�a���\ˌ�4�����a����k�K�L��Y-����6��P���<<���3�t%꾍����N�2>k�`B�$@�<�+=X�&=�U�< �/<��J����3}������ͽ�]��   �   
uw��;i�@7D�������� �;�+�<xd!=��W=�q=2�b=�=`�6;n�i�`��#�������L�;��ˆ��a���?�_6���5�?X�O�z��3���o�����8i��	?��d�z�'Y���6�(`��t�N��c��#>�b���Q敾*���}���Ժ.2=
�Q=��`=��F=d�= ��<�&���	�����~HL��~m��   �   �r0��m#�,�� ᜼�ga�`f<
�=RB=t%q=�=�=��o=�I#= *A; p�n������m��D?�^'���o���I����8�<U\�̭�vF���ٙ�\���ߙ�vf���&���W]�W,:�k��n���򂼿�؊��A�p����&��]�"�%
����Ⱥ$�=�c^=(gs=�0`=�V1=(>�<�p*<0~ڻ\���n�	�2�'��   �   uw��;i�H7D���������;�+�<�d!=H�W=��q=��b=H�=`�6;��i�C��K���n���h�;�@ˆ�(a���>��5��5�>X��z�3���n�����Xh��?>���z�Y���6��_��s��M��rb��3">����q啾���}� XԺx3=��Q=F�`=��F=��=���<@$���	������HL��~m��   �   ��7���/ɽ�Ҥ�tn�����~�80u<j	= �7=��;=`l=�5;z�X�J0��������u1����w��� ��#��,���L���k������Ɍ����^���_`��6�k�U�L�jX-�l��E������;��C�3�#�ㅌ��L�z8k�@�E�<�+=n�&=W�<��/<��J�z��3}������ͽ�]��   �   �'W�k�P��"@��&��o��fŽd&y���� ��9�Z�<��<��< $�8,�@�����:w���о�!��:j��j��Tѿ�"�j���=;��eV�z�m��9}�@M����|���l���U���:�����q�K9ҿ�c��Ql��H#�S�Ӿ�2|�(��F Q� �w���<�s�<�s�<���M��߅�N�ν�
�^ *��B��LR��   �   )g��|汾m���a)��ٿw�5�C�4	� J���G����ԍ;��<�s����&��ٽ�T�vC��[����N��X��0���>G꿝��='&�v�<���O�S\�Y�`�F�[���N�]�;��^%��S�P� ʺ�~Ď���O�����I��VX�*Hཞ�4�����p��;��:`礼��Y��:Ľ�J�|BI�h�|�
d���k��̲��   �   ����������� T˾�򥾍}���6��4ӆ�t����P8�H�E�8R��<��!t.�M�����|/��Hs�造��Vʿ����6�q�!�]�0�S�:���=�A":���/��� ��.����L{ɿz"��24s��i/����͗���0�����m���u�`�l�:�	��C�������<��͂��0��ىξ���9�����   �   ;�T��?P�a*D���1��*������ʾҿ���R��G�85��|2!�,˼�X	��苽DN���n��达 E�k�G��҄����]�̿�y�P��!�*���<��5�� ����!U�>˿SR��:��c�F���v����ko�ڥ	�WE���T��޼�n,�"���q
�� W�yՙ�q�;���8��w3��E��Q��   �   ���둿�≿w {�L�[�V_8����̓ᾂ^����Z����O���m1�f���Y�5�ɽ{�2�Hđ���ܾ)��ºR�Ɇ��Ҥ��i��nڿ����������
���1�nؿ�u��e*�����'�P����)R۾����q2�)`ʽ@�\�����7�
�����
�-�^�P����|����:�L^�.}�����w���   �   @wƿ��¿�_��܄��<j���I{���K������V���<O����l��(�,�ֶ-�����Ψ����Q�>���4�ɂ��0N�5~�����������cÿ�sƿE�¿�\��恨��g���D{��K�ݴ����NR��F7O�#����g���,�,�-�	�������!�Q����l9����z4N�x9~�Z���!��ԯ���fÿ�   �   �������g5�Xqؿ�x���,��5�����P�Ȣ�[V۾�!���u2�eʽԳ\������7�D����
���^�r������H����:��G^�z}�B݊��t��ݔ�*葿�߉�H�z���[�K[8����[~�NZ����Z����J��(g1�~�:�Y���ɽ��2��Ƒ�R�ܾ����R�$ˆ�Nդ��l��>qڿ>�����   �   �>�~7��"�>��1X��˿�T����^�F�=������oo���	�*H���U�h�ݼ8g,�����km
�EW�Vљ�4�;���>5��s3�x�E�	Q�M�T��:P��%D�j�1��&�����.ʾk����Q��B�!.��P)!�|"˼�W	�gꋽTP�J�n��뾾G��G�>Ԅ�$�����̿�|����#����   �   �=�`$:���/�Y� �50�G��}ɿZ$��/7s��k/�I��]ϗ��1�'���o���u�x�l���	�i<������||<��ɂ��+���ξ�ﾢ���9��'�������)N˾o�u� �6�)*��ˆ�|����48���E�TR��>��Av.�������c/��Ks������Xʿ���8��!�E 1�h�:��   �   ��`�u�[���N�#�;�j`%��T�j
꿽˺��Ŏ�țO����L���XX�gK�<�4��������; �:4Ҥ���Y�p1Ľ�D�6;I���|�5_���f��oƲ�wa���౾���w$���w���C���@��BqG�������;��<�a����&�� ٽ�T�E�������N�!Z������I꿸���(&��<���O�&U\��   �   IN����|���l���U�7�:�����r��:ҿ�d��+l�&J#�?�ӾZ5|����Q���w�`��<}�<p��<�z��?�pׅ�J{ν*�
��*���B��DR��W���P�S@�-&��i��\Ž�y�x�� >�9�k�<|�<4��< �8�@�L��h<w��оݣ!��;j��k��8Uѿ�#�V���>;�DgV�9�m��;}��   �   d��.���a����k�f�L�GY-���d�俭����;��T�3��$�ㆌ�N��:k���dG�<V+=��&=�c�<P�/<�J��B%}���;�ͽST��齸���&ɽ[ʤ�en�����R�xTu<0q	=p�7=��;=�n=�F;��X��0�5����澍v1�����w����T$���,�k�L���k������ʌ��   �   S���h���>����z��Y�X�6��_��t�VN���b���">����敾����}� nԺ�3= �Q=J�`=ޝF=��=8��<�i�����0��&@L��um��kw�~2i��.D�ظ�@҉��;�6�< i!=�W=\�q=�b=��= �6;V�i�a��u���������;�mˆ�ga���>��5�_�5�|>X���z�v3��o���   �   ���� ����u�qF]�YA�l�#��o�8�ؿ�u����s�l�(���ھ`́�2j��~5��?5<��5=0`z=���=B�{=^�Q=��=h��<���;��޻��������μXj��@�m���C�`h:<@��<�1=�l=o�=6;�=O͊=�P=l�<B��3���nB{�z�վ��%�mLp�pc��vMֿ�7���"�"6@���\��[u�����   �   �F��v]����p�l�X�J�=�� !��+�Z�Կ����1eo���%�^c־S�}�
��/� <4<��/= o=nD|=��d=�t4=t]�<�	:< ���� ���
�Z��0�&�X�����O����&��3�<0k=��N=��=���=�=��J=��<�=�?��x�u���Ѿ��"�+l������ҿ�a( ���<�u�X��xp�"c���   �   �v��2q�Xjb�'�L���3��
��@���mʿ�1��ڐb�
D��vɾ�m�����h�-<y=r`L=�ZH=$�=�\�< ~�:,���P�.���}��Y���H��F����)���c��
�l��L�� z��c�;$��<(%9=��b=��f=)7=x��<�^�	p�:�e�U[ž�����_�����F�ȿw���D}��X3�0�L���b��mq��   �   � _�jZ�ßM�"�:�2�$�I��x�迂蹿���ƄN���ym���oS�4�ѽT*���<X��<�=8��<<e��y<�iݞ���ݽ��
�j �*�-��
2�~7,�M�4�B�ҽq}��Pb"��� �[{<P=ș(=�d=��s<ă� �Ž�UM�� ��]����L����$���Z����p�$��m;��CN���Z��   �   �C��?��5�-P%�I+��e���4Ͽ�ؤ��z�>5�ԇ��<D��D~3����<ۼ@�;t2�<��U<�������Mԕ�Mｦ�&��:T��|�yH���@��OR���3���O���kw���M�:��/:�B6��d�뼀�:��<���<��1<�������Z�.��噾�,����3��y���pϿ"6��n��^>&�	�5�1K@��   �   �('��#��5��!�����ķ׿����⌿��T��W�^A;�H���k�6���L�� "� �X�����ڋL�ÝýE>��\��
��j���rξDt�2��n��w��	�d.˾Z���&���T��#�C����"5��:I�@�;��i;TA���{��96�ϸ}�]̾����T�4A���ز�f ٿ6���4<�3��~$��   �   �*�@��wl��?�ҿ:o���L��&wg�(--�:���Ң��}G���ڽ�oJ��u�� �9��E˼�xk�wݽ%�2��h���c���n����&��F,��e6���9�y�5��*�f��;���۾�(��NT}��D,��ҽ��X�t���`J�8���dA��׽xmF���������l�-���h�#|������,Կoq��\�	��   �   ���ܿ_ѿe�����������i��6����_»�//t�I0��D��R��4蟼��ݼd?h�>ݽ9�A6����ľ�����"��VB�\1^���s����fՂ��%��A�q�S�[��?�� ��7��`�������"4��|սD\���˼����5������d�u�0>��c��n�7�̊l�.8��	窿�Y���ҿЖݿ�   �   2[��諿𠢿}Z���I���[��b1�
e��ƾ�d���^*�����peA�LgƼ�)ɼ6�E�r�Ľ D-����vɾcd
���3���^�K������#�~���6^���꫿����]���K��	�[�.f1��g��ƾ�g��c*����2kA�@jƼ�$ɼ6�E�a�Ľd?-��{��5rɾ�a
��3�g�^�����T���A����   �   �҂�#��[�q�ԑ[��?�Q ��1���������4��uսF;\��˼ ����g���x����u��A�������7���l�~:���骿�\��,�ҿ�ݿ\���ܿk"ѿ�g������(���D�i��6�ݠ��Ż��3t�R3�rH�����\埼p�ݼH5h�S6ݽ�9��2����ľ���S�"�`RB��,^���s�u����   �   "�9�-�5��*����8��۾.$�� M}�?,��ҽ��X�����0>��9���iA�~#׽HqF�X��������-�2�h�-~�����k/Կ}t￠^��	��,���n��B�Cҿwq���N��3zg��/-��=��>բ�>�G�]�ڽ�rJ��t���~9�p5˼&lk��ݽ�2�e���^���h�p�1"��B,�va6��   �   �g������⾚(˾�T��a"���xT��������5��I�`,�; �i;pD���~���8���}�=̾����T��B���ڲ��"ٿ�����=��4�{�$��*'���#� 7�#�,����׿���0䌿��T�qY��C;9J���m�����L���T!� �R�ح���}L�U�ý.8��\�f�����lξ�m�f���   �   BM���.��K��Bcw�m�M�̳��/��-��,v� :X�<��<��1< ��>�����.��百Z/����3���y�t����rϿR8������?&���5��L@���C���?��5��Q%�z,��g��:6Ͽ7ڤ��z��5�����E���3�����ۼP�;�;�<��U<PP�����?˕���&�3T�6�|��C���;���   �   �2��0,���X
��ҽ�t��zS"�} ��{<�=.�(=g=P�s<4�༉�Ž�WM�s"�������L����n	��6\�����$��n;�EN���Z��"_��kZ�1�M�Z�:�8�$�����进鹿����N�ڰ��n��>qS���ѽ(+���<���<Z�=P��<;<�K��Ni<�	Ԟ�ݩݽ��
��c �N�-��   �   ����i!���[��~�l��?���y�0��;���<�*9=�b=��f=P*7=䈉<�`�r���e��\žo����_�L���=�ȿ�����}��Y3�4�L�*�b��nq�S�v�4q�okb��L�`�3�4��A���nʿw2����b��D��wɾ�m������ȑ-<*{=�cL=�_H=��=$m�<@��:������.�fy}��Q��!@���   �   �&�d�|��(B�� %�H>�<�o=��N=X�=���=��=�J=���<N?�����u�o�Ѿt�"��l�����j�ҿo��( ��<��X��yp�}c���F���]��+�p���X���=�� !�,���Կ퓣��eo���%��c־��}�(��/��>4<(�/=�o=�F|=>�d=y4=Xg�<@!:<ñ�0���4���   �   ��μpj����m���C��g:<���<�1=�l=�n�=;�=#͊=n�P=�<*�������B{���վ��%��Lp��c���Mֿ�7���"�66@���\��[u�������� ��r�u�^F]�DA�X�#�yo��ؿ�u����s�=�(�O�ھ)́��i��}5�xB5<,�5=�`z=���=��{=��Q=8�=���<��;��޻0�|����   �   �&�j�x��B���%�P>�<�o=�N=��=Ъ�=��=�J=d��<�<�����u�R�Ѿ��"��l�ܦ����ҿ��( �A�<��X�Ixp��b��&F��]���p���X�Ɣ=�& !�r+���Կ3���jdo�&�%��b־�}� �(�/� F4<V�/=�o=�G|=��d=Jy4=�g�<�!:<0±����,���   �   ����l!���[����l��?���y���;���<T+9=��b=�f=^,7=H��<�[�Pn��e�Zž�����_�������ȿ�����|�X3�M�L��b�vlq���v��1q�'ib��L���3��	��?���lʿ1����b�C��uɾ�m�������ȟ-<t}=�eL=�`H=b�=<n�<�ɱ:쀫���.�Fy}�}Q��@���   �   �2��0,���\
��ҽ{t��RS"��{ �(�{<&=��(=�i=8�s<dz�C�Ž�SM����u����L������XY�)��r�$�ol;�.BN�d�Z�F_�khZ�?�M���:��$�S�����/繿����N�����k��&mS�H�ѽ�#��<0��<��=<��<0?<J���h<��Ӟ���ݽs�
��c �L�-��   �   FM���.��
K��Hcw�q�M�ʳ�z/ὕ-���t� l:��<ث�<@�1<`��󇤽�.�S䙾\*��&�3�
�y�����%oϿ/4��C���<&�t�5�vI@��C�#�?�B5��N%��)�Oc���2ϿQפ���z�P5�����(B��9{3� ��dۼ�K�;4C�< �U<pB������ʕ���Ȅ&��2T�)�|��C���;���   �   �g��Ē��⾞(˾�T��`"���xT���,���f5��I�PJ�; j;d2���w���3�+�}��̾� ���T��?��ײ�;ٿ�����:�m1��|$��&'�;�#��3�! �����c�׿����ጿ��T��U�T>;^F��|h�����9�� �� �N�8����{L���ý�7��\�T�����lξ�m�e���   �   $�9�0�5���*����8��۾)$���L}��>,��ҽH�X����p&�4'���[A�׽�iF�꺢�����-���h�Dz��U��*Կ�n�`[�Y	�)�����j��<��ҿ�l���J���sg�z*-��5���Ϣ��yG�Ňڽ�dJ�ta��e9��,˼Jik��ݽİ2��d���^���h�j�-"��B,�va6��   �   �҂�#��^�q�֑[��?�Q ��1���������54��tս�7\���˼`	��v�����F��W�u��:����}�7�(�l��5���䪿�V����ҿ��ݿ��࿤�ܿCѿ5b��s󨿱�����i��6�������|)t�,�a>��"���ҟ�8�ݼ61h��4ݽ(9�^2����ľ���K�"�ZRB��,^���s�v����   �   3[��諿�����Z���I���[��b1�e� �ƾjd��h^*����R`A�,WƼ�ɼ2�E�o�Ľ�:-��x��nɾ�^
���3�d�^���������o죿����/X��嫿����W��AG���[�[_1�-b��~ƾa���Y*������XA�<QƼ�ɼ��E���Ľ�>-��{��rɾ|a
��3�`�^�����R���B�����   �   ���ܿbѿe�����������i��6����G»��.t��/��B��D���ҟ�$�ݼ�(h�$.ݽ09��.��5�ľ��س"�SNB�!(^���s�ݯ��Ђ�w ��`�q�2�[��?�� ��+�����F���4��lսX-\���˼�����ų��/��߽u�>��S��b�7�l�*8��窿�Y���ҿҖݿ�   �   �*�B��zl��?�ҿ<o���L��'wg�$--��9���Ң�r}G���ڽ�iJ��c��8Z9��˼N^k�v�ܽ2�2�Da��0Z���b�|�o�{>,�(]6���9�܂5�Ҭ*���55�+�۾K��E}��8,��ҽ��X��������%���^A��׽�lF�P������`�-���h� |������,Կpq��\�	��   �   �('��#��5��!�����ŷ׿����⌿��T��W�EA;bH��k�߉���=�� `� �I�,���PoL��ý=2��	\�������gξcg徭���`����C�⾯"˾�O�����FqT���œ��`5���H��|�; 7j;�2��wy��l5�L�}�5̾����T�0A���ز�c ٿ4���3<�3��~$��   �   �C��?��5�.P%�J+��e���4Ͽ�ؤ��z�;5�Ƈ��D���}3��� ۼ�O�;�I�<��U<�������M��P~&�^+T���|�?���6��9H���)��NF���Zw���M���P$Ὄ$���X뼀	:�.�<P��<x�1<t��������.��噾�,����3��y�쩤��pϿ!6��n��^>&�	�5�1K@��   �   � _�jZ�ğM�!�:�2�$�J��z�迃蹿���ńN���bm��boS��ѽX&���<T��<��=T��<�c<X2���Y<��ʞ�K�ݽ��
�] ���-���1��),�l�[�,{ҽ9k���C"��H �8�{<�=\�(=Bm=��s<�{༰�Ž UM�� ��T���L����"���Z����n�$��m;��CN���Z��   �   
�v��2q�Yjb�(�L���3��
��@���mʿ�1��ڐb�D��vɾbm����
����-<�~=
hL=�dH=
�= }�<��:�j����.��j}��I���7��+�������S����l�82�H�y����;���<�19=��b=x�f=�.7=4��<\�<o���e�B[ž�����_�����D�ȿw���D}��X3�/�L� �b��mq��   �   �F��v]����p�l�X�K�=�� !��+�Z�Կ����2eo���%�Yc־:�}���Ɛ/��C4<��/=�o=RI|=@�d=�|4=�p�<�6:<𑱻d䥼`��F����&�V���3���v#��I�<�t=4�N=��=��=��=~�J=Л�<t<����Z�u���Ѿ��"�*l������ҿ�a( ���<�u�X��xp�"c���   �   "�^�Z�ZM�٦:�]$��w���述����ɍ�hN��J�Ї��kP�¸ƽ4�¼��<��X=YO�=iu�=���=��q=l�@=0}
=4�< p< �L:pc��`q��@!��d�;�v<��<<�,=�Gg=���=�ʠ=���=lN�=��=�"=��e�'��&oF��'��O
�X�J��狿����d����ح#��@:��3M���Y��   �   �>Z��U���I�|N7�|�!�Z
�����g���E���8J��
�A���i{K�����D,�����<�T=�v�=m�=���=�X=�.!=�6�<��)<`J��yB�ا�����8�������hZ;�َ<W=ОG=H��=���=��=�&�=l:~=U=�T�X���V�A�#���u���
G�Ʉ�����X�� V	�L� ��	7��xI�h�U��   �   	"N�{J�ا>�;�-�Mn�<R��gٿ\0������l?��n�s���
	=�\寽`5�����<�D=m=�Xi=�D=�	=@:�<�0\�h̳�,��<�P�r
p��x���g�F�@�����s� �;\9�<PB2=��n=&щ=�W�=(�l=L5=@A"�t4��i54�H��������p<�Ώ��Z̫�b+ؿ���<�Z�-�4�>��4J��   �   k<�r8�|d.��]�����ǿ�Þ��q�ֶ-����J����&��>��؀^����<̰(=*�8=��=|X�< !�9��μmV�� ��`yн�V��6
�Z6	����c����Ľ���d4�������$<�[=�nC=��_=
�M=,� =�緻�̆�T������美�+��8o�����?Mǿ���>�P����.���8��   �   g}&� O#���j��f	���ֿC`��^����S���8�˾T5}���8n�����<D�<$��<0!#<�f��z�G����� ��'�mSJ��We�,v� ${���s�H�`�q�C������～����Q!�p:ֻ|$�<�R=��=y�<������T��I��w�7{ɾ��A S��3��Ô��}�׿c8���g��c� �#��   �   1�E|�51��)��{Gؿ�и��ۗ�K�n��3������p����L��SٽtT,�@K��t<@Pw< p���輡㊽���5�.�a�h������ѩ�Gs��Ľɾ�};�WȾ�ͺ�N2�� s����_��8%�Ic۽�Qr��������;�w�<���<��;�^��DѽݟI�P4���!���3���o�W���	����ٿ������8���   �   ��P��lQ޿��˿F곿���Lz�i)C�����ʾ	郾���%����ۼ Bʹ ��;�Ļ�8��-���
�<~Q�s-��AY��L� \��4����T��R	���
= ��sܾ�S���L���kH�:��.������ �	��n,<`O`;�ü�Ǘ�e`�oԃ��1˾Q��k�D��?|�(�������-vͿ?�߿�p��   �   x���c(��,��5���`xs��=E��]��	߾�����A��/ٽ>;F��zd� �I������҃����x	b�ݩ���׾N�gJ#�LZ;��N���Y��]�,�X��)L���8�!� �xK�q�Ҿ�>��c�Z�f�	�{H��s�5��@-�:�O���D��ڽ�|C�yƚ����j;�T�G��v�����L���z�����   �   ����a����l���{��a\�u�8�"D�>��u)���X����y�����ż�����u����Ѽ&z��@v�e]��q���%澱����;���_���~�-���56��d�������fo����{��e\���8��F�����,��X�(�������żp��Pd���Ѽ�t��Kr���\��m��!澣��;�;�Z�_�C�~������3���   �   l{]���X��%L���8��| ��H���Ҿ�:��u�Z�
�	�lB���c�����:�:��O��D�	�ڽ �C��ɚ���(>���G��v������N��j}������T���1+������������{s��@E�z`��߾� ����A��4ٽNAF���d� lI�����F��,}��8	�b������׾-
��F#�>V;��N�O�Y��   �   �����r���9 � nܾ�N���H���eH�c��~��0�� �hy,<�F`;�ü�˗��c��փ�^5˾���O�D� C|�A�������xͿ�߿�s뿭�:��.T޿�˿�쳿����z�,C�����ʾ*냾ͣ��(����ۼ ʹ ��;�^Ļ�-�0&����
��wQ�=)��,T��#FᾯX�/1�����   �   �w;�QȾfȺ�T-���n���_�j2%�vY۽nBr�@���@0�;���<���<`�;6c�Iѽ3�I��6��?%���3�ݝo������$�ٿH���� �����2��}��2�x,���IؿsҸ�'ݗ���n��3�����s��j�L��Vٽ�W,��K�p't<pew< ����缄ۊ�����.���h�	����̩��m���ɾ�   �   v{���s�E�`��C�\��r��d�B!�@�ջP5�<XX=8�=�z�<�Җ���T�L�J�w��}ɾ���^"S��4��_���b�׿�:��i�*e���#��~&�gP#�;�����l����ֿ�a��8_��n�S�l��'�˾�7}�.�N;n� ����<�<���<�E#<�N���yG�;���Ҟ �L�'��KJ�[Oe�o#v��   �   b0	����T�콢wĽ����4�����h�$<�c=�tC=l�_=�M=X� =�����Ά��U����������+�a:o�	����NǿB��t?�_����.���8��<�Qs8��e.��^���.����ǿ�Ğ�]q��-�2��K��F�&�@����^����<~�(=�9=�=�i�< ��9��μ�\V�s����nнdK��O��   �    x�L�g���@�����r�0^�;�I�<�H2= �n=�҉=Y�=@�l=5=(H"�66���64�`���K����q<�|���2ͫ�d,ؿ|���<�(�-��>��5J�#N�kJ���>���-��n��R��hٿ1��c���)?�Ro�$����	=�:毽P6��`��<ԩD=& m=�\i=��D=�	=�K�<`�[�Դ����"�P���o��   �   ؃��t���p�� �Z;\�<�[=��G=���=ʙ�=^	�=n'�=�:~=�T= T�����D�A�Յ�����G�1����������xV	��� ��	7�yI���U�>?Z���U�"�I��N7�ȉ!��
���h��F���8J�I�
������{K����� ,��Ԏ�<�T=�w�=� �=8��=HX=3!=�@�<�)<���0^B������   �    q��@!�0d�;Xv<���<�,=nGg=���=�ʠ=o��=?N�=K�="=��e�����oF�(��GO
���J��狿Ȍ��������#��@:��3M���Y�"�^� Z�ZM�ʦ:��\$��w�w�迒����ɍ�6N��J�����
P�8�ƽ��¼,��<�X=�O�=�u�=���=��q=��@=l}
=��<�p< �L:�b���   �   Ѓ��\���x����Z;t�<�[=��G=���=㙖=�	�=�'�=�;~=(V=�T�Σ����A�߄��C���
G�����ٌ�����U	�� �+	7�0xI���U�,>Z���U�-�I�N7��!��
�
��Gg��oE���7J���
�����RzK�����0'��,��<�T=x�=� �=q��=�X=d3!=\A�<��)<����]B������   �   x�H�g���@���X�r��^�;�I�< I2=z�n=UӉ=�Y�=�l=�7=�6"��2��`44���������p<�R����˫��*ؿj��n;���-�`�>��3J�!N��J��>�g�-��m��Q��fٿ|/��.���Q?��m�B���O=��⯽�,�����<�D=�!m=^i=��D=��	=xL�< �[�@�������P���o��   �   _0	����W�콡wĽ����4�T���Я$<<d=�uC=�_=��M=R� =`Ʒ�Zʆ�gR�����'��x�+�#7o�����LǿG��=�V����.�e�8�#<��p8�Kc.��\�����:�ǿv�
q�d�-�{�뾁H����&�=;���i^����<��(=�9=��=l�< �9<�μF\V�@����nнMK��F��   �   v{���s�H�`��C�\��h��L|B!���ջ�7�<@Z=@�=8��< 镺��T��G�F�w�>yɾ���uS��2��Z���˨׿f6���f��b���#��{&��M#����-��2��$�ֿ�^���\��n�S�b����˾�1}����/n��n����<L"�<��<�L#<�K���xG�բ���� �,�'��KJ�MOe�h#v��   �   �w;�QȾgȺ�U-���n���_�^2%�=Y۽�Ar������@�;���<P�<`0;4W�+@ѽ��I�2������3�l�o�Ù��!����ٿ.����������/��z��/�['��Eؿxθ��ٗ�_�n�c3�2���\n����L��Mٽ@K,�`~J��>t<puw< @������ڊ����v�.�\�h������̩��m���ɾ�   �   �����u���9 � nܾ�N���H��veH�6��l}�� �漀5���,<��`;x�ü��]�-҃��.˾B��ƐD�N<|�4���l����sͿ{�߿�m뿲�[�꿙N޿�˿�糿����z�{&C����+�ʾj惾�����$�ۼ �Ź�
�;@>Ļ+�4%����
�7wQ�!)��T��FᾪX�,1�����   �   l{]���X��%L���8��| ��H���Ҿ�:��J�Z���	�kA��]�퐻@5�:��O���D���ڽ#xC��Ú�����8�(�G�6�v�r����I�� x��𽿘����%��v������폿ts�:E�1[�l߾�����A�;(ٽ�/F��Rd� SG�`���^���{�����b�����˿׾"
��F#�9V;��N�N�Y��   �   Ò��d����l���{��a\�v�8�!D�7��f)���X�&�����d�ż`������XnѼ�n��>n�d�\�;j��v澿����;�L�_���~�3���1�� ���ɉ��wj��m�{��]\���8�A�N�ᾗ%��X����z��`�ż઎� '���wѼ,s���q�c�\��m��� 澗��2�;�R�_�?�~������3���   �   x���e(��/��7���bxs�=E��]��	߾���U�A�o.ٽ47F��ad� YG� ������u������a������׾+�EC#�KR;�ON���Y��v]�&�X�>!L���8�y �iE�`�Ҿ�6��ހZ���	��:���J�Ð��i�:�O�L�D���ڽ|C�Mƚ����^;�I�G���v�����L���z�����   �   ��P��nQ޿��˿I곿���Nz�h)C������ʾ�胾}���#���ۼ Bƹ��;@Ļ�!�E����
��pQ�+%��?O��c@�qU��-�����������6 �Ghܾ�I���D���^H� ���u����� e�h�,<��`;��ü�ŗ��_�:ԃ��1˾B��_�D��?|�%�������-vͿ>�߿�p��   �   1�F|�71��)��|Gؿ�и��ۗ�M�n��3������p��8�L�DRٽ8P,���J��Ct<��w<  �5��Qӊ�2��M�.���h������ǩ�5h��%�ɾ�q;LȾ�º�=(��j��>�_��+%��N۽f1r�<m�����;ؒ�<��<@1;Z�UCѽ]�I�'4���!���3���o�T���	����ٿ������8���   �   i}&�O#���k��h	���ֿE`��^����S���(�˾5}���4n�`w�d��<�'�<���<pm#<�5��4jG������ ���'�rDJ�GGe��v��{���s�)�`���C�����｢坽�2!�@wջ4J�<�`=h�=��< ���l�T�bI���w�{ɾ��9 S��3����{�׿a8���g��c�!�#��   �   l<�r8�~d.��]���×��ǿ�Þ��q�ն-�����I����&��=���r^�,��<X�(=p	9=8�=�{�< 9�9��μ�LV�E�dнF@��s��n*	���$��FmĽK����3�0���8�$<m=R|C=��_=��M=�� = ʷ��ˆ��S�������羆�+��8o�����<Mǿ���>�O����.���8��   �   
"N�|J�ا>�;�-�Ln�=R��gٿ\0������l?��n�h����=��䯽�0�����<ެD=�#m=�ai=|�D=�	=�\�<��Z�䝳�B��Z|P�0�o�R�w���g��u@����r� ��;@[�<NP2= �n=�Չ=C[�=�l=�8=�7"��3��*54�3��������p<�̏��X̫�`+ؿ���<�[�-�4�>��4J��   �   �>Z��U���I�|N7�}�!�[
�����g���E���8J��
�;���R{K�:����)����<T=px�=�!�=���=�X=(7!=TJ�<�*<`���CB�䋐��u��Xx������-[;��<�`=��G=�À=]��=�
�=�(�=�<~=�V=T�����7�A����q���
G�Ǆ�����X�� V	�K� ��	7��xI�i�U��   �   @�5��42���(��=���e�鿫4��lS�� mh�Z6'�Qg� ύ�L`��ą�����=rDt=i�=���=�r�=���=�}a=6=��=���<���<(Ds<�n<�E�<���<��	=��8=�xl=d�=ٵ�=f�=D@�=��=A˜=n�R=�D(<ZcT�������5Bܾ]$��(e�����q����{�g�_���(��12��   �   F`2��/�׽%����v=�'��h콿�����,d�'�#��ݾ����#�������O�d%=��p=I �=◓=�"�=P�s=LG=X�=HA�<�z{<�*< �o;�SO;��;�K^<0��<x\=��L=�U�=搛=N��=��=Q��=3M�=��Q=�6<$�K�̫�������׾�!�ga�������俄��]q���%�/��   �   �B)��$&�c����M����ڿ�b��Ҏ�F�W����Aо�F�����d�c� ;9��=ޜd=��=�=Rnc=�.2=�<�>X<���� �u�\�̼�^������*�����@�ݻPj<X'�<d�1=>s=���=U��=ܵ�=a��=J�N= �^<�+2���z�w�$˾�#�G^U�����j��4�ٿ��z'�{��{D&��   �   Ph�9��d��9��0����ȿ�u��疂��D����B��g�e�H!����7�٣;��=��N=i[=��A=�v=$7�<g��x���J�u����C�� ��8Z���`����v��}�X�}� 	<��<��J=�Հ=�ƌ=;Ǆ=d.G=��<r��t��N�\�SA��PB
���B�.���D����ȿ2���~��*���   �   �F
�h��T� �z�뿕�п*e��Fi��ff��
,�7W�����<A��Ž�h��}(<~�	=�,=�=<��< �;�μ@�f�����_��0��N-��;�Į>�8�v�'��I�֓�w֝��i1�X�9��q�<�D=R�R=��_=��8=0�<����ɵ��:�%���.��L+��e�┒�,񲿗�ѿL�	=�g��   �   ju�� �}�ݿ(+˿D�������T{y�@�B�Ti�R�ɾ���E���C���ڏ�x)t<���<��<�C�<0�����&��K���m���1��5`�k����֔��ڞ��ɡ��R��ߑ�m���/�U�q�%�p�齗n��|����;D/�<�$=��=�i�<�3�����ȟ�n���QCɾ,~�pOC���z�Z����Ҵ���̿F߿����   �   ��ƿK ÿ����f�������v�{��L�-��ǃ��.���I��8޽
�9�0������<� �<��J<�+C��H���ƽx���_�Pӑ�sݲ��)о��f�����������#�˾"������֢S��e��5��0� ++�<��<�^�<�߿< h[8�@.��(۽��H�������h3�
 N�� ~���(?���湿p�ÿ�   �   r���nu���ᓿ3����l� vF����� �����t�k��*������(����;�Ɠ<��D<�j%��C���ͽ�X+��4|�k���y�پ̈́���='� 1��4�o0��m%��$�Ѽ ���Ӿ�^��d�q���!�]����&��q�����<`��<8<�ˬ�N��� ��S�o��Ĳ�������!�cEI�o�-$��~	������   �   �u�S�p�3�b��M�V�2�/��]-��hRz��L ��밽0O����x�<�[x<��.�ZQ�|�����&����������L���f�5�@JP��d�ӥq���u���p�V�b���M��3��1���)1��:Xz�(Q ���W������<�bx<�M.��H�񖺽�&����������G����5�PFP���d�f�q��   �   �4��0�Yj%��!�� ���Ӿ�Z���q���!�����&��<��`��<H��<<�׬�>���Ғ���o�Ȳ�A�����!��HI�o�X&�������⥟��w���㓿H���El�QyF�������E���;�k�&.�u���h3��P�;Tȓ<��D<0N%�
�C���ͽ�S+�.|����F�پɁ����s9'�+	1��   �   ����̰�7��̯˾k������3�S��`�h-���#���*�ԡ�<�c�<�޿< HN8XG.��-۽��H��㟾t��5�N�U$~�$��iA��鹿�ÿ�ƿ�ÿ󬸿�¨�����ɗ{�LL�g��2��q1��pI��=޽��9�P���̣�<�&�<h�J<�C���G��ƽ���y_�ϑ��ز�*$о羦`���   �   �ġ�N��~ڑ�J�����U�,�%���Of�����0?�;|<�<�
$=,�=�g�<��3�}������v���'Fɾ���QC���z���Դ�0�̿�߿���w�1���ݿC-˿%���!Ø�~y�p�B�k���ɾ�������F�������'t<4��<D!�<�Q�<@���"�&�C��Th�$�1�j.`�*���LҔ�֞��   �   ��>� 8���'��C����%͝�0Z1�8�9���<.L=BS=n�_=N�8=\�<`��3͵���:���B1�N+�^�e�@�����m�ѿW�#>���H
����d� �g��K�п�f���j��bf�Z,�Y�m �F>A�OŽ�k� {(<��	=�
,=F�=\��< y;|μ �f�����T���~�~x-���:��   �   <P��7W��A杽�v��n��}� =	<���<��J=R؀=3Ȍ="Ȅ=�.G=t��< ��~�འ�\�C��yC
�p�B�#�l���ȿ�3����n��'��Qi�2��J�������/�ȿ�v������J�D���	D��)�e�v#���7� ӣ;��=(�N=�l[=�A=�}=�I�<`��P��@�I�����9:��4���   �   x|�4弈����,ݻ��< 8�<L�1=�s=���=�=趤=⍒=�N=�}^<�.2���K�w�i%˾�$�m_U�լ���k��6�ٿ:��(�/��8E&��C)�8%&��c�0��N��x�ڿ�c���Ҏ��W����yBо*G��t����c� �:9�=X�d=��=��=sc=�42=�(�<�aX<���(�u���̼�E���   �   ��O;�0�;�a^<`��<a=��L=W�=4��=R��=���=���=VM�=��Q=��6<�K����������׾-!� a�_��p���:������q���%�k/��`2�</�-�%����=���忹콿9���-d�f�#�<�ݾ䗊�R#�ˤ��`�O��%=��p=� �=ʘ�=3$�=N�s=�G=��=K�<�{< B<�Zp;�   �   �n<�E�<���<l�	=��8=�xl=R�=���=�e�=(@�=i�=˜=��R= B(<8dT�\��뤇�wBܾ�$��(e���������|�t�i��"�(��12�@�5�~42���(��=����H�鿎4��OS���lh�26'�g��΍��_�ą����Z�=�Dt=��=��=!s�=ٚ�=~a=86=��=��<��<�Ds<�   �   @�O; 1�;�a^<���<a=�L=�W�=C��=q��=�=��=�M�=��Q=p�6<,�K�z��ĥ��}�׾d!�a��������J��J��q�H�%��/��_2�t/�q�%�B��=�����뽿���� ,d���#��ݾ���-"�4�����O�j'=��p=^�=��=o$�=��s=HG=�=�K�<А{<�B<�\p;�   �   \|��\���p,ݻ�<08�<��1=s=�=F��=k��=���=��N=`�^< )2� ��<�w�:#˾@#�t]U�����j��h�ٿ ���&�؈��C&�9B)��#&�db���`L����ڿb��Fю��W�!��7@о�E��D����c� �>9�=~�d=��=w�=�sc=�52=�)�<�cX< v���u�$�̼|E���   �   *P��,W��5杽�v��n�X�}� >	<l��< K=�؀=�Ȍ=EɄ=2G=���<,�����d�\��?��eA
���B�fK����ȿ�0�:�����5��Qg�;��q��W����꿘�ȿ�t��ꕂ�u�D�d��@��Ɯe�_���}7���;��=�N=�n[=��A=&=�K�< ����㼠�I����:�����   �   ��>��8���'��C���͝��Y1���9�T��<FM=
S="�_=n�8=�#�<���AƵ���:�{	��L,�DK+�,�e������ﲿ��ѿf��;�G
��E
�A��9� �m�뿼�п�c���g��f��,�hT󾻾��9A�Ž�a��(<��	=^,=��=P �<��;μ�f����OT���~�hx-�q�:��   �   �ġ�N��}ڑ�F�����U�#�%����f�����@H�;4@�<�$=��=�u�<Л3���������@ɾ}|�DMC��z������д��̿�߿���r�K���ݿ�(˿C�������Txy�ȯB�_g�Y�ɾ�������>���ʏ�pFt<��<�(�<XW�< y��l�&�gB��	h��1�9.`����@Ҕ�֞��   �   ����Ͱ�6��˯˾k������#�S��`�-���"� �*�২<�l�<��< hx88.��"۽&�H�Jޟ�>�/1�E�M�x~�.�� =��Z乿��ÿ�ƿ��¿6���)��������{��
L�������+��wI�F2޽��9��L�����<�1�<�J<��B���G��ƽ���y_��Α�uز�$о羟`���   �   �4��0�Yj%��!�� ���Ӿ�Z��׷q�u�!������&��%��`ʇ<��<x8<H�������d��Q�o�;���l���G�!�.BI�`o�"��8��>�����s��Oߓ�����l��rF�$��"��e����k��&���������c�;�ד< �D< ?%�D�C���ͽJS+��-|�����+�پ������m9'�(	1��   �   �u�V�p�5�b��M�Y�2�/�	�U-��HRz��L ��갽�L�������<��x< �-�>����f{&�����й��C���u�5�zBP���d��q���u��~p���b�*�M���2�,����<)���Kz��G ��㰽TC��^����<8~x<��-�JE������&�r��������G����5�IFP���d�e�q��   �   s���pu���ᓿ4����l�!vF����� ������D�k�r*�ߥ���!���I�;ד<�D<P'%���C���ͽrN+�_'|���?�پ�~�=���5'�a1�4��0��f%�9�� ���Ӿ]V���q��!�o	��0�&�P犻hӇ<��<�2<`ì�Ϝ������o�dĲ�������!�YEI�o�+$��|	������   �   ��ƿM ÿ����h�������w�{��L�+������.���I��7޽�9�@l�����<5�<h�J<��B� �G�6�ƽ`��r_��ʑ��Ӳ��о+�nZ��P������C��S�˾�������(�S��Z�E$������)�p��<�s�<x�< 8p8=.�F'۽��H�������[3���M�� ~���'?���湿q�ÿ�   �   ku�� 꿀�ݿ)+˿E�������T{y�?�B�Qi�E�ɾ�����~B��Pӏ��?t<̛�<�/�<\c�<1���&�K:���b���1��&`�󴄾�͔�:ў�𿡾DI���Ց�	���F�U���%���D]�����@��;8O�<d$=<�=�u�<�3�����H��A���2Cɾ ~�eOC���z�X����Ҵ���̿F߿����   �   �F
�j��U� �{�뿘�п,e��Fi��gf��
,�0W������;A��Ž&f�P�(<��	=�,=B�=��<`&;��ͼ��f�]���I���x��q-�e�:�R�>��
8���'��=��}�_Ý��I1�HQ9�P��<:U=�	S=Đ_=$�8=�#�<P���ȵ���:���|.�L+��e�����*񲿖�ѿM�
=�h��   �   Qh�:��d��:��1����ȿ�u��疂�
�D����B��>�e�� ����7���;��=r�N=�q[=b�A=��=�\�<�����㼮�I�����0��U��8F��[M���ܝ�|�u�"_�T}�l	<���<�K=�ۀ=�ʌ=�ʄ=.3G=T��< ������\�:A��FB
���B�+���B����ȿ2���~��,���   �   �B)��$&�c����M����ڿ�b��Ҏ�G�W����Aо�F�����.�c� =9|�=�d=m�=��=xc=�:2=\7�<�X<@K�xu�Dl̼D-���o�h��؉����ܻ@�<pI�<��1=@#s=e��=&��≠�=���=n�N=��^<D*2����N�w�$˾�#�A^U�����j��4�ٿ��z'�}��|D&��   �   G`2��/�ؽ%����u=�)��i콿�����,d�&�#��ݾ����#�N�����O��&=օp=��=���=[%�=4�s=rG=��=\T�<Ф{<pX<�p;@P;p`�;�x^< ��<�e=F�L=aY�=ѓ�=���=⦷=���=AN�=��Q=H�6<f�K����򥄾��׾�!�ea�������促��\q���%�/��   �   �����O�����aTܿ;��\���f�s���6�������S���ܽn���8<ve0=<~=~~�=ݧ�=��=;ć=Xr=RS=��5=��=��=*�=�.=�.=h1=�T=^�}=���=f�=���=��=]��=Ʊ�=Xw�=32�=��=�鍼�?��P�C��<��P���(�3�Q�p������H���ۿ�t��������   �   �:�8��Xy�������ؿG������� o��K3�R���U����M���ս�!�8dK<zk1=��{=��=��=fc�=�x~=�]=,�9=�&=���<hO�<�<���<���<:�=vt2=��_=I�=���=�4�=�w�=�-�=���=C�=V��=�E=(��y&����>�~��������0��l�c햿i5���ؿ-n���u�h���   �   �6����.������6�Ϳ��������Ib��8)�t�Sa���>�l��=�\�<F�3=�:t=���=�˄=��p=AJ=�=$m�<�}w<`w�;�泺"���ל���)�Я�;В�< �=�?=`�{=���=y��=�=D�=,o�=
��=Ҳ=090�X���1����e�}'��i`�a���<���Ϳͺ�������   �   ���62��O�鿠�տ^-��#���̓��7N�����׾kU����&�Uѡ����02�<r�5=��e=v�m=��W=v�+=Є�<@�,<�޻Ԫ��\���jE�J%^�Xa��VM���#�@:м X���TI<�g= Q=Ԉ=���=�a�=�X�=�8�=J�= �`��<���{�,���Ծ}�;!M�H����Pn���eֿ�꿕����   �   �>߿*&ۿ9�Ͽ$��DЧ������6h��4�}��y����o�����t����X	�<��3=�2M=��==~=X[�<p⮻ m����d�j���̟н�1�$�4��;�� v�s������4��[*����<�i =��i=B�=���=&�~=�k)= E�;~tH�&R ��i�ڭ��`��Vx4��h��񎿐{���﾿{пr�ۿ�   �   `"��M���D�����C|��P�r�,�D����V޾�q��-=?���ν���`�;�o�<�+=��'=XM�<��!<�ȍ��L�1i������;T#���C���\��:l��Dp�'uh��kU���8����_sܽ�<��dh��@;�:��<d�D=�zl=X�g=�t/=pan< ]��e�ýL�;�+�����޾�w��E�$Jt�my�����^b��^���   �   hh��KG�����ϑ��2�k��MF��p�����믾7�k��X���W��Lo�<I
=�4=���< �;L�,�}�z�ݽ�4#�x�Y�o
���H���i��]���<𾾗չ��Ѭ��#��z�����J��S�ƺ����;�0��$��<@(=�~E=n�.=�ػ<��K�a󅽊M�+cm�p������<!��|H�(=n�=���ﬔ�0Μ��   �   
~��x��j�=�T�V�9����p��ɻ��E󂾥t(�y%������v;�L�<B�=���<p(1<:��S8��M2񽚮9�<΀�45��sʾM�꾲��\�	������g �ۖ��qľ �����s�T�+�,�ֽhS�`��\�<*=x$=x��<�S�;j��]��6�-��U���ڽ��6��Yu��5<�`\W���l���y��   �   W�A�sH=���1�F� ���
�ֈ�5糾�r���x3�J�սVC� ���J�<dx=��	=�z�<�2���_��4o=�������r�i���&#�5�3��C>��A�L=�E�1�^� ���
����볾�u��J}3�L�ս\C�p<��0C�<w=��	=8��<��1���_���<j=�������z뾎���##���3�B@>��   �   ������ ����Jmľ ���N�s��+��ֽ�[S����*�<
-=$=���</�;>��7��\�-�RX��l޽�;��x��8<��_W�i�l���y�~���x���j���T�^�9�\��Tt��4��������x(��*��t����v;�H�<��=\��<�>1<�(��2���)�&�9��ʀ�
1��*nʾ؍꾽��C�	��   �   "뾾�й��̬��������N�J�SN�%���R�;� c�L�<�(=��E=\�.=�ӻ<��K������P��gm�r������o>!�pH�~@n������DМ�~j��UI����������^�k�;PF��r����T�k��[�����`��xj�<�H
=�6=���<@I�;ܹ�x�}���ݽ2/#���Y����D���d��U����   �   �<p�imh��dU���8�{�-iܽ+4��M��@H ;��<�D=V~l=��g=t/=�Un<h����ý��;�p�����޾�y�r�E�Mt�{�����Rd��g��n$��N���(�������}����r�g�D����OY޾�s��@?���ν�����;�n�< +=�'=@X�<`�!<�����L��`������)N#���C�b�\��2l��   �   0.�)0��,k�	i��߳����H(*�`ʃ<�q =��i=:D�=(�=�~=�j)=P-�;�yH�ET ��i�������,z4��h�5�}��F��|пP�ۿg@߿ (ۿ��Ͽ�%���ѧ�߆���8h���4����S�����o�Q����t�ȓ���<��3=5M=��==l%=�k�<@���$S���d�b�����н�&�d��   �   a��FM���#�tмP���@�I<�p=�Q=׈=���=.c�=�Y�=�8�=�=�a�X?���}������Ծ���"M�<���(���o��Ugֿ�)��������3�������տ�.��$���΃�9N���e�׾|V��#�&�3ӡ�X����0�<ְ5=,�e=N�m=��W=4�+=���<�-<P�ݻ����>��^[E�J^��   �   �����u'���;|��<�=�!?=.�{=࠙=X¯=b�=)�=�o�=���=ȱ=`B0�A����1�͎��g�m'�k`��a���=���Ϳջ�0�����7����4�������Ϳ����B��oJb�79)� u�b����>�?m���?�X�<��3=�;t=���=9̈́=��p=�EJ=�= {�<��w< ��; ��� Ѣ��   �   ���<h��<��=�x2=X�_=�J�=�=�5�=�x�=t.�=<��=0C�=;��=�D=x���'����>�$���o�����0���l��햿�5��Lؿ�n���u�����:�����y����� �ؿ������>!o�@L3�����JU���M�>�ս "��cK<�k1=��{=���=��=Zd�=J{~=�]=��9=�*=\��<�X�<�
�<�   �   /=�.=`1=�T=J�}=y��=U�=l��=��=E��=���=.w�=�1�=0�=덼e@����C��<������Q�3�|�p�����H��3�ۿ�t������������H�����KTܿ�:��E���;�s�o�6�������0S�Z�ܽ���8<�e0=^<~=�~�=���=��=Rć=NXr=�S=��5=��=��=F�=�   �   ���<���<��=�x2=n�_=�J�=��=�5�=�x�=�.�=~��=�C�=Ŵ�=�F=����%��d�>�7���(���Ԙ0���l�&햿5��eؿ�m��Ku� ��W:���	y����2�ؿ���q���  o�`K3�f���ST����M�P�ս^��kK<8m1=��{=��=�=�d�=�{~=D]=�9=+=���<XY�<L�<�   �   �����j'�P��;���< �=�!?=j�{=��=�¯=��=��=Qp�=��=ش=�/0����1�����d��'��h`��`��Q<��R�Ϳ�������i6�`��������>�Ϳ#������NHb��7)��r�0`��C�>��i��h5���<\�3=�=t=i��=�̈́=��p=�FJ=�=�|�<��w<�ö;@����΢��   �   �a��FM���#�мP��� �I<q=�Q=L׈=$��=�c�={Z�=/:�=��=�`��:��Pz�����Ծ~ ��M�y~����.m���dֿ����n����0��ǃ�1�տ,���!���̃�(6N�����׾�S����&�Ρ�����;�<��5=:�e=��m=��W=�+=���<�-<��ݻď������ZE��^��   �    .�0��k��h��ɳ����'*�D˃<pr =��i=E�=M�=z�~=p)= l�;tnH�'P ��i�����#���v4��}h�����-z��	eyп��ۿ�<߿K$ۿk�Ͽ_"���Χ�N����4h��4����1�����o� ��J�t��p�X�<V�3=�8M=��==�'=ho�<P���0P����d�߭��K�н4&�F��   �   �<p�^mh��dU���8� {�iܽ�3��8L�� S ;(��<��D=܀l=��g=�y/=@xn<O����ý:�;������޾�u�ҰE�|Gt��w����z`��^��S ��E��M���D���z��f�r���D���eS޾o���9?�"�ν6�� >�;�|�<<%+=��'=�^�<��!<4���0�L��_�������M#�|�C�9�\��2l��   �   뾾�й��̬��������@�J�>N�񱼽��;�`Z께�<h(=�E=^�.=,�<��K��WJ��^m�����`����9!��yH��9n�u�������%̜�Qf��8E�����􏆿��k��JF�0n����课g�k�WU�}���E��,~�<P
=�;=���<�b�;�ֹ�L}���ݽ�.#�i�Y�a��eD���d��G����   �   ������ ����Fmľ����=�s���+���ֽ�ZS�����/�<�0=�$=���<���;������-��R��I׽�,2���r��2<��XW�ׅl���y�~�
�x��j���T�$�9����bk�����O���p(����0���ew;�[�<��=���<XN1<h"���0���(񽲨9��ʀ��0��nʾ��꾵��>�	��   �   X�A�sH=���1�F� ���
�ӈ�-糾�r��qx3�ڵս�C������Q�<�}=v�	=<��<(�1�ؠ_��Fe=��뉾ƹ���u����� #�V�3��<>��A��D=�o�1�� ��
���㳾@o��Es3��ս�C������[�<�=0�	=���<��1�ة_����i=������jz뾂���##���3�?@>��   �   
~��x��j�>�T�U�9����p������8�vt(��$����� w; V�<0�=���<�`1<P��Q+��3!񽢣9�hǀ��,��fiʾx�����.�	�i�����	 ���lhľʎ��A�s�X�+���ֽ�MS�Ш��<�<�4=V$=���<Pu�;N��(����-�QU���ڽ�d6��Mu��5<�Z\W���l���y��   �   gh��KG�����Б��4�k��MF��p�����믾�k��X�9���Q��,w�<�N
=
==��<0��;�Ĺ��r}�v�ݽ�)#�~Y����@���_��L���澾�˹�Ȭ�'������w�J��H�����6�;��껠�<�#(=�E=$�.=8�<��K��
M��bm�H�������;!��|H�!=n�<�����/Μ��   �   b"��N���D�����D|��P�r�,�D����V޾yq�� =?���ν�����;hy�<�%+=f�'=�g�<��!<����P�L��W������H#�ڳC���\�+l��4p��eh�%]U��8��t�z^ܽ+��,/�� 
;���< �D=�l=ֺg=4z/=8qn<4W��W�ý��;����a�޾�w���E�Jt�ky�����^b��^���   �   �>߿+&ۿ<�Ͽ$��EЧ������6h��4�{��o���ɔo�M����t�����<@�3=J:M=��==�,=~�< 4���7���d�8���x�н}��O(��$��`��^���������p�)�P�<,{ =`�i=lG�=��=�~=p)=�]�;HrH��Q �hi�����U��Mx4��h��񎿏{���﾿ {пr�ۿ�   �   ���82��P�鿡�տ^-��#���̓��7N�����׾_U����&��С�����d7�<J�5=�e=��m=��W=�+=��<�--<0hݻ�w�����KE�^���`��6M�8�#��м����ȭI<�z=�$Q=qڈ=���=�e�=�[�=�:�=V�=��`�$<���{�����Ծt�4!M�E����On���eֿ�꿘����   �   �6����.������5�Ϳ��������Ib��8)�t�La��Ԛ>��k���:��<��3=F>t=��=
τ=��p=KJ=
=���<��w<��; z������2����$��J�;���<*�= )?=��{=���=�į=J	�=��=q�=o��=Ҵ=x30�р���1������e�w'��i`�a���<���Ϳ̺�������   �   �:�8��Yy�������ؿG������� o��K3�Q���U����M���ս6!��gK<�l1=��{=N��=��=ee�=�}~=� ]=�9=�.= �<0b�<��<���<L��<��=.}2=l�_=�L�=���=27�=�y�=r/�=��=�C�=	��=�F=@��7&����>�u��������0��l�c햿i5���ؿ,n���u�i���   �   M����߿�YԿ	`¿N���\����m��E9�~w	������{�(\�e���䅼0��<�I3=�k=Sm�=b�=Z��=�y=vh=�iW=��H=�v>=�-:=�"==�H="%[=�v=��=#Þ=�Ĳ=��=*��= $�=��=M��=2�=@ì=>f=��n<�Z4�q��ej�K������5�6�>�k���F��s$¿qGԿ1�߿�   �   �c*ܿh�п���z����,��6Si���5�'������u�]�8+����k��a�<�R5=�k=�ǁ=Iу=�B~=xm=�yX=b�C=��1=ڳ$=F=�g=��)=��<=��X=<S|=�s�=��=�ͼ=9�=p��=�^�=8��=ˉ�=�1�=h=8��<2%+�4.��"e�n뵾��<�3�U�g�啎�"?��i쾿��п�1ܿ�   �   �տFNѿkƿT~��l��!���2�\���+���������qd������o��I� ��<D�:= �h=y=��t=v�a=v�F=�p'=t8=��<|L�<`j�<�U�<���<���<@��<�R)=�Y=
ʆ=�u�=���=�=D��=���=��=C�=T�l=x�<�v�W�xXU�Y֪�b����)��[�&[���㟿f���h�ƿ�jѿ�   �   �ÿ�S��5��w~��b����x��I�-��\��N���QI���དྷ�:� څ�L��<�A=��b=кe=>�R=r0=��=�A�<�m<�3[�(�O�G��`e���k��` �� ӻ@Q�;Lϯ<��=n�_=t�==�=l�=��=R۽=fO�=�s=`�<�}μ�2���<�]���
�Ᾰ��ԠH�2�w������Ц�c�������   �   ��񬪿q����Z��c��7Z� '0���@pž˃����&�������w(<�=�F=PZV=��F=('=,)�<p��;��1���󼮉B��V���@��X���4��������#�~|:�\�ͼ�%1��e�<&3*=(�v=�֘=���=T˭=ze�=x=H!�<�eP�֖��p�����þAQ�l0���Z��䁿�
������   �   �씿���U����'{�T�[�rn8�������-��$X�FE ��Ir�0�2���<�y'=p�G=��@=R=dȬ< 0ٹ��ҼF�Z������ݽ0������#�Ɠ%�k^���J������?m��[ټ��Y;4f�<BdR=�,�=?r�=���=�_y=B�=��a:��Q��9���OV�E�����8���9��Z]�2�|������d���   �   �@u�h@p�9�b���M���2�s6�9�⋲�T{�U&!��J��� �p��;�n=r*:=|�@=�=��<�/���	�Վ��~߽Y<��A�zd��,��Ї��߉��w��t�u� �V���/�V��|>��$�:�H��t6�<!8=r&t=��=�Ft=��0=x�h<`'�愰���#����.���&�N�s5��oO�1d�q��   �   �A�S=��2��� ������C���߄��n4�ov׽OD�������<� /=`�E=|n/=<��<@��:�������1 �R�7��Hq��k�������&��i̾�mϾ��ɾ*��<��P���P`�W�$�n�ؽ2�f��l�Į�<��*=:�^=��f=��@=�Y�<�|�|�Y�r���=�!���ӹ�vl�4��R#��3��3>��   �   x���0��5�����̾া���=�5��S��i�xIO�`��<j�(=f�O=�3H=��=�?<Df�����k����D�y���𭾋4Ӿ�?��-�S&�Z��z3��8�o��̾�㦾���5�w[�H�i�8jO�,~�<�(=��O=\4H= �=��?<�V��$�������D��u��6�0Ӿ�:��w
�{#��   �   iϾ �ɾ���������
�_�%�$��ؽ*�f�XXl���<`�*=��^=n�f=��@= S�< ��XZ����c�=��#��׹��p뾲��#��3��6>�4�A�)V=��2��� �T�+��+G��Bℾ�r4��|׽"XD��ƕ����<��.=@�E=Rp/=$��<���:��R����- ��7��Bq��g������%"���̾�   �   �ۉ��s���u�A}V���/�2���5��`�:����F�<�&8=V*t=��=�Ft=L�0=0�h<84鼺���b�#����1õ����P�5��rO�`d�iq�Du��Cp�Q�b�҃M��2��8��<����`X{��)!�tO���� �`m�;ll=�):=��@=�=(�<`�.�j�	�XΎ��v߽17��A��d��%��̇��   �   ��%�bX�]~�ç���v/m�|@ټ �Z;�w�<�jR=R/�=�s�=6��=l_y=@�= �`:j�Q��>��xSV����������9�;]]��|�>���>f���<�������*{���[��p8�������3/��[X��G �XPr�h�2��<�x'=�G=��@=&
=�Ӭ< 2չ��ҼZ�������ݽ������#��   �   
�ڷ�����l:��ͼ�a0�tz�<�;*=��v=V٘=Z��=g̭=�e�=vx=��<�uP�Wٖ�a������þ�R��m0���Z�恿sE�������i���Ԉ���[��1d���8Z��(0�R��8ržC�����&������@m(<�=0�F=�[V=d�F=`+=5�<���;��1��~�{B��N��8��Z����   �   �Q��0瀼��һ���;\�<j�=��_=w�=��=�m�=��=
ܽ=�O�= s=<�<D�μ�5��%�<�̍��������Y�H���w������Ѧ�����(���O�ÿU��56�����P���gx�� I�<�����~��HSI�R�� :� ۆ�(��<̜A=��b=��e=,�R=�0=6�=�O�<��<��Z��O��.��(L���   �   D��<���<F =�Y)=|�Y=�̆=Rx�=}��=��=j��=���=���=C�=��l= �<�y���ZU�uת������)�+�[��[��H䟿;���I�ƿ�kѿ�տ'Oѿ�kƿ���������\���+�-���^����rd�T����o��N����<&�:=��h=Dy=n�t=(�a=�F=u'=�==$�<�Z�<�y�<�e�<�   �   ��)=��<=��X=�V|=5u�=�=�μ=�9�= ��=v_�=���=��=�1�=fh=̯�<'+��/��#e�쵾"�ɥ3� �g�G����?���쾿y�п62ܿ���*ܿ��п��ț���,���Si���5�b��j���~�u����+��p�k�Pa�<�R5=k=Jȁ=�у=<D~=Bm=�{X=�C=��1=\�$==pk=�   �   �H=,%[=�v=��=Þ=�Ĳ=��=��=$�=x�=0��=�=ì=�=f=��n<�[4��q��jej����ʢ�W�6�f�k���X���$¿{GԿ6�߿M����߿�YԿ�_¿>���I����m��E9�^w	�����r�{��[����ㅼ���<J3=J�k=qm�=z�=t��=,�y=Dvh= jW=��H=�v>=(.:=�"==�   �   Ƣ)=��<=��X=�V|=Cu�=,�=�μ=:�=@��=�_�=ĩ�=>��=2�=�h=ȳ�<>$+��-��� e�뵾x��3��g������>��쾿��пG1ܿ���)ܿ��п7��	���#,���Ri��5����^�����u����)����k�e�<T5=Dk=�ȁ=B҃=E~=m=�|X=��C=&�1=̷$=j=�k=�   �   ��<,��<� =�Y)=��Y=�̆=ox�=���=��=���=(��= ��=�C�=�l=��<t���JWU��ժ�L��)�)�$�[��Z���⟿������ƿ�iѿ�տ\Mѿ/jƿ|}�����q����\��+�����`����od�3��h�o�P<����<�:= �h=Jy=D�t=��a=z�F=Zv'=�>=�<4\�<{�<g�<�   �   �P��p怼�һ���;��<��=2�_==w�=��=<n�=N�=�ܽ=�P�=�
s=��<�uμ0��K�<�(���p�ᾰ����H���w������Ϧ�>���������ÿ�R���3��P}��V����x�I���T�侾��7OI�e���:� ���(��<ȠA=ܤb=��e=��R=�0=D�=(S�<ؕ<��Z���O�8-���J���   �   �򣽣�����nl:���ͼ�\0�0{�<
<*=v�v=�٘=��=hͭ=ag�=�x=�)�< QP��Җ���遲���þ�O��j0���Z��み�쓿q	������
ﭿo�������)Y���a���4Z�L%0�����mž������&�g�����(<�= G=�_V=��F=f.=t:�<P��;�1�({�,zB�"N���7�������   �   z�%�EX�H~������/m��?ټ��Z;�x�<�kR=0�=�t�=ۂ�=Hdy=F�=�c:�Q��4���LV���<��t����9�!X]�i�|�(��� c��<딿�������%{���[�l8������ᾉ*��G	X�XB ��@r���2�0��<f'=6�G=�@=�=pڬ< �ӹP�Ҽ�|Z�������ݽ�����z�#��   �   �ۉ��s���u�1}V�|�/����5���:�H���H�<l(8=�,t=Ͷ�=�Kt=��0=��h<鼠����#�Q��L�����qL��5� mO�d��q�R=u�=p��b�~M���2�!4� 5����
O{�z"!��D��� �`��;Ju=�0:=��@=��=�/�<�a.�r�	� ͎�Yu߽�6��A�Sd�H%��̇��   �   iϾ�ɾ�����������_��$���ؽ��f��Tl�ܿ�<��*=@�^=F�f=��@=g�< ;���Y���潾�=�O�� й�Oh�ɹ��#��3��0>��A��O=��
2� � �h���� @���܄��i4�o׽�CD��L����<0/=��E=�u/=з�<�+�:h�����- ���7�Bq��g��b���	"��̾�   �   s���0��5�����̾া���&�5��S�*�i�XDO�P��<h�(=֝O=T:H=��=��?<�B����������D��r��q魾�+Ӿ�5����� �����-�:3���I�̾0ܦ������5�zK潠{i�HO�X��<��(= �O=�:H=�=��?< P�������(�D��u����/Ӿ�:��l
�s#��   �    �A�S=��2��� ������C���߄�hn4�v׽�MD�����$�<x/=�E=�v/=��<���:&��!�J) ���7�	<q�*d��I��������˾dϾ>�ɾ��������f�_���$���ؽ��f��)l��ϗ<�*=��^=ʿf=4�@=Hb�<�`绒�Y�2�潐�=�� ��_ӹ�Nl�$��G#��3��3>��   �   �@u�h@p�9�b���M���2�r6�9�܋���S{�/&!�LJ���� � ��;r=H/:=j�@=��=@8�<@�-� �	��Ǝ�bm߽�1��A��d����ȇ��׉��o����u�FvV�N�/�Ƈ��,��*�:��}��Z�</8=(1t=*��=�Lt=��0=0�h<|!鼰���v�#�[��������N�h5��oO�,d�q��   �   �씿���U����'{�S�[�qn8������� -��X�E ��Hr�H�2�`��<�}'=�G=r�@==��< й��ҼppZ������ݽr�� ���#�V�%�0R�vx�ќ�ۙ��Vm�P#ټ@r[;���<sR=�2�=�v�=܃�=�dy=�=�^b:X�Q��8���OV�������)���9��Z]�.�|������d���   �   ��񬪿q����Z��c�� 7Z�'0���<pž����p�&�#��$��((<�=z�F=h`V=��F=2= E�<00�;t1��d��lB��F��1/������飽����(�T\:���ͼ��/�Đ�<E*=��v=�ܘ=��=�έ=h�=x=D'�<`\P�/Ֆ���G�����þ5Q�l0���Z��䁿�
������   �   �ÿ�S��5��w~��b����x��I�.��X��H��}QI���ཤ�:� "�����<�A="�b=��e= �R=�0=L�=`�<`�<@�Y� wO����2��|7��̀��Tһ��;l��<��=��_=|z�=}�=@p�=��=�ݽ=PQ�=�
s=�
�<�zμ2����<�?����ᾰ��̠H�-�w������Ц�b�������   �   �տHNѿkƿT~��k��!���3�\���+���������qd�v����o�F����<J�:=��h=�y=��t=
�a=��F=lz'=�C=��<xi�<���<�v�<��<0��<6
 =4a)=:�Y=�φ=�z�=´�=��= �=&��=Ɓ�=XD�=0�l=H�<�u���JXU�G֪�R����)��[�$[���㟿e���f�ƿ�jѿ�   �   �b*ܿi�п���z����,��4Si���5�'�����
�u�O�+����k�c�<rS5=k=�ȁ=�҃=F~=vm=f~X=��C=��1=�$=�=po=��)=��<=��X=HZ|=�v�=��=м=;�=��=G`�=L��=���=P2�=�h=���<�$+��-��e�e뵾��8�3�S�g�䕎� ?��j쾿��п�1ܿ�   �   ���� ᨿ�ޟ��ґ������W�d.�P���7žk9���M.��,ƽ.0��Բ���<�=~�.=Pk==d�@=��==ү9=�6=޲6=):=�A=��M=.�^=�t=�'�=���=Ǵ�=�=`�=�"�=~��=���=��=���=f��=��=P8�=Կ.= `��Ʌ�<��$�}����d$��,���V�l\�誑�-ӟ�@ᨿ�   �   �
������S��@��Hh{���S��+�r�����Z
���)�k1����%�@l�8�<D�=�_0=T==Z�==��8=v�1=R#,=�)=�)=�.=��8=`�G=��\=&�v=�<�=�=,�=�v�=��=V�=G��="�=m��=2��= ��=���=�+2=@��w��� ���Lx�G���י�z�)�R�R�X�z��%����(����   �   hv�����a����ć��n��LH�ha!�d���ִ���w����誽���@��:�1�<�t=*�4=D%;=0\5=��(=��=�5= |�<8s�<���<��<��=O=��/=^aQ=,5y=���=p)�=T��=fT�=�k�=�+�=�Q�=�g�=h��=��=��;=�4;�sb���p�g��a��4u���G �ŹG�$�m�qЇ����铝��   �   v��
=��@U��. x��Y�s56��H��߾�ܡ��Z��W�}.��4r��h'$<@��<��(=�P9=��5=��$=8�==�<T^�<��W< �;@�m;�D�:��*;P-�;@P<8�<VC	=�-?=�8x=e<�=��=�9�=*��=ʂ�=~��=43�=6��=��I=��< D3��轑_N�蝾)~ݾ����36�KgY��x�E���*d���   �   �݁��~�Ubp��PZ��u>��;��H�������ԉ��A6��ֽ�E����o�<
�=�7=��;=�0*=�N	=�"�<��3<��ƺ��_��ɼ�Z�f����'��$��������Vػh?)<\�<LL@==C�=\��=���=~��=xx�=2ں==��Y=ȷ�<<�J�2T.�D䇾�|��@���I��p\?��A[��-q����   �   v�\��@X�|�K�|�8�WZ �M�\&Ӿu:��Љ]�V�X����Լ��<F=̾4=��D=�F8=X�= ۽< �;�@��K �DJP��J��؝���5ý��ν<Bͽ˓��5E��X�z��.���l��(<
=t�^=Po�=b�=D��=���=�I�=;h=�V�<�ka����ɰ
���^�m���վ��t�!�'�9���L���X��   �   J4�y,0���%�	c�#���Ծ�p��N�t��V%�O2Ľ8�/�@z2����<��/=<`O=�L=�,=|��<h	<�o{���,�>\���ͽǺ��%���-�<8�o9��E1�a �8A���ѽꎽ.��P蟻ĺ�<z@=��=�ә=e7�=$ϕ=��r=$=@��:�91�z�̽`{,��|}�sX���پ�Y��T��'���0��   �   l��	��i ��Z��Iž2���bv��.�qݽf'`���D�\v�<��)=��Y=:gd=zbL=�=��<�5<���4�E�������^�&�T�N�`r�FԆ����q���k>��AG��{b��9���������U�Xi� ��<�-=��s=�Ћ=�g�=H,v=�.=��<�����
���O����=�&���������˾�u��5��	
��   �   �о��ʾ홼����������Ka��W&��Lܽl�n�چ����<N�'="e=�z}=�q=F{B=��< [�P��z��Fh�?�;���t��Օ�+)������̾Qо3�ʾ������������#Qa�b\&�PTܽ6�n�0솼�r�<n�'=�e=$y}=��q=�|B=��< �����t���d���;�*�t��ҕ�q%�������̾�   �   ���:���C��2b�i�9�'�������U� �h�覐< �-=��s=>ҋ=�h�=,v=&�.=�<薧����U���=�����ʹ��t�˾(z�38�
�un�	�l ��^澉MžO����v�@�.��
ݽF1`�XE��k�<&�)=��Y=Zfd=cL=>�= �<�<���4�[���S�����&���N��Yr��І�b	���   �   i9��?1�� �<��ѽ#⎽���p����˿<@=P��=�ՙ=j8�=|ϕ=�r=�!=@M�:�@1�^�̽�~,��}�=[��O�پ�[�W�@'�<�0��4��.0��%�5e����Ծxs����t��Y%�n7Ľ��/�`�2����< �/=�^O= �L=�,=t��<�,	<�S{�`�,�+V���̽V��� �$�-�d8��   �   �8ͽ����x<��0�z�N � �l���(<�
=|�^=r�=b�=���=�¯=J�=�9h=hQ�<�~a�����O�
�)�^��
����վ���s�!�e�9���L�	�X��\�xCX���K���8�@\ ��N�)Ӿ�<��&�]��
��[����Լ �<�|=6�4=�D=XG8=b�=L�< 9�;��?�rB ��>P��C������,ý��ν�   �   ��Җ�4���P�׻�k)<Po�<�T@=�F�=��=��=��=uy�=�ں=ܔ�=t�Y= ��<l'�����V.��凾���������N^?�	D[��/q�@��ށ�6�~��dp��RZ�_w>�=�8K������n։��C6��ֽ�E����i�<f�=T�7=Ƨ;=�1*=Q	=`*�< �3<@�ź8r_�tɼO����&�'��   �   �{�;�AP<��<L	=�5?=�?x=]?�=v��=�;�=���=ރ�=,��=z3�=��=��I=H�<6H3���轲aN��靾�ݾ ���46��hY�Ѡx�6���%e��q�� >��'V���!x�"Y��66��I���߾�ݡ���Z�SY��0��x�� $<T��<�(=�P9=D�5=��$=Ϊ=DD�<�g�<��W<�X�;�<n;@f�: f+;�   �   JU=��/=RgQ=�:y=7��=�+�=>��=�U�=m�=�,�=YR�=Fh�=x��=⺜=��;=�^4;2wb����g�c���v���H �˺G�Q�m�ч�=������w������ ��nŇ��n�uMH�b!����״���w����q骽������:�/�<ht=�4=�%;=]5=��(=ʶ=�8=ă�<`|�<D��<l�<��=�   �   ��\=0w=Q>�=_�=X-�=�w�=���=�V�=���=��=���=P��=���=���=�*2=��ﺅ�������Mx�񟺾C����)���R��z�U&��v�������
���������]@���h{���S��+�������
��^�)��1��>�%�`$l�T�< �=�_0=�==��==p�8=��1=�$,=p)=>�)=��.=��8=d�G=�   �   �t=�'�=���=Ǵ�=�=Z�=�"�=p��=p��=|�=���=N��=���=$8�=h�.=�#`�ʅ�|��v�}����$��,���V��\�򪑿5ӟ�Fᨿ����ᨿ�ޟ��ґ����i�W��c.�6���7žF9���M.�a,ƽ�0��Ѳ� �< =��.=~k==��@=��==��9=@�6=�6=B):=�A=��M=F�^=�   �   ��\=vw=i>�=u�=j-�=�w�=��=�V�=���=��=���=���=^��=��=D,2=���쀀����>Lx�ힺ����,�)���R���z��%���������;
��;�������?���g{���S�+�������	��$�)�0��d�%�� l��<��=a0=�==(�==��8=��1=�%,=`)=
�)=*�.=.�8=��G=�   �   �U=8�/=�gQ=;y=[��=�+�=b��=V�=Hm�=�,�=�R�=�h�=4��=�=��;= �4;qb���*�g�&a��t��+G ��G�&�m��χ����;����u��6������1ć��n��KH�`!����xմ���w�����媽*�� $�:7�<�w=�4=L(;=�_5=��(=�=�:=4��<h�<���<l�<v�=�   �   ���;�DP< ��<�L	=<6?=@x=�?�=���=,<�=��=]��=���={4�={��=��I=��<�?3��轪]N��松�|ݾ���V26��eY�m�x�`���6c��y��<��KT��cx�Y�46��G� �߾ۡ���Z�V��+���h��P7$<��<H�(=�T9=��5=�$=�=8J�<@m�<X�W<0i�;�Xn;���:`x+;�   �   ��
�����P�׻0m)<p�<�T@=�F�=\��=r��=���=Dz�=�ۺ=���=��Y=���<����Q.��⇾�z����������Z?��?[�}+q����܁���~�`p�pNZ��s>��9��E������Ӊ��>6�)ֽ:�E�@��x�<��=��7=��;=`6*=@U	=2�<0�3< vź�f_���ȼ�L����Ԏ'��   �   q8ͽ?���(<����z���@�l���(<^
=�^=wr�=�=���=�ï=�K�=�?h=ta�<�Qa�憊��
�>�^�8��a�վ`����!���9�"�L���X���\�l>X�
�K�4�8�IX �RK�]#Ӿ8����]�Q�aS����Լp�<��=��4=��D=�L8=D�=@�<�Z�;0�?��> ��;P�bB��񔬽,ý�ν�   �   �h9��?1�� ��;�I�ѽ�Ꮍf�����TͿ<@=���=}֙=�9�=�ѕ=Ĉr=�)=@��:�01���̽�w,�x}��U����پ�W��R�h'�#�0��4��)0�+�%��`��$�Ծ�m��p�t��R%�8,Ľ��/���1���<f�/=�eO=
�L=X,=l��<?	<�B{�t�,�hT����̽���L ���-�8��   �   �𐾸:���C��b�R�9���`���nU���h����<F�-=��s=�Ӌ=xj�=�1v=�.=$�<�x�� ���H����=�w���l�����˾�q뾝3�D
��i�F	�g ��V�Fž؈���v���.��ܽ�`���D�t��<V*=��Y=2md=�hL=��= �<�
<���4�{���������&�4�N�LYr��І�;	���   �   �о߇ʾ♼�韧�����vKa��W&��Lܽ޳n��؆�Ȃ�<��'=�$e=�~}=<�q=��B=\��< ����	n���`���;�M�t�2ϕ��!��o��k�̾�о��ʾ�������D����Ea��R&��Dܽ�n��Ć����<��'=\(e=̀}=�q=��B=���< ������r���c���;���t�Tҕ�<%��h����̾�   �   �k��	��i ��Z��Iž)���Qv��.�0ݽ�&`���D�Dy�<
�)=��Y=�kd=�hL=�=��<�;���4����������&���N�=Sr�L͆�����쐾7��C@���b���9�
������ U�P�h��<��-=\�s=.Ջ=Sk�=�1v=�.=4�<������.N��B�=�ء��_�����˾�u��5��	
��   �   F4�v,0���%�c�!���Ծ�p��:�t�pV%�2Ľh�/��g2�X��<<�/=$dO=��L=2,=,��<�O	<�){���,��N��s�̽t��k�L�-�E8��b9��91�� ��6�ٹѽ�َ�z���0���߿<R!@=���=xؙ=;�=ҕ=��r=8(= M�:t61��̽�z,�|}�4X����پ�Y��T��'���0��   �   v�\��@X�|�K�z�8�UZ �M�V&Ӿo:����]�8��W����Լx�<b�=��4=�D=�L8=Ģ=H�< ��;��?�L6 ��0P��;��h����#ý��ν2/ͽ���S3��.xz��@el���(<�!
=��^=cu�=:�=��=�į=aL�=?h=�]�<`a�ŉ��4�
�1�^�3����վ���e�!��9�{�L�}�X��   �   �݁��~�Wbp��PZ��u>��;��H�������ԉ��A6�NֽX�E�0��Lr�<l�=��7=b�;=>7*=<W	=�8�<8�3<��ĺ�F_�D�ȼ�A������'��P��t߫���׻8�)< ��<h]@=gJ�=:��=���=K��=|{�=�ܺ=ږ�=�Y=��<��J��S.�䇾�|�����=��f\?��A[��-q����   �   v��=��@U��/ x��Y�q56��H��߾�ܡ���Z��W�?.���p��0,$<��<�(=T9=<�5=4�$=.�=�P�<�u�<��W<���;��n;���: ,;���;`kP<��<BU	=J>?=*Gx=�B�=H��=J>�=���=���=���=�4�=���=D�I=X�<jB3�;��@_N��睾~ݾ����36�FgY�
�x�D���*d���   �   hv�����c����ć��n��LH�ha!�c���ִ�z�w�����窽4�����:�3�<�v=h�4=V(;=4`5=�(=�=�==��<���<���<<'�<N�=
\=^�/=�mQ=�@y=���=.�=_��=�W�=�n�=.�=�S�=Xi�=���=��=h�;=`�4;�rb�j�;�g��a��#u���G ���G� �m�pЇ����蓝��   �   �
������S��@��Hh{���S��+�q�����W
����)�W1��B�%�@l�D�<�=�`0=�==`�==�8=��1=',=�)=�)=j�.=��8=��G=ھ\=fw=�?�=��=�.�=y�=��=�W�=���=I�=[��=���=���=2��=D,2=���2������Lx�=���ә�v�)�O�R�W�z��%����'����   �   �x��Qs���e��P�m�5�d�wn�ι�������7�X��Rj��Pr��(�����;x�5<�Y<p�Z<PyU<�)\<�zz<�V�<4j�<8C�<b0=��<=�;`=���=�i�=���=��=���=�<�=l��=��=��>8c>��>���=��=��=���=<1�<|�������V����z�C���+�����sK5�PP�t�e��Rs��   �   F�s���n�6�a�<�L�Nn2��"�\x˵������2�kH὎�|��7�p�ɻ0&�;��L< ^k<�~g<X�[<P�Z<h�o< #�<��<��<&�=�1.=�<P=R't=�Ҍ=�3�=�ٳ=�4�=}��=���=���=Ř >��>�c>5�=��=�=,m�=2=(�u�X������u�������� ���1�6�L��a�7�n��   �   l�f�S!b�LPU�QoA��g(������)��եt�0�$��%˽>Z�09���K���7<��<O�< (�<��j<��Q<rL<0_<��<�n�<���<��=h#=�f@=�e=�d�=�I�=g��=~+�=/�=�q�=��=��=�M�=�=s��=z:�=2��=�T=x�%����A��G5e�sa��"hݾh��5>(��A��{U�8Ab��   �   $WR��$N��AB���/�����-�ɾ9
���X�4g��z��^�#���*�@<ٗ<h��<�o�<���<�~x<�q8<�u<���;Ј�; �;�<�fM<T)�<��<@
=�3=8b=Ȧ�=�g�=$�=|��= �=���=�}�=�=�u�=�=��=��=`]7�fc������L�s���Ⱦ]����OZ0���B�@fN��   �   O�8��4��*�a�������۾�D�����ĳ3�佪|x������S;,$�< ��<���<L��<���<H�u< .�; %+:pV��@�0��fm�L텼d�����V��~�� Bw:��C<�U�<C"=�.`=�T�=Z�=�S�=\��=>��=Y��=���=�k�=��=P�/=���;��(��z̽�-.�L���?>����ݾ/ �ј���*�P-5��   �   ���������~ �Aݾ�����N���_N� �
�&���p�� Pg�d��<E=��=�=��=<�<�Q< k�:h�7��C��r��q4��cR�n�c��e�$;U���3��� �d��� y";��<̕(=`r=[2�=S�=���=��=���=�^�=ސ=�RA=�y<��Ӽ���ړ���S�<��t����*�4(�@��Ǿ��   �   ����T�����e�̾�	���ۍ��QX�.��ᓿ�T�@� (����<�B=v�5=�,@=D�1=�R=|ֹ<���;HZ#����VD��}��¡��>�Ƚ�ܽm��EL�eZѽ�鳽*���|9�tk��0��;0��<��M=�ى=m�=�.�=��=1֧=b��=�N=\��<P"4�l�[���ս�&���f��̔��3����Ѿ�辌����   �   K���|��CV��W����?���N�!����ǽx�V��	n� �z<&�=�%N=F�f=2�b=BiF=��=���<@H캨�ԼP%W��줽�i޽�5
�va!� �2�<���<��3�"�����'ս���������̧<K2=(�y=���=�=�Q�=�7�=�U=��<�r;rS�N�����x.�^c��)��᪡��,������   �   	����,����x�l4Y��`2�����Y����K���d�P�<L%!=H�c=�]�=��=��~=HuR=*�=��H<P�y�L�A��Q�������$�0�J��l�Uׂ�Uq��3����/����x��9Y��e2�$���`��L���d�`A�<�!=ސc=�[�=�=P�~=�tR="�=��H<��y���A�M��u���}$���J�pl�jԂ�?n���   �   3�<�ٻ3��"����yս�z�����@��0ݧ<�Q2=0�y=���=|�=�R�=M8�=ZU=p��<�;;�X�N�����{.��bc�0,��䭡��/��������������Y��_����B����N������ǽ|�V�X)n�(�z<B�=�!N=v�f=L�b=bhF=��=���<���@�Լ�W��礽yc޽�1
�]!��2��<��   �   �C��Qѽ�᳽���9��S����;��<n�M=I܉=� �=20�=�=�֧=���=�N=���<�24��\�;�ս�&���f�dϔ�n6���Ѿ���K����������<從;a��]ލ��UX�q�����t�@��5(����<�>=b�5=H*@=��1=`R=�׹<���;K#�<�꼐D��x������3�Ƚ5�ܽ���   �   �-U�@w3�� �D����'#;��<�(=�fr=.5�=FU�=���=��=z��=b_�=�ݐ=NQA=(y<��Ӽ���4����S�@�����-��)�
�����m������ � ��Cݾ%����P��cN���
�!ţ������g���<�A=H�=R�=��=t�<HQ<���:(�7�L8������g4�YR�Jwc��e��   �   �-����y:��C<h�<tK"=�5`=�W�=�=�U�=��=���=L��=��=�k�=[�=ď/=�v�;r�(�H~̽�/.�ϓ��*@����ݾ��]��n�*�/5��8���4�-*�ܙ������۾�F�����3���N�x�t���`�R;@�<@��<���<���<м�<��u<@:�;��+:06��h�0��Km�P݅�L邼�YV��   �   0�<n
=�3=�"b=ʩ�=Tj�=t�=p��=V��=:��=�~�=��=Bv�=���=͗�=��=��7�0jc������L��	����Ⱦc�����[0��B��gN��XR�T&N�ICB���/��������ɾn��tX��h�;}����#�h�*�P6<�ԗ<��<lm�<L��<�~x<�t8<�|<�	�;0��;�3�;H�<�M<7�<�   �   Lk@=e=�f�=�K�=]��=A-�=�0�=�r�=��=���=N�=~�=���=k:�=߯�=�S=8�%�����h���6e�wb��giݾ,��?(�چA��|U�JBb�~�f�]"b�BQU�.pA��h(�����ྯ*�� �t�.�$�Q'˽�Z�0=������7<\�<0M�<'�< �j<��Q<�uL<�#_<|��<�t�<���<̊=�'=�   �   �)t=�ӌ=�4�=�ڳ=�5�=X��=���=H��=� >Ŀ>d>15�=��=Ϯ�=�l�=H=؎u�b��X���u�����h��m!�h�1���L�y�a���n�֐s�v�n���a���L��n2��"��x��˵�A���%�2�I὘�|�\9��ɻ0 �;�L<P\k<(}g<0�[<P�Z<P�o<�$�<�< ��<��=�3.=0?P=�   �   ���=�i�=���=��=���=�<�=p��=���=��>4c>��>���=��=���=x��=D0�<�������������z�i���U�����K5�&PP��e��Rs��x��Qs�t�e��P�Y�5�N�Pn�\ι�������7���j���q��������;��5<HY<��Z<�yU<*\<@{z<W�<�j�<�C�<�0=ҵ<=�;`=�   �   (*t=Ԍ=�4�=۳=�5�=u��=���=a��=� >п>-d>f5�=n��=<��=�m�= =(�u����4��,u���1�꾲 ���1�˅L�l�a���n���s�[�n���a���L��m2�"��w��ʵ�r����2�G�l�|�4�`�ɻ01�;(�L<dk<��g<`�[<@�Z<��o<�'�<��<���<�=�4.=�?P=�   �   Nl@=�e=Eg�=1L�=���=h-�=�0�=�r�=G��=��=�N�=��=>��=@;�=��=�V=��%�p��@���3e��`��gݾ���s=(��A��zU�0@b�Y�f�@ b�?OU�SnA��f(�=�f྿(���t�Ȱ$��#˽�Z�3�� ��0�7<$�<�T�<@.�<�j<0R<��L<@/_<���<ly�<���<\�=)=�   �   ��<�
=��3=t#b=��=�j�=��=���=���=���=�=V�=w�=,��=w��=��=�7�>ac�
����L�7���Ⱦ�����Y0�T�B��dN��UR�e#N�~@B�0�/�������a�ɾ���4X�Te��w��|�#���*�(O<L��<ؼ�<�w�<d��<��x<ȇ8<p�<�)�;0ø;�L�;��<��M<�:�<�   �    !�� z:��C<�i�<L"=z6`=,X�=F�=LV�={��=��=��=��=Jm�=_�=j�/=p��;��(�w̽+.�Đ��]<��]�ݾ���T�� �*��+5���8�Q�4��*�̖�3��D�۾�B������3��佚ux������gS;X-�<��<���<h�<�Ȳ<��u<�f�;�$-:���h�0��<m�ׅ�$䂼@QV��   �   �+U��u3��� ������2#;� �<��(=vgr=y5�=�U�=&��=��=���=�`�=-��=�WA=x�y<T�Ӽ����j�S�&
�������'ᾓ&�y���������#���| �>ݾ���gL��4\N�,�
�j��������f�� �<2J=�=v�=��=�&�<*Q<��: �7��-��F���c4��UR�|tc���d��   �   �B�1Qѽ3᳽&� 9�`R����;D��<�M=�܉= !�=�0�=9	�=sا=��=^�N=<��<4���[��ս9&�d�f�mʔ��0����Ѿu�达������}���	���̾}��Hٍ�{MX�������@���'�辉<�H=��5=(2@=:�1=tY=��<@(�;2#�p��FD��v��������Ƚ��ܽ����   �   В<���3��"����)ս�z��H����ާ<LR2=Z�y=���=��=JT�=�:�=�U=d��<��;�I�n��}���s.�Yc��&������)��e𽾛���xx���R��#���=���N�����ǽ�V�H�m��z<��=�+N=�f=�c=�oF=��=$Ɯ< �0�ԼHW�?夽@a޽�0
�A\!�z�2�Q<��   �   �����,��n�x�E4Y��`2�ښ��Y���K�H�d��Q�<P&!=��c=�^�=���=��~=�zR=��=��H<��y�J�A�JF������sx$�b�J��l�Pт��j�������)��j�x��.Y��[2�|��>R����K���d�xa�<�,!=��c=k`�=ᵈ=x�~=�{R=x�=H�H<X�y�,�A�~J��0���
|$���J��l�#Ԃ�n���   �   +��� |��1V��I����?����N���F�ǽ�V� n���z<^�=n'N=̔f=��b=FnF=��=dȜ<���Լ�W��ऽW[޽#-
�X!���2�2
<���<�?�3��"�����սs������b���<FY2=��y=� �=)�=^U�=;�=�U=��<`�;`N����`��w.�9]c�3)������L,�����   �   ����D�����Z�̾	���ۍ��QX���������@�@(����<"D=��5=�/@=��1=�X=D�<�5�;(%#�l���C��q��쓫���Ƚ0�ܽ���7:⽕Hѽ�س�c鋽
�8��9���]�;$��<d�M=�߉=t#�=�2�=�
�=H٧='�=�N=���<4�&�[���ս�&��f��̔�O3����Ѿ��m����   �   ���������~ �Aݾ�����N���_N��
�������� Cg����<�F=0 =|�=��=$&�< -Q<���: �7�X#��Z��[4�NKR��hc��d��U�|h3��� �~��`�#;�4�< �(=�nr=r8�=X�=��=
�=���=�a�=W��=�VA=��y<P�Ӽ�����#�S����5����*�!(�2������   �   M�8��4��*�_�������۾�D������3���4|x�\����%S;�&�<���<���<���<�ǲ<8�u<0p�; �-:@󷻰�0��#m��ǅ��҂��+V���� �|:��C<0|�<�T"=
>`=t[�=�=�X�=T��=���=��=���=�m�=a�=��/=��;�(��y̽�,.�
���>��q�ݾ �Ę���*�J-5��   �   $WR��$N��AB���/�����)�ɾ5
���X�%g��z����#��*��C<�ۗ<<��< u�<���<x�x<��8<��<`<�;0ݸ;�n�;�
<��M<�G�<�&�<�"
=��3=*b=��=Jm�=�=���=I��=���=��=�=�w�=o��=o��=��=�97�
dc�0�����L�F���Ⱦ?����FZ0���B�<fN��   �   j�f�T!b�KPU�PoA��g(������)��ϥt�%�$��%˽�Z�T8�� &�8�7<P�<XR�<�,�<��j<�R<��L<`4_<t �<x~�<���< �=0-=�p@=X e=zi�=EN�=���=,/�=;2�=Lt�=e��=֘�=�O�=l�=���=j;�=��=pV=��%�_������5e�Xa��hݾ_��.>(�݅A��{U�7Ab��   �   G�s���n�6�a�;�L�Mn2��"�Zx˵������2�cH�^�|�7� �ɻp)�;ؖL<pak< �g<`�[<�Z<��o<�(�<X�<���<Z�=<6.=�AP=0,t=Ռ=6�=#ܳ=�6�=K��=e��=��=V� >�>`d>�5�=���=c��=�m�=�=`�u���|���u�������� ���1�3�L��a�5�n��   �   My)�v&�tG��#��p����ʾ溠�^Ts���/�$��������P��������] �|K�%���+�X�$��#��/ҼH�a� ��8`v<��<�d9=�s=e��=	�=΅�=d��=���=>�=��>]>��	>�U>�F>\��=���=I��=�~k=���<(��� ������a�	1��M�Ǿ���3��e8�&��   �   �@&�y�"�n?��X
�rx�lƾL#���nm���*�|�˅����E�z���BԼ��Ѽ���P���&��'%���8�
�5мp�g��h�(]<�r�<�p/=��h=٢�=��=޳�=��=��=̿�=C�>b�>	q>7;>Xn>��=�'�=&{�=r�l=� �<T���_=�����d5\����+�þ�B�^*
��?��"��   �   ������Ut�	@���������RS\�6��eӽ᳆��I%�0�мx��ޜ��h���o漪��~-��;��X�L�̼��}� #��P�<���<Ң=n�F=�={=��=^��=�]�=2��=.�=�>�=N�>JE>>�>���=���=���=��=�{p=_�<�-��XB��r��86N��㎾�N��Ŧ�R\�ߤ�6���   �   �Y�$K�����F���ʾ����Ay��{�A�;9��쯽xKR����Ȫj�f�R�( Y�=����ʼ���8:��h��(�ͼ�R���&� ����,<�g�<��
=Z�<=��n=�t�=���=
��=z��=�0�=�N�=|U�=�=�Z�=���=\�=X�=t=��<�0��ap��콺�8��׀�`���r�˾���F�!���   �   c���w;����]˾O2�����p�[����_$׽P������8
D� �ζ`4�;`�d;@䭺N�hx�\����м���T޼,3ʼ����@Vk�p���$�:h�E<�w�<\J=��G=�l~=��=���=�k�=,��=p��=("�=ؠ�=[E�=^�=��=��v=��= �^�z�=��ƽ�d���^�"ϐ�9��ξ[��xP��   �   ��ξyɾ�񻾲���3F��Ne�0S-����K��0���E@����;���<�,�<�9�<��><`�i;Ͱ��hg������3弈�lE����H���F���ּ(���i�����;�<��=0JO=Ո�=�[�=ǅ�=U��=�z�=��=�u�=��=�)�=.t=H:=�	r;
�w���f��\�8� Yq�}���N��cU���:˾�   �   hp�������ړ����N�Z���+�����
z��r�,�(GC���-<@'�<j�=
�= �=�G�< �n< /N;��<�������o.�~�S�_q�7����Y�����@)n�N\F��N��w�� <�8���<��=�1e=��= ��=���=�U�=��=��=ɶ�=��j=��=��<0���:�p�k̽�����@�(�l��鉾����^%���   �   -�w��ln�%pZ���=��q�<;��M����&��&�X�n<��=��6=��M=��L=Hm8=�=�z�<��< ڻ!¼�(�\�o��ݙ�!���Cн-��X�X�޽��˽u����݅���.��e��Х�;X��<�7A=��="ҕ=U��=��=�U�=�Ǉ=2�W=��=�0M<(v\��/��R��������v5��R�z�h���u��   �   �l.��8%�|�|=���
������T��J��8a�<ā"=�)]=V\�=���=�V�=�Vh=�:=�N�<��N<�(��S���c��饽^ٽ�������'�"/�Uq.�R=%���6E������"��`_�0����R�<�{"=�$]="Z�=ݷ�=U�=�Sh= �:=L�<�N<x$�`N��H�c�楽PYٽ������Ҁ'��/��   �   ��޽9�˽W���6ׅ���.�lP����;ؒ�<j>A=N�=hԕ=C��=4�=W�=�ȇ=��W=��=.M<�~\��/��U����ཟ���y5��R���h�R�u�(�w��qn��tZ��=��u��A轋S��<�&���&��n<�=�6=f}M=�L=j8=0=�v�<��<~ڻ�¼��(��o��ٙ�a��>н�ཱིQ��   �   Zn�LPF��B��a�� D�8P��<\�=X8e=��=W��=p��=fW�=��=��=���=p�j=��=��<T���4�p�̽I��	�@���l�)쉾8����'��s��B���^ݓ�N���^�Z��+������~����,� bC���-<h�<�=�=|�=A�<��n< N;h��h������(l.��S��Wq������T��]����   �   �������@G�;dў<��=dQO=���=�^�=��=B��=�|�=	�=�v�=��=>*�=F.t=x9=@�q;�
�>���\����8�K\q�u	��Q���W��G=˾��ξ�{ɾ>�������8H���e�V-�ٽ��O�����x[@�0[�; z�<�$�<�1�<�>< oi;�߰� og�����p2�Z��A��������>�|�ּ�   �    �E< ��<LQ=��G=�r~=s�=��=�m�=���=���=e#�=ڡ�=F�=��=V��=��v=��=��^�T�=�ݺƽ�f�-�^��А�c;��(ξ����R������=�
���_˾.4������[�Ͻ��'׽A�������D� @&���;�d;@N�� Z�xx� ����м�ἰR޼t.ʼ����`Ck������:�   �   ��
=\�<=��n=0w�=è=��=E��=2�=�O�=�V�=\�=�[�=@��=�\�=X�=>�t=l��<(0�.ep����x�8��؀�¼���˾ކ��G�.���Z�,L����dH뾄�ʾ����Zz��I�A��:�ﯽ|OR����طj�xr�@^��Y�hB��<�ʼx�켨<��|��\�ͼ�O����%� s��h-<xp�<�   �   ��F=�@{=N�=���=n_�=���=T �=�?�=��>�E>��>$��=���=���=��=F{p=�\�<�1���C��x���7N�y䎾�O�� ��]����������S��u��@�����l����T\�9���fӽE���TL%�� Ѽ�|���✼�l���s�`���.��<�HY��̼��}����P�<���<��=�   �   $�h=���=\ �=���=D�=���=_��=��>��>1q>Z;>qn>5��=�'�={�=��l=$��<슯�O>�����66\�?��ɲþsC��*
�$@���"��@&���"��?�Y
��xﾃlƾ�#��Hom� �*�>	�n���ζE����PEԼP�Ѽ\��`���'�r(%�t��x�
��4м��g� �g�x]<@u�<`r/=�   �   <�s=v��=�=څ�=j��=���=>�=��> ]>��	>zU>�F>F��=���=*��=\~k=���<0��!������a�%1��k�Ǿ���A��n8�&�Ly)�r&�kG��#��p��ߴʾʺ��.Ts���/�������z�P��������] �pK�
%���+�:�$�z#�L/ҼP�a� `�8Xv<L�<�d9=�   �   ��h=���=� �=ش�=d�=���=���=��>��>Aq>l;>�n>u��=D(�=�{�=B�l=��<�����<��t���4\�a����þ6B�*
�_?��"�(@&��"�?�iX
��w�lkƾ�"���mm���*�9꽾���ֳE���@Լ �Ѽ����$��%%�ȓ���
�L0м��g� qg��]<�w�<js/=�   �   �F=(B{=��=D��=�_�= �=� �=�?�=ϫ>�E>��>~��=`��=h��=���=�}p=�c�<T(���@��f���4N��⎾�M����ྯ[�-��v��5��˪��s�P?������������Q\�����bӽ����F%�\�м�r���؜��b��`i� ���)�t7�vT�\�̼��}�����ȝ<T��<��=�   �   ��
=��<=�n=�w�=xè=\��=���=L2�= P�=�V�=��=�[�=���=�]�=fY�=̈t=(��<��/�l\p�����8��ր�����ٖ˾5���E���|X�J�����D�4�ʾ"����w��P�A�r7��鯽rFR��传�j�`V�0B�P�X��3����ʼ �켐.����,�ͼE����%� x���-<�u�<�   �   �E<ԉ�<�R=��G=�s~=��=Y��=�m�=D��=H��=�#�=n��=�F�=��=࿧=�v=�= y^���=��ƽ_b���^�q͐��7���ξ����M������8�?�⾇[˾@0��&��]�[���' ׽Ι�����@�C�  ŵ�Z�;�e;�=��87�x�w�����м��D޼�!ʼ<���x0k�p�ỀW�:�   �   d������ T�;�Ӟ<��=&RO=R��=�^�=d��=���=�|�=�	�=�w�=��=�+�=�2t=�?=�sr;R
�͒������8�8Uq�T��sL���R���7˾.�ξOvɾ﻾;����C��oe��O-����oG�����P+@�@��;���<X7�<�D�<x�><@j;P���0Ig�@���$!�n���:��������:���ּ�   �   �n�>NF�dA�4_�� <�8�<
�=9e=��=���=���=X�=��=��=N��=H�j=<�=@<����(�p��̽c����@���l�}牾����"���m��؄��7ؓ������|Z���+�&���{t��2z,��'C���-<`3�<4�=��=�=hT�<��n<��N; ��̓�� ��$d.��S��Qq�)����R�������   �   ��޽?�˽�����օ���.��N��0��;��<?A=�=�ԕ=校=�==X�=cʇ=N�W=^�=XPM<�Q\���/��L��ɖ�����q5�B�R�]�h�*�u�ʿw��gn�kZ��=��m��3轊G���&��&��n<6�=��6=V�M=��L=Zs8=��=���< �<4ڻ0¼0�(�p�o�f֙�q���;н��P��   �   jl.��8%�*��<��7
��n��TT�0F��xb�<|�"=�*]=�\�=���=�W�=�Yh=h�:=XZ�<��N<����9����c�kߥ��Qٽ���3��"|'�
/�h.�*4%����5�� ����dI�����q�<��"=P0]=@_�=���=�Y�=�\h=��:=�]�<��N<��>����c��⥽GVٽj������'�2/��   �   ��w��ln��oZ�^�=��q��:轖M��4�&���&��n<T�=��6=��M=��L=�o8=��=0��<x�<�6ڻ�	¼|�(���o�ә���36нd�߽,I�r�޽��˽i����υ�x�.��8���@�;T��<�EA=��=Vו=�=��=�Y�=�ˇ=��W=:�=�OM<PX\���/�rO��������t5��R���h���u��   �   <p������ړ�񊂾0�Z�k�+������y���,��DC�`�-<�(�<��=��=h�=�M�<��n<@�N;���ȓ�����
a.��S��Jq������M��$����n�JBF��5��H�� ��8(��<�=�?e=��=0��=�=�Y�==�=�=,��=T�j=v�=�<����F�p��
̽�����@�B�l��鉾{���#%���   �   ޽ξ�xɾ�񻾢���&F��6e�S-�׸��K�����PC@�0��;p��<0/�<=�<��><��i;����HPg�쐲�p 弸��~7����Z~�43���ּX攼�������;x�<��=zYO=���=�a�=���=���=�~�= �=y�=��=�,�=�3t=�?= ^r;
����M��b�8�,Xq�%���N��*U��w:˾�   �   O���j;����]˾G2�����\�[����6$׽$��� �� D�  ���<�;`�d;����hC��x������м�ἼB޼�ʼ ���Xk��v�  ;`�E<���<�Y=B�G=�y~=��=ֹ�=,p�=��=���=)%�=���=�G�=��=L��=<�v=
= �^���=�?�ƽ�c���^��ΐ�>9���ξ6��]P��   �   �Y�K�����F���ʾ����;y��n�A�,9��쯽KR�̫优�j�c�PN���X�D9����ʼ�켄1�����$�ͼPC��x�%� ��`*-<~�<*�
=̝<=��n=z�=�Ũ=`��=S��=�3�=zQ�=�W�=��=�\�=���=,^�=�Y�=܈t=��<8�/��^p����&�8�j׀�+���I�˾���F����   �   ������Qt�@���������HS\�-���dӽǳ���I%���м$w���ܜ��f��Pm���J+��8�2U���̼��}�p����<h��<�=ںF=(E{=G�=���=a�=��=�!�=�@�=D�>F>��> ��=���=���=��=�}p=�b�<<*��|A�����5N�v㎾�N�����H\�פ�/���   �   �@&�x�"�n?��X
�qx�lƾK#���nm���*�v�����v�E�N��dBԼX�ѼD��¶��%��&%������
��0м��g� bg��]<py�<rt/=,�h=���=N!�=���=�=���=��=Ћ>޲>oq>�;>�n>���=l(�=�{�=h�l=��<t����<�����65\�����þ�B�[*
��?�~�"��   �   7پ��Ծ�8Ǿtв�إ���|�>G�z<��L䦽R��Ryn�@oy��[��������˽�~�����A� �Y����]���ýn��h�N��μ �i�|{�<�n9=槄=>��=���=�y�=�Y�=9V>$<>J�>5!>��>��>���="��=���=s�=$�P=hd�<(��2-���,���t6�,s��n��5���[	Ǿ5�Ծ�   �   ��Ծ5.оb
þ��b0��c�v��B�����ؽrK��`�|�n�b�n�m�>=��M9����Ľig�`��9��X���_$�m���z�����K��]μ 2I�h�<��3=7�=4��=��=X��=j��=�� >��>�~
>��>�
>8�>pE�=lx�=���=�Ý=�P=��<th��,v��ڙ��2��n�`���f���þ�Eо�   �   Ⱦ$�þ�붾_���)��}:e�_3�,�P�½����aY� �@�4�K���p�i�������˽lV߽������oFѽ��������D���ϼ�X.��Ĝ<w!=�m=O_�=M6�=T �=T��=L�=�>`>�B>6|>g�>&��=<��=�
�=by�=|�O=(š<f��N�y�3��K�'�s3`��������z����þ�   �   �3��Qү�����S���y���I�h���e�.v����]��"�P��H���$9�vl��Y������,���ʽvȽ�'�������ƃ�F=�Ȱټ ٻ��R<@� =�BG=�%�=��=*��=���=h��=Ȇ�=L��=B�>X�>��=ܕ�=T��=LH�=�ݖ=<�L=���<�\�� [���ɽ{���VJ��|�
5�����������   �   V������P��ǝx�\�Q��W'�u���ؗ���oi�l��,$��|���8����/���!�^�W�;W���������򱨽�e��f4����s�b�:��.��Ȯa� �.;�Ě<6�=�L=w�=2ў=�y�=���=���=^y�=��=e �=���=���=��=إ�=��=�D=��<�~���8�
٭����K�/�Q�Z��}���i��寘��   �   Fe���v�M~c��;G�%��K ����Иo��|���`������:��;� H����������4�t.`�����އ������Ph��D�j����м��O� �b:��u<���<�4=(�n=`�=���=��=
��=ۇ�=I��=�w�=p��=���=uH�=�g�=�4=(M�<�ٻ���Ց��q۽��ͦ6���U���m��5|��   �   �G��c>�T�,�FQ�5���H��H
d���� Q޻<|m�< l�<��< �I<@��:��)�e���A�`_6��T�Ryf��n��k��X`���L���0�f�ح¼Xx8��9;�< 2
=�/I=	��=ᮚ=�F�=�c�=V�=���=���=�=�t�=��`=rE=t��<0ӻ�t�s�ץ��AK�o,�q�*���<�.WF��   �   ��a����<ƽ�_��g?�x�� �):\1�<�=z-#=�Q,=!=�{=��< �!<`�_���������$��L�,l�A��tB��c�����f����xd��B7��m����i��wh;�<r[=N�[=m�=���=�d�=٠=��=�=�pg=2�/=���<h�<P5!�����޻R�k8��໿�8{潾G�J}�8���   �   mýaE��ۉ��t.X�6_�H@-�xG%<�9�<l�1=�?]=��u=��z=^�m=�zP=NB&=�M�<�E]<��躸y������D�4��(ٚ��ñ���½�̽�+ͽ�rý+K������.9X�
i��c-�X(%<�+�<`�1=J:]=~�u=��z=��m=FvP=�=&=E�<6]<�H�|~�������D����ך�������½�̽f&ͽ�   �   $od�(97�pZ����i�  i;��<Xb=^�[=�o�=%��=�f�=:۠=��=�ĉ=�tg=��/=���<h�<`0!�������R�N:��ɾ��$�*J���T��O��fd�{���BƽLe���p?�T+����':h$�<�=(#=�L,=!=�v=�u�<��!< `��È����<�$��L�^l��?��=@��`��Q܊�����   �   ؞¼�X8���9;�ѓ<>9
=R6I=���={��=0I�=f�=�W�=w¿=4��=��=v�=J�`=|G=�< /ӻN�p�s�Q����Nｰ.�/�*���<��ZF�LG�g>���,�nT�����M��d������޻P�<pb�<La�<$��<P�I< C�:@�)��o���F��c6�T�b{f�Tn��k��U`�4�L�
�0�� ��   �   �d:�u<H��<��4=��n=�=��=�=���=���=���=,y�=���=9��=�I�=�h�= 4=�M�<0ٻ��ב��t۽��<�6���U���m�29|��h�N�v���c��>G��%��M �F���,�o�V����`��Z� ��:�F=��]�Ȫ�����L�4��3`�X������������\h�D����d�м�O��   �    ͚<��=6L=my�=lӞ=�{�=���=���=�z�=B��=��= ��=���=��=���=%�=��D=���<Ѓ�T�8�ۭ�t��:�/���Z��~��k�������W��d��R����x��Q�"Z'�^���6���^ui�����-��Ŏ�؋���9� �!�ƐW��Y��Ù�_������[g��k5��n�s��:�|+�� �a��/;�   �   "� =�EG=�'�=���=� �=J��=���=���=`��=��>��>b�=���=���=�H�=Cޖ=T�L=l��<�\�z#[���ɽ����XJ�!|�B6���������]5���ӯ����U���y���I���[h佖x�� �]��"�F��V���(9��l��[��g����.���ʽ�wȽV)������sǃ�P=�,�ټPٻH�R<�   �   �x!=�m=e`�=b7�=^�=V��=3�=4>v`>�B>~|>��>���=���=�
�=�y�=N�O=�á<�h����y�ɰ�X�'��4`�a���t��{����þ$Ⱦ,�þ�춾;£��)���;e�3�$ ���½(���dY���@��K���p��j��K����˽X߽4��X�⽏Gѽ���(����D���ϼ�H.��ǜ<�   �   �3=�7�=���=B�=��=��=� >*�>
>��>=�
>U�>�E�=�x�=���=�Ý=��P=��<pj���v��ښ񽨝2���n��`��Wg���þSFо&�Ծ�.о�
þ=����0���v�FB�;����ؽ2L��Β|���b� �m�>��;:����Ľ_h�M��������$�ڋ��������K�X]μ�
I� 
�<�   �   �n9=��=P��=���=�y�=�Y�=<V>"<>L�>8!>��>��>v��=��=���=�r�=ڌP=�c�<��y-��-��u6�Xs� o��G���g	Ǿ;�Ծ7پ|�Ծ{8Ǿcв�ǥ����|��=G�^<���/䦽�Q��Vyn�Zoy��[��������˽�~�����D� �M����]�ߛý�m���N�h�μ <i�|�<�   �   �3=�7�=��=��=��=��=�� >7�>&
>��>O�
>g�>�E�=�x�=��=.ĝ=��P=0�<�e��`u����r�2�:�n��_��`f��~þ5Eо�Ծ�-о�	þ@��/��{�v��B����~ؽ|J����|���b��m�y<��{8���Ľff�D�������#����!���"�K��Xμ �H��<�   �   *{!=�m=a�=�7�=��=���=p�=P>�`>�B>�|>̯>���=��=��=vz�=��O=�ʡ<�_����y���	�'�2`������y����þ�Ⱦ
�þ�궾[���(���8e��3���H�½����^Y���@�&�K���p�Wg�������˽>T߽P�罉���CѽB��5��ʼD��ϼ`.�4͜<�   �   2� =*HG=q(�=p��=J�=���=��=D��=���=��>��>��=��=���=�I�=�ߖ=��L=¬<x\�T[���ɽ����TJ��|��3��B������^2���Я����R��y���I����^b�ls����]�~
"��� ���9��l��V��)~��q)��}ʽ�rȽT$�����]Ã�D=�@�ټp�ػ��R<�   �   �Ԛ<�=hL=?z�=Ԟ=n|�=.��=���=0{�=���=�=x��=]��=r�=ʧ�=��=�D=��<�e���8��ԭ������/�\�Z��{���g�����FT������N����x�k�Q�JU'���������hi����L��(����w���$���!�ބW��S�������������ha���/����s�t�:�T����a��f/;�   �    e:h�u<��<ȗ4=>�n=��=x��=}�=L��=��=D��=�y�=���=,��=�J�=Aj�=�4=�Z�< �ػr��Б�rl۽�
���6�^�U���m��1|�>a���v��zc�)8G��
%��H �)���j�o��u�Ȅ`�����R�:��:�P/�D��������4��%`�R���ه��������g��D������м��O��   �   Ж¼XL8�@�9;hՓ<�:
=p7I=i��=ݱ�=�I�=ef�=oX�=ÿ==��=Tw�=޸`=VL=�Ȉ<��һ���s�����D��(���*��<�SF��G�z_>���,��M���� C��r d����@޻� <�y�<x�<4�< �I<���:8�)�0T���8��U6�2�S�Nnf�Zn�H�k��L`�d�L���0�t���   �   Rkd�(67��U����i�`i;��<,c=&�[=p�=���=>g�=�۠=��=�ŉ=wg=.�/=@�<0�<(!�D�����R�f2��a���=t�D�gy�A����@]���� 6ƽ�Y��4\?�L�� �+:@�<��=�3#=�W,=J!=8�=��< �!< @_�h�������$�$�K��l��:���;��J\��Cي������   �   XkýD��و���,X�^��<-��J%<�:�<�1=p@]=T�u=��z=��m=�|P=�D&=T�<�V]<@*�k��6��Z�D�����К����½̽̚ͽ�eýD>������!X��S�-�k%<I�<R�1=F]=p�u=V�z=F�m=.�P=I&=�\�<@g]<��纔e�����F�D����mҚ�����\�½Y�̽0$ͽ�   �   R���`�B��@<ƽ__��>f?���� �):�2�<��=4.#=�R,=B!=,}=�< �!<��_�4�����$���K��l��9���9��vY���Պ�e�bd�z,7��B����i�@�i;x�<Bj=b�[=�r�= ��=�i�=�ݠ=��=�ǉ=�zg=��/=��<��<�	!�l����R��3��㷿��w�NF�|�G���   �   .G�c>���,�Q����mH���	d�����L޻H<�n�<pm�<��<��I< *�:�)��^���=��Y6�� T��pf�V	n���k�pJ`���L�j�0�
��P�¼�-8��(:;��<�A
=>I=f��=���=�K�=�h�=fZ�=�Ŀ=���=T�=�x�=��`=�N=̈<��һ2�.�s�����G�+�D�*���<�lVF��   �   �d�i�v�~c�u;G��%�[K �Ê��X�o�v|�Ȝ`�`�����:��;�0D� ���$��8�4�*+`�>���ۇ�������l�g�D������мX�O��mf:��u<��<4=��n=1��=���=��=D��=���=���=0{�=���={��=L�=Lk�=p 4=H\�<��ػ��bґ��n۽����6��U���m� 5|��   �   �U�����kP����x�<�Q��W'�F�������8oi���\#���������4.���!��W�NV��M���Y��د��)c��11���s���:�4��X�a���/; ܚ<�=�L=y|�=1֞=q~�=��=���=�|�=���=B�=���=j��=o�=���=z�=�D=ĺ�<�g�V�8��֭�޺�P�/�|�Z�<}��Di�������   �   �3��?ү�|���S��ty���I�W��ze�v����]��"��������#9��l�&Y��l����+���ʽ�tȽ�%��a���5ă��=���ټ��ػX�R<�� =KG=�)�=���=��=%��=n��=~��=���=d�>h�>��=���=`��=_J�=��=z�L=¬<X\��[��ɽ���VJ�a|��4������k����   �   Ⱦ�þ�붾X���)��r:e�T3�#�<�½����aY���@��K�f�p��h��B��~�˽�U߽����?EѽI�������D�|�ϼ�	.�,Ϝ<�|!=4m=�a�=�8�=��=���=J�=�>�`>BC>�|>�>r��=���=��=�z�=D�O=�ʡ<�`����y���ɕ'�3`�f���f���y����þ�   �   ��Ծ/.о]
þ��^0��`�v��B�����ؽnK��L�|�N�b�D�m�%=��.9����Ľ<g�"���������#ུ���������K��Yμ��H���<��3=Y8�=���=��=���=���=(� >j�>R
>�>t�
>��>F�=y�=T��=aĝ=F�P=x�<�e���u��J��Ɯ2���n��_���f���þ�Eо�   �   �E�Dy�DQh�}�N��80��P��彳϶�Ł��=��o���϶�.��7P�80��N��Ph��Cy��E��By���g��,L��e)�PM������!I�0�X��#�<f2@=��=Z�=�q�=@��=�>�H	>�>�<>�>�H	>-�>���=Lr�=��=>��=*4@=(�<��X�I�T����L�e)�2,L�V�g�NBy��   �   ��y���s���b�ǨI��~+����O޽����Q$���ه��#��F����N޽d�?~+�L�I���b�~�s���y�%�s���b�[�G�c�%��Z��,����E���R�$��<J�==*�=�¶=��=PS�=��>�>��>�>��>�>��>�S�= �='ö=��=�==X��<(�R�E�����hY����%���G�T�b���s��   �   Bi�K�b�&�R�͠:����4����SȽ����7���k�"7�8���RȽ1���{��[�:�θR��b�@i�-$d��yT���;�����r������9��E�x��<��5=�/�=���=H��=���=R��=�w>�V>,�	>�V>x>���=2��=���=<��=�0�=t�5=p��<(�E�0�9������q�c��,�;�ZyT��#d��   �   q�O��[I���9��<#�d��ٽ.䥽��y���D��2�f�D���y�d㥽ٽ�c�_<#���9��[I�l�O�GL�ػ>��)�?
��eڽ����Z�+��6=� ΃<
]&=��}=��=>��=���=C��=p�=�@>ڒ>A>��=���=B��=���=���=��}=�^&=�у<�.=�$�+�~����dڽ�	��)���>�L��   �   �:0��[)���������ڽ(��B�s�@�)�����|�Ӽ����<�)���s�='����ڽN��Z��X[)��:0�fa.�v$�u�5�������S���U��K� �E<6N=2]=ҿ�=<ޯ=���=\�=n�=9��=0��=P��=4n�=V\�=��=�ޯ=Y��=p]=�O=��E<��K��S��R�����L����t�3$�Ga.��   �   f��v��ۘ�L]ɽ�z���ya�����^��x���.������\�����xa�z���\ɽP��K��Z��}	�`r��j���[ҽ�ب���w����
��p��;з�<�-=�ep=ȕ=�=�k�=�^�=�|�=?��=�|�=(_�=�k�=`�=xȕ=�fp=8�-=T��<ྜྷ;�����w��ר�J[ҽ�i��.r�j	��   �   ��ս�.Ľn���yb���^<�tvۼh����;�X<LK�<P�X<p��;0���sۼp]<��a��狨�@.Ľ��ս�ܽ�h׽��Ƚ[[�������k�T�'�|�ü`�ܻ &<�D�<�,=��g=�$�=t�=�.�=I�=ǵ�=.I�=(/�=��=E%�=T�g=��,=G�<�&<��ܻ~ü�'�h�k����Z��B�Ƚ�h׽�ܽ�   �   �5������T�I�������� �t:��<L��<=h�=Z=���<��< �t:\������^�I������5���ޡ�>y��ĩ������0��0ks�P�G�N����� �P{�;(׭<j�=��K=n�{=B�=ׅ�=jp�==p�=�{=J�K=6�=�ح<���;X�����M�l�G�Jjs�E0����������+y���ޡ��   �   z:�n?	�@P��pL���j@<�O�<n#=�;M=p�g=:�p=��g=V<M=�n#=�Q�<�n@<`D��tN���>	��y:���a�X�~��ӈ�_u���u��#Ո���~���a���:��F	��^�������O@<�B�<.h#=06M=�g=��p=V�g=�6M=�h#=hD�<�R@<`~���\���E	��:���a�d�~��Ԉ��u��Bu���ӈ�v�~���a��   �   $��� �����;L�<J�=4�K=��{=��=<��=�r�=X��=��=Z�{=�K=4�= �<���;�������4I��G�fis��0���������|���⡽�9�������I����������r:@ӂ<H��<N=��=�=D��<�Ԃ< s:���������I�����t9��N⡽�{����������0���is�X�G��I��   �   ��ܻ&<�N�< �,=h�g=D'�=��=1�=(K�=ҷ�=BK�=O1�= �=�'�=:�g=ڡ,=hP�<�&<��ܻ0yü��'���k�"���\���Ƚ?l׽� ܽJ�ս3ĽҐ���f���f<���ۼ��� S�;@hX<�?�<hiX<pW�;����ۼ�e<�:f��m����2Ľ�ս� ܽGl׽-�Ƚ	]��j����k���'��zü�   �   �ȝ;d��<ʞ-=tip=�ɕ=��=�m�=�`�=H~�=��=X~�=�`�=�m�=F�=dʕ=Njp=��-=8��<`Н;���(����w�|٨��]ҽm��t���������T�ｈaɽ�~����a�H���j��X
��[����`i��d���a�6~��aɽ�｛�������&t�dm��^ҽ�٨���w�������   �   �E<�P=�]=E��=�߯='��=�]�=do�=���=���=���=�o�=�]�=r��=�=���=�	]=�Q=p�E<��K��T��S��p��ً��Tv�$�Rc.��<0��])�Ė����-�ڽY+��,�s���)������Ӽ$��� �)�.�s��*����ڽf������])��<0�^c.�6$��v�`���	��XT��V���K��   �   Ѓ<�^&=��}=��=N��=���=N��=m��=vA>S�>{A>���=���=@��=���=���=~�}=�_&=�҃<�/=�`�+�����cfڽ�
��)�)�>��L�H�O��]I���9�r>#��e��ٽ�楽\�y�FE�V�2��E���y�楽ٽIe�(>#�o�9�e]I�E�O��L�]�>�8)�:� gڽt���܋+��5=��   �   ���<��5=z0�=\��=���=���= ��=Hx>�V>��	>�V>Zx>2��=���=X��=���=�0�=��5=x��<X�E�l�9������r�L��D�;��zT�R%d��i���b�l�R���:�������UȽt���:�Ȑk�V:�����TȽl��������:�0�R���b��i�o%d��zT���;�����s�����9���E��   �   ��<��==��=�¶=�=�S�=Ø>>��>>��>&>ߘ>�S�=f�=^ö=�= �==�<0�R��E�s���MZ��M�%�s�G��b���s�b�y�h�s���b�`�I�O+�d�sP޽����%��Nڇ��$��C����O޽��~+��I�Z�b�B�s�e�y���s�H�b���G���%�5[��d����E���R��   �   �$�<�2@=���=t�=�q�=N��=�>�H	>�>�<>�>�H	>(�>���=Kr�=��=&��=�3@=l'�<�X�hI������L�:e)�K,L�j�g�ZBy��E�Dy�6Qh�l�N��80��P���形϶�����G������/϶�[��TP�-80��N��Ph��Cy��E��By���g��,L��e)�2M����2!I���X��   �   h��<4�==��=Hö=J�=�S�=٘>">��>>��>2>�>)T�=��=�ö=��=h�==8��<��R�DE�����OX��&�%�&�G���b�)�s�ڍy��s�'�b��I�~+�J�zN޽����u#���؇�:#��|����M޽���}+���I���b���s�܍y�K�s�۳b���G���%�7Y������E��R��   �    ��<6�5=g1�=��=}��=���=L��=fx>W>��	>W>xx>���=4��=ڲ�=x��=�1�=h�5=ԋ�<�E�H�9�����9o���ɢ;��wT�u"d��i���b���R�h�:��������QȽ���4���k�4����*QȽ5���\���:�g�R���b��i��"d�xT��;�|��	p�s�����9� �E��   �   �؃<�a&=�}=��=��=���=���=ŀ�=�A>z�>�A>��=���=���=^��=���=�}=c&=�ۃ<0=�F�+�M���)aڽ���)�l�>��L�>�O��YI���9��:#�Xb��ٽ_᥽��y�h�D���2���D��y��ॽ)ٽb��:#���9�fYI�9�O�L���>��)�.��aڽ�����+��=��   �   @�E<�T=�]=p=��=���=^�=�o�=���=ۭ�=���=�o�=>^�=��=��=�=�]=�U=��E<��K�PL�{N��0������=r��$��^.�80��X)�3��i��_�ڽY$����s�F�)�l�����Ӽ������)���s��#��Ɉڽ$������X)��70��^.��$�vr�%������O���M�p�K��   �   @��;X��<6�-=�kp=�ʕ=��=n�=/a�=�~�=M��=�~�=Za�=Zn�=��=R˕=�lp=�-=@��<0��;�������H�w��Ҩ��UҽHd��Do�s�x�����s��KXɽCv��Rqa�t��xQ��������p��P�����Bpa��u���Wɽ��u��e��u�Vo��d��8Vҽ,Ө�H�w���������   �   P�ܻ0+&<�U�<��,=Z�g=(�=G�=�1�=�K�=3��=�K�=�1�=��=Z(�=$�g=r�,=XW�<�.&<��ܻ jü��'�t�k�U	���T��,�Ƚ�b׽�ܽػս�(Ľۆ��V]��nU<��eۼ0�� ��;@�X<�W�<��X<���;����cۼlT<��\��n���_(Ľ��սrܽ�b׽N�Ƚ!U���	���k�R�'��kü�   �   Ԩ��x��@��;H�<&�=��K=ȣ{=-�=���=(s�=���=f�=h�{=d�K=�=�<��;X��|���
B��G�|^s�=*���}��X����r���ء��/��5�����I����t�����v:��<��<b=��=�=��<T��< �v:���������I�Ձ��}/���ء��r��N����}��M*���^s�`�G��B��   �   �t:�x;	�4J��`:���q@<4R�< o#=�<M=0�g=��p=t�g=(=M=�o#=T�<xu@<�2��tH���:	�vt:��a�2�~��Έ�~o��o��͈�N�~��a��n:��4	��;��@�� �@<_�< u#=0BM=|�g="�p=��g=�BM=�u#=�`�<x�@< ����9���3	��m:�T�a���~�C͈��n��\o���Έ�L�~�^�a��   �   �3��C�����I����ȧ����t:��<���<�=�==��<��< u:�������ʍI�셀�g3��ܡ��u��w����~���*���]s��G��>���������;@��< �=2�K=�{=��=���=|u�=��=��=��{=��K=��=��<@��;@��(����=��G��\s�Z*���~��A����u��'ܡ��   �   �ս0-ĽZ����a���]<��tۼp�� ��;��X<dL�<p�X<P��;H��rۼH\<�a��ڊ���,Ľ��սvܽf׽�ȽW���
����k�>�'��fü��ܻ<&<�^�<b�,="�g=Q*�=|�=�3�=�M�=2��=�M�=�3�=��=�*�=��g=\�,=�`�<�@&<�ܻXdü�'�T�k�
���V����Ƚ�e׽bܽ�   �   ������
�ｬ\ɽ^z���xa�:���]������*������[�����Twa��y���[ɽ|�ｾ�������8q��g���Xҽ�Ԩ�ֵw����������;0��<��-=�op=�̕=��=�o�=�b�=S��=��=j��=c�="p�=��==͕=�pp=¦-=���<0�;p�V��0�w��Ө��Wҽg��q�~��   �   $:0�[)�Z��y��:�ڽ�'����s���)�̦����Ӽ̥����)�d�s��&��]�ڽ�����Z)�:0��`.��$�	t������	��9P��~N���K���E<~V=X]=�Ñ=��=1��=^_�="q�=6��= ��=M��=Lq�=�_�=���=e�=Lđ=�]=�W=x�E<0�K��L�7O����������s�V$��`.��   �   �O�k[I���9��<#��c��ٽ�㥽��y���D���2��D�p�y�7㥽�ٽ�c�6<#�]�9�<[I��O��L�<�>�3)�X	��cڽ=����+� =��ك<�b&=��}=���=���=z��=���=���=B>�>B>��=���=���=l��=���=�}=�d&=�݃<�=�Ѓ+�����bڽ���)��>��L��   �   i� �b��R���:��������SȽ����7���k��6� ���RȽ���g��?�:���R���b�i��#d�RyT�1�;�d��|q�y���4�9�X�E���<��5=�1�=���=��=���=��=�x>PW>�	>\W>�x>)��=���=���=!��=�2�=^�5=��<��E���9�,���0p������;��xT��#d��   �   ��y���s���b���I��~+����O޽����J$��vه��#��5����N޽\�6~+�B�I���b�l�s���y��s���b��G��%�Z��i����E�P�R�䫙<4�==�=vö=��=*T�=��>F>��>6>�>]>�>�T�=�=Ķ=��=��==��<��R�ZE�����X��z�%���G�&�b���s��   �   @� �%����"�˽���/\���oy�,yn��Q���㦽� ླྀ;�*=G�$�|�b���в�:8ǾX�Ծ7پ[�Ծ�	Ǿ����ho��8�s��u6��.���.��0��`_�<�P=;r�=B��=���=.��=x�>��>4!>R�>4<>TV>Z�= z�=^��=ĺ�=���=p9=�~�< �g�t�μ��N�Nm��I�ý]�����   �   ?������g�w�Ľ�9���=��ֲm�P�b���|��J���~ؽ
���B�x�v��/��k�
þ
.о��Ծ�EоIþ8g���`���n�	�2�����w��`n����<�P=�=��=�w�=E�=�>�
>��>�~
>
�>Ħ >���=���=%�=���=�7�=b�3=��< �H�lZμ�K����������#�����   �   ��罤V߽O�˽���i����p���K���@��`Y����9�½x��3��9e��(�������붾��þȾ��þVz��������j4`�>�'���὎�y��k��x��<��O=�x�=�	�=���=���=P�>(|>�B>$`>�>��=���=� �=�6�=�_�=�m=vx!=�ǜ<�?.�<�ϼ
�D����!���Eѽ����   �   �ʽ�,��u���Z��ll�<%9����0��@"�|�]�,u��Ld佧����I��y��S��G��-ү��3������𦥾c5���|��WJ�^��x�ɽ�#[�("\�P��<j�L=9ݖ=�G�=��=���=j�=P�>D�>c��=��=���=��=���=���=_&�=�CG=�� =8�R<�ٻ�ټ�=�Fƃ� ���~'���uȽ�   �   �������W��6�W���!�1�䂢�L����"��.���mi�������� W'���Q�$�x�DP�����V�� ����i���}���Z��/�ļ�~ڭ�j�8�����<b�D=��=R��=J�=n��=���=T �=��=zy�=��=2��=5z�=�ў=�w�=�L=>�=ǚ<��.;�a�D,��0�:���s��3���e��ױ���   �   Ћ�/`�n�4����0����J� <����: ��H�`�R{���o�щ���J �l%�;G��}c��v�9e��5|���m�s�U�f�6���s۽�֑�6�0ٻ�I�<p4=�f�=�G�=���=3��=�w�=A��=��=5��=4�=�=��=��n=4=���<`�u< �b:�O���м����D�� h��������އ��   �   �_6�nB��f�� �)� ��:��I<4�<l�<hn�<�	<0F޻0��Nd��G��%���P���,�Gc>��G�HWF�̃<���*��,�JL�⦴���s����=ӻh��<*D=��`=t�=��=H��=���=V�=d�=G�=$��=d��=�0I= 3
=Lē<�9;�t8�@�¼�� �0��L�,X`���k��n�Lyf��T��   �   ��|���@�_�г!<�~�<,{=�
!=�Q,=�-#=��=�3�< *:��<e?��^��<ƽ|���`����D��r}�H��{潪���;9��l�R������:!�p�<���<@�/=�og=Q=��=٠=�d�=ڄ�=Hm�=��[=F\=��<��h;��i��k��B7��wd�*����ߊ��b��dB��A��Rl�L�h�$��   �   <{����躐B]<0L�<�A&=VzP=�m=��z=Ғu=X@]=V�1=�;�<�L%<X:-��]�-X�O���E���lýe&ͽB�̽	�½"����ך�����D��������@k�82]<\C�<=&=�uP=Z�m=��z=��u=�:]=�1=x-�<@,%<X_-��g� 8X�����J��rý�+ͽئ̽��½�ñ�]ٚ������D�X���   �   84!���<,��<��/=�sg=Tĉ=��=0۠=�f�=c��=p�=J�[=rc=��<`i;0�i��X��l87��nd�����U܊� `��v@��@��l�jL��$����dň��#`���!<Pt�<v=�!=�L,=T(#=��=�%�< #(:�(��vo?��d��IBƽ���7d�8��P��,��MJ�y�5����:����R������   �   `8ӻ���<�F=l�`=�u�=n�=��=k¿=
X�=0f�=yI�=ر�=k��=R7I=@:
=�ӓ<��9;�U8���¼8 ���0��L��U`�&�k��n��{f��T�Rd6��G�Pq���)�@/�:8�I<���<Da�<�b�<��<�~޻t�뼰d�M��,��T�u�,��f>�;G��ZF�φ<�h�*��.�fO�������s����   �    ٻlK�<4=h�=4I�=���=���=y�=���=���=2��=h�=a��=i�=��n=ږ4=��<��u< @d:��O�t�м8���D�6h�����������Ȑ�Z4`���4�X������_��X=����: V�в`�@��Ğo�w����M �r%�s>G�n�c�#�v��h�H9|���m�(�U���6�8��u۽gؑ����   �   @��ȫ�<f�D=��=>��=P�=���=���=��=Z��=	{�=���=��=D|�=�Ӟ=�y�=
L=~ =�Κ< (/;0�a� *��T�:���s�?5��Og���������bÙ�BZ��j�W���!��:�h���Ŏ� -��̮�$ti�k���p����Y'�|�Q�H�x��Q��M���W������:k��*��$�Z���/����ܭ�,�8��   �   �$\�`��<
�L=�ݖ=dH�=���=a��=H�=��>��>���=0��=��=���=�=��=�'�=�FG=�� =��R<P�ػP�ټ�=�ǃ�h���,)���wȽ�ʽ/������I\��� l�F)9����>��|"�:�]��w��yg佁���I�*y��T������ӯ�[5�����3���~6���!|�YJ�l����ɽ�%[��   �   �l��t��<��O=�x�=f
�=J��=^��=��>z|>�B>�`>J>d�=���=��=�7�=�`�=�m=�y!=�ɜ<�8.���ϼ��D����/��VGѽ@��=��PX߽��˽���k��x�p�t�K���@�dY����;�½���3�8;e��)�������춾�þ#Ⱦ��þA{���������p5`��'�����y��   �   �n��,�<B�P=Ý=J��=@x�=hE�=D�>9�
>��>&
>?�>�� >.��=1��=��=(��=�7�=�3=(�< �H�[μ��K�/���h����$������z��h�L�Ľ�:��g>��V�m���b�N�|��K���ؽ����B�e�v�r0���󮾭
þ�.о&�ԾpFо�þ�g���`��a�n�]�2�%��x���   �   0��4`�<j�P=`r�=^��=���=A��=y�>��>7!>U�>4<>SV> Z�=z�=R��=���=u��=�o9=8~�< h��μ��N�qm��k�ý.]�(���D� �!�����˽����(\���oy�Hyn��Q���㦽-��;�S=G�V�|�z���"в�G8Ǿ`�Ծ7پW�Ծ�	Ǿ����Uo���s��u6�V.���.���   �   �i����<��P=�Ý=���=�x�=�E�=W�>G�
>��>0
>N�>� >T��=e��=��=���=q8�=�3=�<�MH��Vμ�K����������"������u��f�i�Ľ�8���<��<�m���b��|��I���}ؽ���]B�ڷv��/���򮾛	þ�-о�ԾREо�þ�f��`���n�&�2�1��v���   �   �c��Xǡ<��O=�y�=�=���=���=��>�|>�B>�`>e>��=ܪ�=�=<8�=sa�=^m=|!=,Ϝ<@ .��ϼԻD��������Cѽu��[��pT߽8�˽���g��2�p���K���@�^Y�c����½��j3�D8e��'������궾�þ�Ⱦ��þ>y���������2`���'�L����y��   �   �\��<��L=ߖ=WI�=`��=��=��=��>��>η�=x��=X��=���=��=Ұ�=�(�=�HG=� =X�R<`�ػ��ټ|=�Ã�ր��3$���rȽ�ʽ�)��}~��TW��Tl�� 9�J����
"��]��r��~a�����I��y�FR������Я�\2��!���k����3��|�=UJ�<����ɽZ[��   �    l�L��<��D=C�=i��=)�=,��=]��= �=���=\{�=$��=~��=�|�=jԞ=�z�=2L=X=֚<�r/;�a�����:�D�s��/��^a������������T����W���!��%�Hx��$����������gi�<�������T'��Q��x��N�����CT��$����g��&|����Z�*�/�.���խ�f�8��   �   0�ػX�<�4=�i�=�J�=潼=U��=�y�=O��=��=���=��=҉�=��=�n=��4=���<p�u< Be:P�O���м����D���g����(��ڇ�̂�h&`�d�4�R������h1���:�@Q�:�����`��t� �o�Y���DH �w
%��7G�>zc���v�2a��1|���m���U�ݣ6�J�Lm۽�ё����   �   0�һ�ƈ<^K=�`=�v�=h�=Ɣ�=�¿=�X�=�f�=�I�=<��=׭�=\8I=�;
=Hד< �9;pI8���¼��j�0�R�L��L`���k��n��nf���S�V6�X9��U���)����:�I<��< x�<pz�<0#<�޻,���c�aB����jM�=�,�L_>��G�!SF��<���*�4)�yEｯ���8�s����   �   �!���<��<d�/=lvg=Aŉ=o�=�۠=Wg�=���=yp�=�[=@d=�<`(i;X�i��S��p57��jd����Hي�m\��<���:���l���K���$�`��0����N_���!<���<��=�!=�W,=�3#=��=�A�< ,:���Z?�Y���5ƽH��]����<��vy�*D��t�ĵ���2����R�����   �   �l�� C��S]<�R�<�C&=|P=V�m=x�z=��u=A]=��1=8=�< P%<�6-��\��+X�P����C��(ký5$ͽ��̽��½+����Қ����t�D�����g��@��Hc]<[�<hH&=��P=�m=2�z=��u=dF]=��1=�J�<�n%<�-��R�� X������=��veý�ͽ̽��½����К�X����D�����   �   0������_���!<���<�|=�!=�R,=�.#=F�=�4�< @*:���zd?�^��y;ƽ���X`�?��T��G|��F�zx潫����4����R�p���X!�h�<h
�<��/=zg=4ǉ=q�=�ݠ=�i�='��=!s�=�[=k=D�<��i;�i��@���+7�pad��zՊ�XY���9���9���l���K�"�$��   �   `Z6�>>�``���)� �:��I<�<�m�<�o�<�<PB޻�뼸d�[G�����P���,��b>�G��VF�ق<���*�{+��H�(���<�s��p�һ�Ȉ<\M=��`=rx�=��=q��=�Ŀ=dZ�=�h�=L�=̴�=���=�>I=�B
=x�< 7:;*8���¼N����0��L��I`�T�k�$	n��pf�� T��   �   ����+`��4���������F���;�@��:`��x�`��z�N�o������J �D%��:G��}c�-�v��d�H5|��m���U�H�6�:�&p۽�ӑ�"�p�ػ�X�<�4=�j�=�K�=!��=���={�=���=ċ�=m��=��=,��=���=��n=��4=���<��u< �f:X�O���м���8D���g�m������ۇ��   �   q�������V����W���!��/似���p���"��Ҩ�nmi���������W'���Q��x�0P��w���U��ʯ��{i���}��2�Z��/���� ح��8�Xq����<<�D=��='��=�=#��=y��=2�=��=�|�=���=S��=�~�=�֞=�|�=�L=�=Hޚ< �/;Pa����p�:��s��0���b�������   �   �ʽ�+��̀���Y���l��$9�2�����"�>�]�u��-d佔����I��y�~S��9��ү��3����������'5��3|��VJ������ɽ�[��\����<��L=Wߖ=�I�=���=���=t�=^�>e�>ڸ�=���=���=v��=2�=m��=w*�=$LG=�� =��R< �ػ��ټ�=��Ã�ׁ���%��otȽ�   �   ��V߽��˽���Ii��0�p�L�K���@��`Y����#�½n��3��9e��(�������붾�þȾ��þ;z�����ڑ���3`�'����y��f���š<J�O=�y�=Q�=��=$��=��>�|>@C>�`>�>��=ѫ�=�=N9�=b�=`m=�}!= Ҝ< �-��ϼ��D�2������Dѽ����   �   ���W��g�X�Ľ�9���=����m�,�b�t�|��J���~ؽ���B�o�v��/��h�
þ.о��Ծ�Eо<þ(g��y`����n�˝2�,��Gw���k��|�<@�P=�Ý=���=�x�=�E�=r�>f�
>�>Z
>|�>B� >ʷ�=��=o�=
��=�8�=
�3=��<�'H��Uμ�K�Ъ�����V#འ����   �   ��+�@%��K�*^ �<�<���0�P�����~�񽡛/�Ss�2���?�ʾ6p��F#�<G�X&�Ky)�,&��8����O���Ǿ�1��a�����"���� ��<~|k=p��=F��=���=�F>pU>��	>]>��>?>�=��=���=*��=g�=ӂ�=�s=�e9=��<�v< �8��a�.Ҽ#��$��   �   �'%��&�������8�Ѽ�BԼ���&�E������꽠�*�~mm��"��\kƾ�wﾄX
�6?�Z�"��@&���"��?��*
�pC��þv���6\���t?��,���P��<D�l=Tz�=P'�=���=;n>);>q>j�>Q�>���=]��=��=2��=��=G��=~�h=�q/=�t�<�]<��g���g�t3м��
�����   �   �-����lp�,i��dޜ��w����мlH%�Ų���cӽ<��#R\����k���_��?� t�x�����Q�����\�m��uO��M䎾�7N����YD���4���Y�<�yp=F��=
��=:��=���=.�>GE>X�>�>�=b�=v��=F^�=���=�=�>{=V�F=ƣ=���<8�<���p�}���̼DX�N;��   �   ��,�ʼ�=���Y��R�@e��j����lIR�K믽T8�e�A��x�����\�ʾF뾑��	K��Y�8��G�����˾���M؀���8���Jep�0���<҃t=TW�=�[�=`��=�Z�=i�=�U�=�N�=�0�=���=L��=/��=(u�=��n=(�<=|�
=4i�<-< �����%�lQ��,�ͼЪ�:���   �   ����x��O�@�`�d;P5�; ���xD��������"׽���Z�[�b���1��[]˾]��E;�^����P���rξ:���ϐ���^��e��ƽ��=�@�^���=:�v=p��=� �=E�=���="�=���=V��=�k�=޴�=��=^m~=��G=K=Ty�<p�E<�;�:P���Sk�����P2ʼTT޼@���м�   �   xjg�Ѱ���i;��>< 9�<�,�<���<p��;?@�����J��X��BR-�Se��E��J���t��xɾ��ξ�:˾�U��;O������Yq�R�8�P������
�@�q;R8=�,t=0)�=��=�u�=��=�z�=x��=���=9\�=2��=�JO=��=���< �; d�������ּFF������TE���44�,����   �   x���%N;��n<�F�<��=�=��=�(�<8�-<�?C��,��x��1�����+���Z������ړ�z���`p��u%������Bꉾ��l���@�����̽��p� �����<2�=\�j=M��=B�=[�=�U�=���=8��=�=�2e=��=t��< 4�8�u���M��[F��(n������Y��3���4_q���S�p.���D����   �   p�ڻ��<ty�<P�=�l8=��L=ԁM=��6=��=x�n<0�&�b�&��L���9�*q��=��oZ��ln� �w���u���h�}�R��v5�k�����S��F�/�~\�0*M<�=�W=5Ǉ=`U�=r�=Y��=Kҕ=j�=�8A=\��< ��;<c����.�S݅����:�˽!�޽�X�;��Cн]���ݙ��o���(��"¼�   �   0-�ДN<�L�<h�:=$Vh=�V�=ҹ�=�\�=�*]=��"=Xd�< <���R�����	���<��%��8%��l.��/�
�'����$��=Zٽ�楽&�c��Q���*�P�N<�I�<�:=,Sh=�T�=η�=9Z�=H%]=l|"=�T�<�����]�"������D��g�"=%�@q.�&/�܄'�I�����^ٽ!꥽8�c�@V���   �    �\�`)M<��=βW=iȇ=�V�=4�=n��=�ԕ=F�=�?A=̕�< ��;�L���.�}օ�ş����˽̽޽�Q��ཇ>н���qڙ�d�o���(�� ¼ �ڻ �<�t�<n~=~i8=��L=d}M=\�6=��=�n<8�&���&��R��A�<u���=��tZ��qn��w�f�u�+�h�Z�R��y5���ʢཀྵV����/��   �   ����8�<t�=t�j=6��=x�=��=~W�=���=���=��=z9e=��=���< �8X_��B��OF��n�P����T������vXq�ΚS�m.����P������N;��n<�?�<�=ܝ=0�=P�<`�-<]C���,��}��������+�لZ����0ݓ�'���s��(��[���^쉾s�l���@����̽�p��   �   �
���q;8=.-t=�)�=��=�v�=	�=�|�=���=h��=_�=p��=ZRO=��=\Ӟ<N�;`������ �ּ�>����B����3�Т���qg� 尻�ei; �><d1�<\$�<pz�<�_�;�W@�>���N�����yU-�e��G����������{ɾ��ξ[=˾X��`Q���	���\q���8����d����   �   �>�@_� �=��v=ὧ=��=�E�=Ρ�=z#�=��=6��=n�=h��=��=�s~=F�G=R=8��<�E<���:�ỠBk�x����.ʼ S޼0Ἠ�м����x�\��[���{d;p�; �!��D�Z��k����&׽%��]�[�,���3���_˾����=�����S����wξ�;��ѐ���^�yg�0�ƽ�   �   �gp��0� �<�t=�W�=p\�=
��=n[�=b�=�V�=P�=T2�=���=^��=tè=�w�=z�n= �<=�
=|q�<(-< A����%��O��0�ͼ���=�����ʼ@C��Y��^��r�0�j�$��2NR�*:���A��y�������ʾH뾚��L��Z�@���G�8���˾3���9ـ�H�8�����   �   0E��X6��Y�<�yp=w��=d��=���=��=��>�E>̫>�?�=� �=Ҡ�=�_�=<��=��=�A{=&�F=H�=���<x�< ��0�}���̼(Y��<�(/�����t�|m���✼�|��  ѼzK%������eӽ����S\�����������y@��t�@����������3]�t��IP���䎾u8N�D���   �   �?������\��<t�l=�z�=�'�=��=\n>T;>6q>��>��>���=��=��=���=� �=���=��h=s/=�v�<�]<��g��g�04мF�
�n���(%��'�������Ѽ$EԼ0���E�����)�l�*�rnm�.#��lƾ�x��X
��?���"��@&���"�G@��*
��C�J�þ���*7\�`���   �   w"�� �����<�|k=���=e��=��=�F>rU>��	>]>Ā>H>�= ��=���=&��=b�=Ƃ�=��s=�e9=��< v< ��8`�a��.ҼH#�(�$���+�J%��K�4^ �`�x�����P��������ӛ/�VSs�S���c�ʾTp��T#�FG�_&�Ly)�*&��8�u��1���Ǿ�1���a�����   �   >���������<��l=�z�=�'�=/��=un>f;>Eq>��>��>���="��=��=$��=� �=K��=��h=t/= y�<�]< Pg�ȅg��/м��
�����%%�:%������l�Ѽ�?Լz����E�����&�2�*��lm�E"���jƾBw�6X
��>���"�(@&�0�"��?�C*
��B�<�þ����5\�J���   �   B���,��`�<b|p=^��=
��=$��=^��=��>�E>�>"@�=� �=��=`�=���=�=�B{=��F=0�=l��<؟<������}�̼̐^T��7��)�r�� j�Lc���؜�xr����м�E%�Z����aӽ7���P\�<������H� ?�ms����5�����N���[���HN��L㎾�5N�3���   �   �^p� �/�Ȉ�<��t=�X�=`]�=���=�[�=��=�V�=OP�=�2�=���=���=�è=x�=��n=��<=.�
=�v�<0-< H����%��D���ͼP��/��t�켔�ʼ�4����X�C��V�(�j�d��*ER��诽�6���A��w������ΗʾWD뾕���I�|X�"���E����A�˾o����ր���8�9���   �   �=� �^� =Чv=l��=��=�F�=a��=�#�=r��=���=Tn�=���=5�=�t~=n�G=�S=��<�E<�b�:����/k�8����!ʼtD޼`���м���x�w��9�@K���e;pZ�;  ��x�C�j������׽g����[�����/��:[˾���8�����N�-��ξ�7���͐���^�c�U�ƽ�   �   B
� Yr;�>=�1t=�+�=��=�w�=�	�=}�=ޤ�=���=`_�=Ό�="SO=��=�՞<�Z�;���t���<�ּ�:�������;����`"弈����Kg����� �i;��>< D�<(7�<���<���;`'@���{F��h��FO-��e��C�������0vɾ*�ξ�7˾�R���L������Uq���8�>��铞��   �   H����<�=V�j=���=��=��="X�=.��=��=U�=*:e=J�=���< ̟8�\��n@��MF�Jn������R��f���TRq���S�e.�������������N;`�n<S�<��=��=H�=<4�<�-< #C��x,��s������+�Z|Z�Q���ؓ������m���"��@����牾,�l�t�@�����̽��p��   �   HW\��KM<^�=��W= ʇ=X�=�=��=:Օ=��=R@A=��<@�;�K��8�.��Յ������˽��޽&P���<н��י���o���(��¼@>ڻ��<���<ć=�r8=<�L=V�M=0�6=ڴ= �n<��&�v�&��F���2�,m���=��jZ�zgn���w�>�u���h���R�r5�L����ཏM���/��   �   �8�N<�X�<:=>Yh=�W�=���=']�=�+]=��"=�e�<`7��PR�]��2	��<����T8%�Yl.�G/�'�'����֏�4Wٽ�㥽��c��A����дN<[�<��:=�[h=TY�=x��=N_�=�0]=��"=t�<���G�P��H��^4������3%��g.�/�<|'�`����vRٽ�ߥ���c��;���   �   =ڻ��<ȃ�<"�=�o8=��L=>�M=~�6=l�=�n<��&���&�NL���9�q�ϒ=�soZ�]ln���w��u��h���R��u5� ���཮P��,�/�0`\��HM<��=ָW=ˇ=eY�=��=�=wו=f�=�FA=`��<�I�;�6��B�.�Pυ����˽9�޽I�k�߽_6н>��Sә�r�o�@�(��¼�   �   ��@�N;P�n<�L�<�=��=�=�*�<��-<h=C���,�`x��������+�e�Z������ړ�Z���6p��?%�������鉾��l���@�b��-̽�p�p���� <��=��j=���=��=�=�Y�=�=f��=�=�@e=��=0��< ��8G���4��AF�tn�����M��𔂽Kq�>�S�^a.����Ĕ���   �   �Qg�������i; �><�<�<P/�<|��< ��;�<@����`J��*��*R-�<e��E��<���a��xɾؽξ�:˾oU���N�����'Yq�\�8�6�������
� 7r;�==
2t=�+�=v�=�x�=�
�=�~�=Ŧ�=���=b�=珆=BZO=��= �< ��;н��唼خּ�2��}����R7����� �d����   �   `���x�E�@�����d;`=�;  ���D�J�������"׽���J�[�Z���1��R]˾T��8;�I����P���Aξ�9��hϐ��^�e�&�ƽ��=���^���=~�v=���=,�=vG�=Z��=%�=���=F��=bp�=��=��=�z~=��G=rZ=��<X�E<  ;0q��k�����ʼ0B޼P���м�   �   @���ʼ:����X��N�`b�إj�D��IR�/믽E8�W�A��x�����Y�ʾF뾎��K��Y�/���F�f���˾ѻ��؀�[�8�̓콊bp�x0���<�t=�X�=�]�=*��=�\�=��= X�=�Q�=4�=���=���=ƨ=gz�=��n=��<=�
=��<�--< �����%�B��,�ͼ��T1���   �   R+�:�� n�tg��ݜ��v����м0H%�����ncӽ1��R\�����g���[᾿?�t�t�����J��
���\�T��VO��)䎾,7N�6��|C���0���]�<�{p=P��=&��=b��=Ĝ�=��>F>O�>A�=�!�=P��=na�=��=��=�E{=ƻF=�=`��<�<�탻X}�x�̼�T��8��   �   �&%� &������ѼBԼ����E������꽞�*�xmm��"��Ykƾ�wﾃX
�8?�Y�"��@&���"��?��*
�dC�۲þe���6\����?��\���<��<@�l=�z�=�'�=@��=�n>�;>kq>�>ۋ>>��=���=`�=��=�!�=��=�h=~u/=�{�<]<  g���g�X/м �
�F���   �   �yU<��Z<pY<��5<�Ɯ;P��Tn���h��T��k�7�稆��͹�pm�����5���P�2�e��Qs��x��Rs���e��PP��K5�z��:��>���l�z��������ƈ�d+�<���=:��=p��=t��=��>2c>��>��=���=/=�=���=��=ꧨ=,j�=څ�=b<`=B�<=1=�D�<\k�<�W�<|z<h*\<�   �   ��[<�~g<�^k<�L<�+�;P�ɻ�3弬�|�mF�l�2�-���ʵ�Ww�"��m2�ЮL��a���n�D�s�\�n�3�a���L�e�1��!�������hu�������u�T=l�=$��=���=�4�=�c>��>ɘ >ʊ�= ��=���=5�=4ڳ=�3�=�Ҍ=�'t=�=P=H2.=ĥ=<��<��<�#�<x�o<�Z<�   �   ��j<$(�<(O�<t�<h�7<��\5��xZ��#˽��$�V�t��(���ྊ�\g(��nA�PU�,!b�j�f�\Ab�7|U�D�A��>(����iݾ]b���6e����B�����%�*R=.��=�9�=���=��=�M�=��=)��=�q�=:/�=�+�=���=J�=e�=e=Lg@=�#=>�=���<�o�<��<`_<�rL<P�Q<�   �   X~x<D��<�o�<���<ڗ<PD<��*�֋#�4y��f�/X�j	��L�ɾ!�����,�/��AB��$N�"WR�`fN��B��Z0��G���ȾK	��t�L�����6jc���7���=0��=M��=ru�=��=�}�=���=��=���=b�=�g�=��=�b=��3=�
=��<P*�<XhM<��<`�;���;p��;v<�q8<�   �   0�u<4��<��<���<���<�%�<`/S;�����yx��佈�3����,D����۾?����P*���4�L�8�l-5���*�!��� �o�ݾ?������..�@}̽��(� v�;�/=��=k�=&��=,��=:��=r��=T�=��=U�=D/`=�C"=0W�<@�C< fw:�z��V����� 텼�fm�X�0�`W�� +:P,�;�   �   �	Q<x�<��= �=�=�E=��<�0g����e����
��^N��M��
���s@ݾ=~ ���������߾�r��y(�q+�'������#�S��������Ӽ�y<�PA=Rݐ=^�=`��=x�=���=;S�=�2�=�`r=��(=x�<@�";����4� ��3��:U��e�j�c�dR�Hq4�����D�� �7��Y�:�   �   ���;4չ<RR=�1=�,@=��5=�C=贉< (�Z�@����"���PX�Wۍ������̾[�"�����������a��F�Ѿ4���͔�ܲf��&���ս�\�@-4����<:�N=�ߎ=�է=��=�.�=��=�ى=h�M=<��<���;i��R9�����|鳽ZѽL�h��.�ܽz�Ƚ���>~��.D�4�꼀]#��   �   �j��<�=�hF= �b=��f=x&N=r�=p�z< n���V���ǽ4���N�q?�������U���{��C�������,��9����)���^c�y.�L�����2V��N;X��<^
U=k7�=�Q�=�=��=��y=�K2=Tϧ<��l��E����&ս4���"���3�u�<�<�#�2��a!��5
�pj޽i��&W��Լ�   �   ��y��H<8�=�tR=h�~=%��=�]�=L�c=�&!=�S�<P�d���K�nX��:��6`2��3Y�*�x��,�����Rn���Ԃ��l�7�J��}$�����\N���A�0�y���H<��=�sR=��~=Ʊ�=�[�=R�c=j !=�C�<`�d�<L��_�����Ee2�n9Y�7�x��/��,���aq��qׂ�l���J�P�$������R����A��   �   �Z��#;��<�
U=8�=�R�=��=H��=T�y=�R2=��<�����y��[սj���"���3�$�<��<�]�2�k]!�,2
�|d޽�褽�W���Լ �(��<��=�gF=��b=f�f=:"N=��=Їz<#n���V���ǽY��
�N�FB�����bY��|�����������/��!���w,��cc�@|.�4��Y���   �   �\�0:4����<�N=+��=�֧= �=k0�=� �=�܉=ЋM=@��<��; P��9�����#᳽xQѽC�#�彃�ܽ��ȽJ����y�� D�$�꼰P#����;�չ<�Q=T�1=*@=z�5=>?=���<�/(���@��������6UX��ݍ���M;�
���������e���׌�b�Ѿ�6���ϔ�d�f��&���ս�   �   D
�� �Ӽxy<�OA=�ݐ=$_�=h��=��=���=�U�=�5�=hr=R�(=h"�< =#;����� ��v3�h-U��e��wc��YR��h4����4:��0�7� ��:�Q<��<`�=��=D�=6B= �<��g�����ã��
�AbN�-P������Cݾ� ����n�l�����-��*�%.�f��������S� ���   �   �̽�(��f�;6�/=��=�k�=���=L��=���=\��=]V�=u�=gX�=�6`=rL"=�i�<��C<��y:@+��YV��邼�݅�XMm���0� ;�� �+: 5�;��u<���<0��<���<|��<0�<`�R;����@�x�A�@�3����CF��n�۾������*���4��8�$/5���*��������ݾ�@��T����0.��   �   ���� mc��7�<�=*��=���=v�=��=�~�=^��=���=���=��=�j�=0��=�#b=��3=�
=��<�7�<X�M<p�<�2�;स;@�;{<@s8<H}x<l��<�l�<��<\՗<�8<�*�`�#�|���g��X��
���ɾB�������/�CB�<&N��XR��gN�H�B��[0�' � ��V�Ⱦ[
���L��   �   [��1�����%��Q=/��=�9�=X��=V�=�N�=Η�=J��=s�=�0�=�-�=���=<L�=<g�=�e=�k@=(=��=��<u�<d��<`#_<HuL<��Q<��j<t&�<�L�<��<`�7< ���:���Z�&˽\�$��t�*��$�V��Dh(��oA�QU�D"b���f�fBb�.}U��A�f?(����jݾc���7e��   �   V������u�F=.l�=L��=ǧ�=5�=d>̿>� >���=���=���=6�=D۳=5�=Ԍ=
*t=�?P=4.=4�=x��<H�<�$�<��o<ЁZ<x�[<�|g<�[k<��L< #�;�ɻ�6弼�|��G�G�2����M˵�&x"�Xn2�b�L��a�[�n�֐s���n���a�
�L���1��!���_����u��   �   ��������Ĉ�T,�<���=`��=���=���=��>:c>��>#��=���=<=�=��=��=짨=%j�=υ�=@<`="�<=�0=D�<�j�<dW�<({z<�)\<yU<X�Z<�Y<`�5<0Ŝ;��� o��!i����轪�7�����͹��m����5�P�B�e��Qs��x��Rs���e�rPP��K5�f�������$�z��   �   2��O��`�u�=�l�=���=��=:5�=)d>ۿ>"� >���=���=���="6�=g۳=>5�=<Ԍ=�*t=2@P=�4.=6�=���<��<�'�<��o<��Z<ؘ[< �g<�ck<��L< 4�;��ɻ�1弔�|��E��2��~��Hʵ��v��!�ym2�g�L�p�a�>�n���s���n���a��L���1�!����f���Vu��   �   0�������%�U=[��=�:�=���=��=�N�=��=x��=8s�=�0�=�-�=���=|L�=�g�=`e=�l@=h)=��=���<xy�<���<�._<��L<R<�j<�-�<HT�<0�<��7<�t��0���Z�O"˽�$��t�((�����~��f(�nA�OU�& b�Z�f�J@b�.{U�I�A��=(����gݾAa��5e��   �   ����dc��C7���=Ԙ�=���=�v�=:�=�=���=ܢ�=���=
�=�j�=u��=.$b=V�3=
=��<�:�< �M<��<�K�;0��;�'�;Ќ< �8<ؐx<���<`w�<ļ�<���<pQ<��*��#��v���d�BX�5��ɦɾN�������/�P@B�M#N��UR��dN���B�SY0���$��"�Ⱦ����L��   �   �x̽H�(�P��;��/=��=�l�=���=���=9��=���=�V�=��=�X�=p7`=
M"=\k�<��C< ;z:@���PV�`䂼�ׅ��>m�`�0������,:�a�;@�u<�ǲ<� �<l��<@��<4.�<�uS;����sx�B�,�3�U��UB����۾�������*�:�4���8��+5�I�*��������ݾ�<��F����+.��   �   p����Ӽ��y<,VA=�ߐ=�`�=���=��=b��=V�=�5�=�hr=�(=�#�< G#;`���� �Bu3��+U���d��tc�8VR��d4�6���/��8�7��`�:�&Q<0%�<,�=$�=�=~J=�<@�f���A���s�
�][N��K�������=ݾ�| ����������������&�Y(�p����
��J�S�ۑ��   �   �[�x
4�P��<P�N=s�=Mا=A	�=21�=�!�=B݉=t�M=t��< �;�N��t 9�j����೽�Pѽ�B���#�ܽ��ȽJ���@w���D�p�꼘7#�p�;|�<�X=��1=�1@=�5=I=���<��'���@�����̃��LX��؍�����̾��Z������٩�������Ѿ�0���ʔ�*�f��&�)�ս�   �   �K���;��<�U=H:�=8T�=��=��=h�y=�S2=�< ����ty��ս<��d"�V�3���<�n<���2��\!�<1
�Kb޽K椽VW��Լ�K�DÜ<��=�nF=�c=җf=�+N=h�=h�z<�m��V�^�ǽF��n�N��<��ޢ���R��[x������y�=)��󧡾�&���Yc�xt.��	��u���   �   (�y�8�H<�=`zR=��~=���=�^�=��c=�'!=TU�<��d�^�K�0X����`2��3Y���x��,������n��RԂ�Gl�c�J��|$������K����A��y�ȩH< �=�zR=��~=���=v`�= �c=l-!=�c�<x�d��K�?Q�����H[2�A.Y��x�k)������k��jт�l�ȩJ��x$�s���+G����A��   �   ��꺠Ɯ<��=�mF=��b="�f=2(N=��=�z<`�m���V���ǽ���N�e?��奚��U���{��$����󽾋,��򪡾�)��"^c�x.� ��~��Q�@�;x��<FU=�:�=U�=�=� �=f�y=.Z2=<�<�W����Or���ս���b"��3�n�<�:
<�ؐ2�:X!�f-
��[޽E᤽�W�p�Լ�   �    /�;��<4X=H�1=�/@=�5=0E=ඉ<(�Σ@�ߑ�����PX�Nۍ������̾N������������8���Ѿ�3��8͔��f��&���սr�[� 4�p��<P�N=��=�ا=X
�=�2�=�#�=�߉=P�M=<��<�f�;7����8��苽tس�FHѽ	:⽬��L�ܽ��Ƚ5���Br����C����h(#��   �   H+Q<`%�<T�=��=| =nG=d��<`$g�"��)�����
��^N��M�����k@ݾ9~ ������}��վ�d��e(�@+�籹����o�S�8�������ӼP�y<�TA=�ߐ=a�=N��=��=��=FX�=�8�=|or=�(=�6�<`�#;`|��6� ��g3�6U���d��hc�dKR�H[4����4$���7�@��:�   �   �u<ǲ<\��<���<���<�(�<�=S;ԥ��yx���t�3����%D����۾=����N*��4�I�8�h-5���*���} �@�ݾ�>��ɒ��I..��{̽��(����;B�/=��=m�=t��=��=���=m��=�X�=[�=�[�=�>`=VU"=�}�<��C< �|:��� *V�`҂��ǅ�`#m���0� �����-:n�;�   �   ��x<l��<u�<���<�ܗ<H<0�*�j�#�y��f� X�e	��F�ɾ�����*�/��AB��$N�!WR�^fN��B��Z0��)��́Ⱦ	���L�����6hc��n7�X�=x��=���=&w�=��=
��=���=j��=���=L�=�m�=j��=�*b=@�3=(#
=�'�<�H�<p�M<H<0q�; ߸;p=�;��<h�8<�   �   ��j<�,�<�R�<��<��7<����4��8Z��#˽�$�L�t��(���ྉ�Zg(��nA�PU�,!b�g�f�[Ab�5|U�@�A��>(����	iݾCb���6e�X�������%��S=��=�:�=��=�=^O�=̘�=|��=lt�=n2�=l/�=ʈ�=�N�=�i�=� e=@q@=�-=��=���<l�<P�<�5_< �L<�R<�   �   ��[< �g<�ak< �L<�.�;��ɻ43弈�|�dF�h�2�,���ʵ�Ww�"��m2�ЮL��a���n�D�s�\�n�2�a���L�b�1�~!�������Ku����_��`�u�=�l�=���=��=\5�=Hd>�>_� >&��=���=���=7�=jܳ=R6�=ZՌ=�,t=`BP=�6.=��=���<L�<�)�<��o<��Z<�   �   ��@=�k==��.=�=��< ò��0��*ƽBL.�z8���6ž���Sc.���W�����ґ�mޟ�ᨿ����Zᨿ_ӟ�.���]�a�V���,�%������}�ԍ�;̅��V`� �.=N7�=O��=���=���=|�=���=���=�"�=��=B�=��=Չ�=(�=�t=��^=��M=0�A=R):=�6=:�6=�9=��==�   �   z�==�==`0="�=�<��k�L�%�9/����)�k	���������+���S��g{��?���������
��B���H��>&����z��R�-�)�~��o����Nx����䃀� ��(2=©�=X��=���=2��=�=T��=>V�=:��=�v�=X,�=D�==�=��v=�\=��G=�8=(�.=0�)=�)=z#,=��1=��8=�   �   4\5=n%;=��4=�u=p4�<��:���檽�����w��մ�+���`!��KH�&n��ć�0������hv���������Ї���m�q�G��H �rv��c��J�g�$��xb�@G4;P�;=/��=Ȟ�=�g�=�Q�=�+�=�k�=�T�=���=�)�=���=�5y=�aQ=��/=nO=��=P�<4��<hs�<D|�<�5=��=��(=�   �   ��$=��5=�P9=D�(=� �< /$<�l���,���V�`�Z��ۡ���߾+H��46�Y��x�U���<��t��@d��q�����x��gY�,46�u��Pݾ靾GaN����jH3���<��I=b��=�2�=5��=���=8��=":�=N��=�<�=l9x=�.?=�C	=P�<�P< 0�;��*;�H�:��m;��;H�W<�]�<�<�<�=�   �   ZN	=�0*=��;=��7= �=Xr�<�𻘝E�?ֽ-@6�ԉ������G��;�u>�PZ�bp���~��݁���-q�`B[��\?����X����}��*凾�U.����%�ܱ�<��Y=7��=�ٺ=Ax�={��=��=���=�C�=M@=�]�<�B)<�Pػ0��
��R$���'�����Z�|ɼ(�_� �ƺ�3<�!�<�   �   �ٽ<��=xF8=��D=��4=��=8�<��ԼV���N�]��9��n%Ӿ�L��Y ��8�5�K��@X�t�\���X���L���9���!�}���վO	��D�^��
�9���@ya��Q�<@9h=PI�=���=.��=��=�o�=L�^=
=��(<��l��-�^�z��D������Bͽ��ν�5ý����J��KP��L � @� 	�;�   �   �	<��<(,= �L=�`O=��/=4��<�R2��/�10ĽHU%�ۊt��o����Ծ���b�h�%�V,0�G4���0�'�!U��Y���پ<Y��~}��|,���̽R=1� ��:�!=@�r=�Ε=:7�=�ә=�=X@= ��<Pݟ����B鎽��ѽ�@�" �gE1��n9�L8�Ջ-�&���6ͽ�\���,��t{��   �   8;<�h�<`�=$bL=jgd=��Y=,�)=Tz�<��D��#`�bݽ�.� v�����GIžMZ澤i ��	�l��	
�6�qv�R�˾D���Ȣ��*�=��Q��l������(�<\�.=2+v=�g�=�Ћ=�s=��-=|��<�i�U�����m����9�b�G��R>��k�����fԆ�j`r���N�ٖ&�����3���B�4��   �   2�� ��ܺ�<�zB=�q=B{}=�"e=μ'=���<�Ԇ�2�n��Jܽ�V&��Ja�=�����������Çʾ�о��̾����%��	ӕ�&�t���;��e�Xv��|�����|��<>{B=��q=�x}=e=4�'=|u�<�膼�n�Sܽ�[&�uPa�����`���ĝ���ʾMо%�̾���l)��,֕�e�t��;��h�&{���   �   K��̚��,��<.�.=�+v=�h�=�ҋ=֤s=��-=��< �h�U����^����9��b��C���:����y	��
ц�ZZr�z�N�n�&�������J�4�H%<���<�=*bL=�ed=��Y=��)=�m�<�E�/`��	ݽz�.��v�ߎ�� Mž�^��k �	�sn�&
�R8�z�ڜ˾:���*�����=�`W���   �   ��̽�B1�@�:R =*�r=Yϕ=�8�=�ՙ=���=�@=�Ͽ<p����������g�ѽ�;�o �y?1��h9��8�f�-�9!�Ҷ��̽8W��n�,�p[{�H&	<���<�,=|�L=�^O=d�/=���<@�2���/�6ĽY%���t��r��u�Ծ�� e�ߛ%��.0��4�P�0�h'�HW��[�ٻپ�[���}��,��   �   5�
������a�N�<�8h=�I�=�¯=ť�=��=�r�=��^=l
=h�(<P�l���ćz��;��S����8ͽ��νM-ý����[D��(@P��C ���?�`.�;�߽<��=�F8=��D=j�4=6}= �<�Լ�Z��
�"�]�<��k(ӾjN��[ �d�8���K�aCX��\�"�X��L���9���!�����վI��>�^��   �   �W.�m����,�4��<�Y=t��=�ں=|y�=?��=h��=���=+G�=�U@=�q�<`p)<��׻����D����8�'����O�ɼv_���ź��3<�(�<XP	=\1*=p�;=^�7=ؔ=�k�<��أE�jֽ�B6��Չ�E���}J���<�w>�?RZ�Kdp��~��ށ�^�0q�UD[��^?�H����������懾�   �   �bN����0K3�H�<�I=���=03�=��=���=���=D<�=���=�?�=�@x=�6?=�L	=D��<�CP<�}�;@f+;�_�: 8n;�T�;p�W<�f�<�B�<0�=�$=��5=hP9=�(=���<p#$<�t��C/��|X���Z�'ݡ��߾aI�D66��Y��!x�V���=��r��6e��V���&�x�IiY�]56�n��рݾ6Ꝿ�   �   \�g���dzb��74;�;=P��= ��=$h�=`R�=�,�=Ym�=EV�=���=,�=���=^;y=�gQ="�/=�U=��=L�<��<�{�<��<�8=`�= �(=�\5=|%;=
�4=�t=X1�<@��:���誽�����w��ִ�����a!�MH�^n�AŇ��������� w������^��Fч���m�C�G�0I �zw���c���   �   Ox�ҕ�/���  ��(2=꩛=���= ��=���=��=��=W�=>��=.x�=�-�=��=�>�=�w=�\=��G=��8=x�.=�)=8)=�$,=J�1=(�8=��==t==�_0=t�=�<@l�6�%��0��h�)��	��E��@��g+��S�Vh{�/@����������
����������&��v�z�g�R�y�)���������   �   ��}�����˅��L`���.=�7�=|��=��=���=��=���=���=�"�=��=P�=	��=㉖=(�=�t=n�^=��M=�A=$):=޲6=�6=��9=n�==j�@=jk==��.=�=��<�Ʋ��0��*ƽ�L.��8���6žƅ�rc.���W�����ґ�xޟ�ᨿ����VᨿYӟ�%����\�D�V��,��$�̀���   �   �Mx�����������n*2=v��=���=g��=���=��=%��=6W�=R��=:x�=�-�=��=�>�=�w=:�\=��G=4�8= �.=�)=()=�%,=d�1=V�8=��==�==2a0=�=��<`�k�^�%��.��,�)�+	��5������+�|�S�+g{��?�����*���<
����������%��S�z�k�R���)��������   �   s�g���@tb�`}4;
�;=_��=ޟ�=�h�=�R�=-�=�m�=pV�=���=.,�=���=�;y=LhQ=��/=8V=��=T�<���<�~�<���<|:=��=l�(=F_5=(;=�4=�w=�8�<�L�:B���䪽���z�w��Դ���`!�KH�&n�ć�����%���u��M�����Ї���m�d�G��G ��t���a���   �   �^N��轠B3���<F�I=���=14�=���=p��=F��=�<�=��=@�=Ax=*7?=RM	=T��<�FP<Є�; x+;���:�Sn;e�;ثW<�k�<�H�<b�=��$=��5=dT9=v�(=��<�;$<Le��Y*��:U�}�Z�[ڡ�\�߾*G��36��Y�x�-T���;��z��Fc��~�����x�CfY��26�D��X}ݾ�睾�   �   �R.�R﻽$�м�<0�Y=<��=�ۺ=Qz�=���=΅�=܇�=jG�=.V@=�r�< r)<��׻@���~�����'�^���M�H�ȼ�j_�@�ź�3<40�<zT	=�5*=8�;=��7=��=�z�< �� �E��ֽ�=6��҉����6E���9�[s>�$NZ��_p�r�~��܁����+q�F@[�[?�,�������{��Vㇾ�   �   ��
�_����Za�(^�<x>h=�K�=�ï=���=^�=�r�=v�^=�
=@�(<��l�>�H�z��;��艾�S8ͽ�νj,ýs���C��=P�v@ �8�?� P�;��<L�=�K8=��D=.�4=Z�=X�<�}ԼR��|��]�n7���"Ӿ K��W ��8���K�S>X���\��X�R�L�>�9���!�����վ���P�^��   �   R�̽<31����:�(=��r=[ѕ=�9�=�֙=���=�@=ѿ<0|��������.�ѽ};�J �J?1��h9�-8���-�� �*����̽~U����,�XJ{��8	<���<`,=��L=�eO=Ĭ/=��<��1���/��*Ľ�Q%�t�t�<m����Ծ�
��`��%��)0��4�6�0��'��R��W��پ1V��y}��x,��   �   5���|��H�<$�.=41v=wj�=�Ӌ=��s=��-=���<��h��U�����H����9�ub��C���:����S	���І��Yr���N���&�$���䌦�<�4��<���< �=hL=�ld=��Y=�*=���<��D�z`���ܽ��.��v�i����Ež&V�^g �3	��i�S
��3�r�e�˾֮��⟂�`�=�"J���   �   Į��C�8��< �B=�q=�~}=|%e=j�'=�<0ӆ���n��Jܽ�V&�sJa�4�������������ʾ�о��̾����%���ҕ���t��;��d��t����������<��B=P�q=��}=�(e=6�'=P��<,����n�HCܽR&��Da�񈍾Л������p�ʾ�о��̾����!��ϕ���t�h�;�<a�!o���   �   ��;�@�<b�=�hL=�kd=��Y=P�)=(}�< �D�F#`�'ݽ٠.�v�����@IžEZ澞i ��	��k��	
�6�Gv��˾���z���t�=�MP���
��������<4�.=�0v=k�=(Ջ=Īs=��-=|��<سh���T��������9�2b�@���6���쐾���h͆��Sr�_�N��&���������P�4��   �   �K	<���<�,=��L=�dO=H�/=���<@@2��/��/Ľ/U%�Ȋt��o����Ծ���b�d�%�T,0�C4���0��'�U��Y��پ�X���}}�|,�9�̽:1� ��:&= �r=�ѕ=�:�=�ؙ=���=0"@=<�<�%�����؎��ѽ^6�� �n91��b9�V8�r�-�������̽hO���,�P.{��   �   �<Z�=�L8=\�D=��4=��=��<ĈԼ�U����;�]��9��f%Ӿ�L��Y ��8�4�K��@X�r�\���X���L�|�9���!�k����վ	��­^���
���ma��X�<>=h=�K�=�į=��=W�=�u�=j�^=�"
=`�(<p`l���0wz��2��ʀ��/ͽ��ν�#ý����:<���1P�7 �8�?�0z�;�   �   �V	=7*=v�;=
�7=f�=�u�<p���E�ֽ@6�ԉ������G��;�u>�PZ�bp���~��݁���-q�ZB[��\?����8����}���䇾IU.���t!� ��<��Y=%��=$ܺ=D{�=F��=އ�=���=�J�=@^@=���<��)<��׻(ޫ�҇���j�'�����A���ȼhH_���ĺX�3<�7�<�   �   �$=N�5=`T9=ƃ(=��<�3$< k��P,���V�T�Z��ۡ��߾)H��46�Y��x�U���<��u��@d��p�����x��gY�%46�k��4ݾ�蝾�`N����F3��<��I=Ĳ�=j4�=h��=|��=���=r>�=���=�B�=�Gx=�>?=�U	=��< mP<���; ,;���:`�n;@��;��W<�u�<8P�<��=�   �   >`5=�(;=Б4=dw=�6�< !�:"���媽�����w��մ�)���`!��KH�%n��ć�2������gv���������Ї���m�k�G�H �bv��c���g����wb� [4;��;=��=��=i�=^S�=.�=�n�=�W�=���=`.�=8��=8Ay=0nQ=ư/=n\=��=�'�<���<��<4��<�==޺=�(=�   �   z�====6a0=�=�< �k��%�$/����)�h	���������+���S��g{��?���������
��A���G��>&����z��R�)�)�z��e����Nx�v������ �~)2=7��=���=���=��=7�=���=�W�=4��=Dy�=�.�=�=@�=�w=B�\=��G= �8=��.=$�)=)=.',=��1=.�8=�   �   x�=�m�=ڥk="K3=���<Tޅ� ���Z���{�п���v	�E9�"�m�潑�㏫��_¿�YԿ��߿L��S�߿�GԿ�$¿������,�k��6�q������*gj�Rt���_4���n<�;f=d¬=�~�=��=u�=*$�=I��=��=.Ų=`Þ=R��=v=r%[=�H=�"==.:=�v>=��H=�iW=�uh=�y=_��=�   �   \у="ȁ=rk=�S5=f�<�k��(�����u�ՠ��g����5�MRi�,�����U��&�п@*ܿ��1ܿ=�п�쾿�?��X���@�g��3�t��쵾1e�_1���)+�8��<�h=�0�=D��=���=�^�=���=29�=�ͼ=�=�s�=�S|=T�X=�<=О)=�g=V=س$=p�1=H�C=~yX=\m=�B~=�   �   ��t=Ry=țh=��:=���<�=�F�o����od�_�������+�+�V�\��������}���jƿ%Nѿ�տ�jѿ��ƿ�����㟿�[���[���)�����ת�kZU�_�0{���<��l=VB�=��=ȅ�==��=6�=İ�=.v�=Yʆ=��Y=2S)=��<8��<p��<(V�<Xj�<PL�<8�<08=\p'=@�F=J�a=�   �   �R=�e=<�b=��A=���< ~����:�B���OI�5����o���I�x����'~���4���S��
�ÿ�������Ѧ�������w���H�y��`��}�����<�|5��P�μ` �<�s=�N�=�ڽ=b�=l�=p�=Tt�=(�_=p�=�Я<�V�; ӻ����4k��Xe��TG��P�O��:[��k<�@�<B�=0=�   �   �&=��F=�ZV=��F=��=��(<���*�� �&�т��ož^��j&0�I6Z��b��<Z��<���Ԭ���� �����`$偿��Z��l0��Q���þq������ؖ��tP���<Fx=�d�=˭=���=�֘=ֺv=4*=�g�<�1�H�ͼ�{:�:#��������e����@���V��f�B�X��H�1�p��;�'�<�   �   �Ƭ<�=��@=�G=�z'=���<h�2��Er��C �rX�
,�����T���m8���[�z'{�&�������씿�d��أ����|�.[]�I�9���:��L����QV��<���Q���`:�=F^y=(��=+r�="-�=�dR=Ph�<�Z;�Xټ,>m�X������܃�H^���%�ϫ#���n��~ ޽?����Z���Ҽ �ٹ�   �   �"/�0�<��=��@=6+:=Np=���;�� �|H���$!�PR{�튲� 8��5��2���M��b�>@p��@u�9q�|d�bpO��5�"O�0	�'���o��l�#�:����.� �h<2�0=�Et=별=�&t=�!8=�8�<0��^�:�{=��ґ��/���V�%�u��w���߉��Ї�:-��d�kA��<��߽�Վ�B�	��   �   �����:���<6n/=��E=�/=��<��tKD�$t׽(m4��ބ��B��9�很�|� ��2��R=���A��3>�I�3��#����Mm�jԹ��!����=����@Z����|U�<f�@=�f=D�^=0�*= ��< yl��f�9�ؽ��$��`�������������ɾ�mϾ̾�&������k���Iq���7��2 �� ���   �   ���j����?<��=�3H=��O=��(=x��<0>O�^�i��Q��5�T��mߦ�*�̾��5��0�v���#��
�k;���0Ӿ���v����D��������\��ؑ?<��=�3H=��O=z�(=P��<xcO���i�Z�F�5��
��R㦾��̾�~8�h3�Y��b&�M�A@���4Ӿs񭾉y��|�D�(���   �   S���Z���综P�<�@=��f=ʲ^=҆*=8��<�Ml���f�>�ؽ%�$��_�)������Q����ɾiϾ�̾j"������dh���Cq��7��. �����n� m�:ث�<Ho/=ܽE=��.=���<0����UD�,{׽�q4��ᄾ�F������N� ��2�V=�3�A��6>�@�3�W#����Pq뾬׹�l$��V�=��   �   _�#�N����8鼰�h<b�0=�Ft=K��=L+t=x(8=�J�<8����:�o4��q��؝/��|V���u��s���ۉ��̇��%�5d��A��7��w߽�ώ���	���.��$�<��=��@=�):=m=�w�;�� �N���(!�@W{�����;�B8���2���M��b��Cp�Du��q��d�6sO�n5�>Q����õ�z���   �   �TV��@��N�Q� `:��=�^y=1��=�s�=�/�=HlR=${�<��Z; <ټF-m�����ڦ�~�1X���%�Х#�L�L���ݽ� ��(�Z���Ҽ ֹ�Ь<	=��@=��G="y'=�<P�2��Mr��F �:X��.�����H��'p8�l�[�p*{�����,���Mf��]���t�|��]]�]�9������T����   �   ɯ��{�ۖ��P���<~x=�e�=|̭=���=�٘=�v==*=�}�<@H0��ͼlk:��������򣽂���c8��JO��}B����H�1����;�2�<`*=��F=R[V=V�F=��=�r(<X�������&�����mqž݇�A(0�v8Z��c���[������V���򭿙���h���A恿u�Z�fn0�(S���þ�   �   ����a�<�q7���μX��<�s=CO�=�۽=��=,n�=�=�w�=�_=��=��<0��;�һP怼�Q���L���/����O�@�Z���<�M�<<�=�0=��R=:�e=z�b=2�A=��< ��L�:���� RI�����侺��d I��x����N��6���T��O�ÿ=�������(Ҧ�忒���w��H�{�����   �   Mت�k[U��ὦ|���<�l=�B�=T��=Ɇ�=���=��=䲷=�x�=L͆=\�Y=�Z)=� =\��<���<�e�< y�<�Y�<��<.==dt'=R�F=��a=�t=y=h=��:=̤�<�G���o�d���qd�����6���'�+���\�d�������~���kƿOѿ�տ�kѿt�ƿv����䟿\��ƚ[�\�)�����   �   �쵾�e��1��Z*+�4��<�h= 1�=���=���=�_�=h��=M:�=ϼ=|�=�u�=NW|=(�X=��<=��)=lk=�=�$=4�1=��C=T{X=�m=�C~=�у=>ȁ=Jk=>S5=�c�<��k�"*����+�u�����߹�V�5� Si�|,�����������п�*ܿ��O2ܿ��п��?��������g�a�3����   �   d����fj��s��
_4��n<�;f=�¬=�~�="��=��=D$�=c��=��=@Ų=rÞ=_��=*v=x%[=�H=�"==�-:=�v>=��H=�iW=�uh=��y=C��=`�=gm�=��k=�J3=���<�߅�����Z��{�����v	�*E9�K�m����������_¿�YԿ��߿L��P�߿�GԿ�$¿���m���k���6�S���   �   �뵾e��/���'+���<4h=�1�=���=���=�_�=y��=b:�=%ϼ=��=�u�=fW|=N�X=*�<=�)=�k=8=x�$=��1=0�C=|X=|m=�D~="҃=�ȁ=�k=�T5=�g�<��k��(������u�����-��r�5��Qi��+�����������п�)ܿ��_1ܿ��пN쾿?��������g���3����   �   c֪��XU���w�@�<��l=�C�=���=+��=���= �=��=�x�=`͆=��Y=�Z)= =���<d��<�f�<dz�<D[�<��<R>=�u'=ʗF="�a=ܓt=y=�h=��:=��<5���o�@���nd���������u�+�o�\�&���b��C}��jƿFMѿ�տjѿĎƿ苵�*㟿�Z����[���)�M���   �   틙���<��1���{μ��<v	s={P�=�ܽ=n�=�n�=X�=�w�=V�_=ز=�<���;@�һx值�P��K��.��H�O�`�Z���<<Q�<@�=0=
�R=�e=¤b=,�A= ��< Ђ���:����NI� ��n��e���I�nx����}���3��|R����ÿÉ��f����Ϧ�����-�w��H�4��\���   �   ������pԖ��ZP�X&�<�x=-g�=vͭ=L��=Cژ=��v=�=*=T~�<`C0���ͼ"k:�z�X���������7���N��x{B�~���1� ��;�7�<d-=�F=J_V=, G=��=�(<l���	����&�S���mž���$0�Z4Z��a���X��م��\���	ﭿ�����	��퓿�みk�Z�k0�rP���þ�   �   �MV��6����Q� �b:��=�cy=Ԃ�=u�=�0�=6mR=`|�< �Z;P;ټ�,m��������}�X�n�%���#�������ݽ�����~Z�X�Ҽ �Թ�׬<�=F�@=�G=�'=8��<��2�L>r�wA �*X��)��Ĝᾑ���k8�F�[��${��������;딿c��F�����|��X]���9����������   �   ��#�1������h<��0=�Kt=���=�-t=�)8=�L�<����:�B4��^��ǝ/��|V���u��s��~ۉ��̇��%��d�5A�o7��v߽gΎ���	� �.�L,�<f�=h�@=�0:=�u=���;ܫ �bC���!!��M{����o4��3���2��}M�Ҏb��<p�R=u��q�Hd�imO�C5��L�C���������   �   ;��z�Y�`I��d�<�@=`�f=�^=�*= ė<�Il�J�f��ؽ�$���_�"������J����ɾ�hϾ�̾M"������4h��Cq���7�. �����@����:`��<�t/=x�E=d/=��<0@��xAD��m׽�h4�܄��?��!��"��� ��
2��O=��A��0>�=�3��#����h뾳й������=��   �   ����F��p�?<�=>:H=n�O=��(=T��< 9O���i��Q���5�L��fߦ�'�̾��5��0�q���#��
�L;���0Ӿ��dv��d�D������,V����?<r�=�9H=��O=�(=t��<�O�Zyi�J��5�I���ۦ���̾&�3��-����� ���P6��$,Ӿ�魾Hs��s�D�T���   �   ������:d��<hv/=l�E=�/=�
�<�q��hJD��s׽m4��ބ��B��4�径�z� ��2��R=���A��3>�B�3��#����&m�8Թ��!����=����b�Y�Px�^�<��@=(�f=��^=��*=җ<�"l�T�f���ؽ��$���_�z񌾃�����!�ɾdϾ��˾�������xd���<q�G�7��) �7��   �   �.��6�<d�=��@=0:=�s= ��;V� �H���$!�<R{�劲��7��5��2���M��b�=@p��@u�7q�vd�YpO��5�O�
	�����6����#�	����(鼀�h<��0=�Kt=���=`1t=�/8= ]�<�w�d�:��+��B��җ/��uV�6�u��o���׉��ȇ�>�d�.A�G2�Un߽�ǎ���	��   �   ��<�=b�@=��G=�~'=0��<��2��Dr��C �WX��+�����P���m8���[�z'{�&�������씿�d��أ����|�'[]�=�9����� ���PQV��;����Q���a:��=Xcy=x��=�v�=�2�=�sR=���<��[;| ټ�m�)���8��;x�R�K�%���#�H����X�ݽ�����qZ�`�Ҽ �й�   �   �1=��F=�`V=J G=��=h�(<@�������&�Ȃ��ož[��i&0�H6Z��b��=Z��<���Ӭ���� �����_"偿��Z��l0��Q���þJ���B��ז�XkP��!�<Bx=�g�=�έ=��=�ܘ=R�v=�E*=В�<��/�p�ͼp[:�z �c����飽"���[/���F���mB�,f�Pw1�0*�;�C�<�   �   ��R=��e=��b= �A=��< ȃ���:��ཾOI�.����n���I�x����'~���4���S���ÿ�������Ѧ�������w���H�r��I��`�����<��4���μ��<�s=�P�=|ݽ=��=Pp�=��=�z�=��_=~�=���<��;�Pһ\̀�7���1��8��@xO���Y���< _�<ڎ=80=�   �   ĕt=Hy=��h=��:=���< :���o����od�[�������*�+�U�\��������}���jƿ&Nѿ�տ�jѿ��ƿ�����㟿�[���[���)�����ת�@ZU���z���<��l=�C�=S��=���=���=��=�=3{�=%І=ҿY=�a)=�
 =���<���<�v�<���<Li�<\�<�C=$z'=d�F=��a=�   �   �҃=Ɂ=�k=�T5=Tg�<h�k��(�����u�ՠ��f����5�LRi�,�����V��&�п@*ܿ��1ܿ>�п�쾿�?��X���=�g��3�p��쵾e�*1��n)+����<�h=z1�=��=��=1`�=-��=C;�=@м=��=!w�=�Z|=��X=��<=Ҧ)=�o=�=�$=��1=��C=D~X=Pm=
F~=�   �   �=�~�="=~=Jg0= �8<<���ܽ�S��������6�P�s�Ȯ��~:���Sܿ����%���������ƭ�Yu����ۿtI������j�p�#�3������=��\�C��B��t򍼬�=(1�=�v�=p��=?��=(��=���=��=���=��}=T=�1=�.=/=(�=��=��=~�5=�S=�Wr=ć=w�=�   �    �=^��=��{=Jm1=`oK<����ս��M��S������K3��o�P������:�ؿ���0y�!���:�~���u��n��Iؿ�5���햿�l��0�0���ͼ����>�{)��`���B=U��=sB�=���=�-�=�w�=�4�=ʋ�=^I�=�_=�t2=��=0��<��<�<O�<��<b&=Э9=�]=�x~=Sc�=�   �   �˄=н�=�;t=��3=��<`5�Hi���>�`���rﾜ7)��Hb�(��u�����Ϳ@����������6����a��8�还�Ϳ�=���a���j`�g'�Bg����1�2����I0���=��=�n�=�=��=���=Ǟ�=��{=v?=��=쓖<0��;��)��֜��"���pt�;�{w<l�<`=�@J=��p=�   �   ��W=��m=J�e=ر5=�6�<����Ρ���&�IT��w�׾A���6N�A̓��"���,��<�տ��2������������Nfֿ�n��������/"M�X�|ԾR����}��?�� 'a���=�7�=GX�=�a�=���=`Ԉ=�Q=�h=�XI<Q���8мF�#��VM�6a�t%^�kE���P��� !޻�,<h��<��+=�   �   �=h�==.3M=��3=8�<@}���t�����o�5������*�4�6h�5����ϧ��#����Ͽ&ۿ�>߿��ۿ]{п�﾿�{��U򎿖�h�2y4�#��"����i��S �$yH��*�;�i)=�~=���=$B�= �i=�j =ķ�<�V*������xr���u�Y;�� 4�6��1�D�н������d�lo��@뮻�Y�<�   �   x�!<(L�<��'=t+=�r�<��;�����νp;?�op��DU޾W��e�D���r��{�����
���.���]"��x���b�����y���Jt�ҳE�Mx�Ҍ޾G����;��ý�d��hVn<
s/=t�g=�zl=֧D=���<@e�:@e���;��srܽ���=�8��kU��th��Dp��:l��\���C��T#�����j����L��ˍ��   �   ��@�;���<�4=
J
=0s�<�P������W�g�k��꯾����o��LF���k�����ּ��0G��fh��GΜ��������=n�4}H��<!�A�������em�O�������K�Ի<6�.=H~E=�(=���<���л;�����S�,�J�,����#��\Ѭ�}չ�:�t����i��*I���
���Y�`5#���ݽ6�}��   �   z9��p=��H$1<��<��=xO�<  w;|��&#��1s(�c�Ⱥ���n��7��Ԋ9���T���j���x�
~���y��l��\W�66<��u��7���۽�hV����-�������?�;<��<�$= *=� �<`���eS���ֽ��+��s������qľ���F ������l�	�������osʾ�5���΀�k�9��3��   �   ��b�_��2��x�<��	=2y=0N�<P��C��ս2w3��q��[泾��很�
�� ���1�NH=�U�A�^@>���3� $#����e{뾑�����k=��V�_���1�p~�<��	=�v=pD�<01��,C�ۻսb|3�'u��~곾��g�
�$� ��1��K=���A��C>�`�3�'#������[¹���(p=��   �   `�-��������#�;���<P$=.=8.�<P��zXS���ֽ��+��s�Z����lľ��O ������Z�	����X���nʾ�1��sˀ�X�9�,��3��4.���61<ܑ�<>�=lI�<`�v;b���)���w(�O��������s�� ���9�]�T�g�j���x�~���y���l�7`W�=9<�yx��;��߽��X���   �   �hm��Q�%����L�Dѻ<�.=R�E=�(=�<�N�:�;�h���bM�Y�J�6���4���̬�pй�뾾w����d���D�������Y�!0#�m�ݽ��}�\Ṽ�8�;���<�5=�H
=l�<l]������Z��k������xr��OF���k�j���־��EI��~j��UМ����F����@n��H��>!�×��6����   �   4�����;�� Ľ$m��POn<Zs/=��g=�~l=F�D=���<@l ;H���2���gܽfz�\�8�4dU�1mh��<p�3l���\�8�C��N#������a����L������!<pU�<0�'=�+=�o�<���;T����ν�>?��r��lX޾\��ޛD�v�r��}����� ���8���n$��z��zd�����R{���Mt� �E�z�w�޾�   �   㰷�4i�TU ��|H���;�i)=p�~=:�=�D�=�i=js =΃<� *���ﲆ�Bh���j��/��-.���'�f�нF����d��V��𝮻<h�<"$=��==�4M=��3=|	�<Ȍ�Љt�T��7�o�y���:���4�R8h�����fѧ�j%����Ͽ�'ۿg@߿h�ۿ}п��]}���󎿎�h��z4�V���   �   �ԾQ����~�A���>a���=W8�=mY�=]c�=!��=�׈=�Q=*r=؅I<����м��#�rFM�a��^�\E�<��𓾼@�ݻ@-<���<�+=�W=��m=(�e=\�5=3�<����ѡ��&��U��p�׾���v8N�>΃��#��7.����տ��鿦3������B���6꿙gֿ�o���������t#M�Q��   �   4h꾨����1�+���0M0���=��=do�=5�=��=�¯=Z��=8�{=�"?=�=$��<0�; ^'� ���Ӣ�@������;p�w<0y�<�=�DJ=��p=�̄=r��=�;t=T�3=P�<;�wk����>�5a��tﾙ8)��Ib����Q�����ͿR�����v���7�"��f�� ��b�Ϳ.>��/b���k`�'��   �   ����
����>��)�����C=���=�B�=4��=�.�=y�=26�=\��=2K�=&�_=ly2=^�=��<���<�
�<$X�<D��<�)=�9= ]=�z~=d�=x�=���=��{=�l1=�jK<��]�ս��M�lT�������K3�� o�����8��ǣؿ�����y�s���:�ȹ��u�o���ؿG6��2d�l�S�0��   �   �����=��
�C�vB������:�=`1�=�v�=���=]��=B��=�=��=Ҝ�=�}=>T=�1=�.=/=�=��=n�=L�5=�S=�Wr=�Ç=^�=ק�=�~�=�<~=�f0=��8<	�l�ܽ�S����&����6���s�ᮚ��:���Sܿ����-������������Iu����ۿ_I��q���>�p���3��   �   J��������>��'��0���D=-��=>C�=p��=�.�=$y�=F6�=m��=:K�=8�_=zy2=p�=8��<��<�
�<�X�<���<T*=L�9=�]={~=_d�=��=��=��{=&n1=�rK<��l�սp�M�uS��N����J3�go����i��٢ؿ�����x�ٳ�W:�/��gu�	n���ؿ5���햿P�l�{�0��   �   �e�捘�c1�Á���:0��=���=p�=��=��=�¯={��=r�{=�"?=�=\��<��; R'�0���pТ��������;Мw<�z�<�=�EJ=��p=�̈́=H��=>t=(�3=��<�0��g���>�]_���q��6)��Gb����Ŷ����ͿV������T��i6���H��/�迩�Ϳ�<���`���i`�r'��   �   �Ծߩ���{�V<����`��=�9�=`Z�=�c�=���=�׈=2Q=vr=��I<@����м��#�8FM��a�4^��[E����D�����ݻ0-<̓�<��+=�W=*�m=�e=>�5=�=�<x���s̡�b�&�0S����׾<��5N�õ��!���+����տ��鿉0��n���(���F��dֿm��h���~��� M���   �   ެ��`i�4Q ��qH�P[�;�n)=
�~=d�=ZE�=�i=�s =�΃<P*���߲��/h��~j⽸/��.�g��&��н®����d�T��P���0l�<x&=��==X8M=��3=$�<�i��}t���,�o�X���|����4��3h����tΧ�$"��@�Ͽ4$ۿ�<߿��ۿ�yпEvz�� �O~h�Tw4�����   �   ܷ��m�;���ý T���qn<*y/=��g=��l=�D=���<`v ;0G���2���gܽ[z�S�8�*dU�"mh��<p��2l���\���C��N#�?���a��̟L�̳����!<�[�<�'=%+=�}�<�H�;���z�νg8?�_n���R޾���-�D�߬r�[z����%���/��S ��r���`��H��"x��Ht�^�E�Lv���޾�   �   -`m�XK�
�����K���<
�.=N�E=�(=d
�<�F껞�;�/���PM�M�J�3���1���̬�lй�뾾i����d���D�����^�Y��/#��ݽ|�}�8ܹ��Q�;���<:;=
P
=��<B��'��jT�1�k��篾��m�!JF�l�k�Ǐ��溓�'E��Of��6̜��������g:n�DzH�4:!�<���a����   �   �-��������;���<$=�1=03�<����WS���ֽ��+���s�U����lľ��N ������U�	����@�꾦nʾ�1��Dˀ��9�+�2��((���E1<��<&�=�\�<�ww;.����#o(��Z����j�����·9�f�T�ܥj���x�
~���y��l�9YW�3<�s��2���׽�iS���   �   ��6�_���1����<`�	=�~=<U�<`෻^C���սw3��q��V泾��很�
�� ���1�OH=�T�A�\@>���3��##����D{�h���Y2k=�罢�_���1�Ї�<,�	=�=�\�<����tC���ս]r3��n��~⳾O����
�ة �F�1��D=��A��<>���3�� #���]v�Z���쉾4f=��   �   y,������\1<���<��=�X�<`1w;����"��s(�X������n��7��Ԋ9���T���j���x�
~���y�މl��\W�-6<��u�y7���۽�7V��@�-��������`�;���<�$=�4=L>�<آ�zKS���ֽ��+�j�s�Z���hľ���j	 �y��h�<�	����Έ��iʾb-���ǀ�r�9��"��   �   ȹ����;��<H==�O
= {�<�K����OW�E�k��꯾����o��LF���k�����ռ��0G��eh��FΜ����}����=n�+}H��<!�"���d����dm��N�X���K��ݻ<ޖ.=t�E=$(=x�<���D�;������G���J�g�������Ǭ�r˹� 澾a���`��[@������~Y�1*#���ݽ�t}��   �   ��!<�f�<d�'=Z&+=x|�<�3�;���_�νD;?�bp��<U޾U��b�D���r��{�����
���.���`"��y���b�����y���Jt�ɳE�Ax���޾!�����;��ýH_��(fn<tx/=��g=�l=l�D=p��<�;�+��5*���]ܽtt���8��\U�leh��4p�5+l�/�\�/�C�tH#�����~X���L�h����   �   b,=��==�:M=\�3=��<�s��t����ɒo�-������(�4�6h�5����ϧ��#����Ͽ&ۿ�>߿��ۿ^{п�﾿�{��S򎿏�h�*y4������xi�US ��vH� C�;�m)=��~=��=qG�=�i=| =��<��)�������F^���_�U$��H(������нƥ��F�d�8:���<��P|�<�   �   D�W= �m=��e=��5= <�<����GΡ���&�=T��s�׾@���6N�@̓��"���,��=�տ��2�� ���������Nfֿ�n��������("M�O�eԾ8���c}��>�� a�º=�9�=([�=re�=���=�ڈ=�%Q=t{=��I<`��� м��#�`6M���`�>^�PLE�t��y��`nݻ�*-<���<~�+=�   �   τ=:��=&?t=h�3=�
�<D3��h����>�`���rﾛ7)��Hb�'��t�����ͿA����������6����a��8�还�Ϳ�=���a���j`�c'�3g������1������C0���=���=�p�=��=:	�=�į=ӣ�=�{=�)?=ڨ=췖<0N�;��$��1�� ��� �����;�w<���<�=�JJ=��p=�   �   ��=���=��{=xn1=�rK<"���ս��M��S������ K3��o�O������9�ؿ���/y�"���:�~���u��n��Gؿ�5���햿�l��0�*���ļ����>�5)������C=��=aC�=���=Z/�=�y�=V7�=���=�L�=�_=�}2=��=���<���<��<�a�<��<B.=��9=t ]=�}~=Ne�=�   �   ��=��=�Et=<�=P�������r^��͍��e�U5'��kh��R���3����鿱���=�W�(�d42�=�5��12�O�(�������|�$���@����)e�d$��Cܾ�������hT��5(<��R=�ʜ=,�=@�=f�=��=��=Zyl=X�8=��	=���< F�<�n<�Cs<<��<܌�<,�=�6=x}a=���=�r�=�   �   �=� �=�p=�'=��O����G!�t���I�ݾ#�#��+d�U����뽿{��$=�[����%��/�E`2� /�Ѷ%��q����T�俟������� a��!�r�׾;������X�K���6<��Q=yL�==䤷=c��=��=V�=��L=]=8��<�L^<��;�TO;��o;�)<y{<d@�<Ҏ=�G=��s=�"�=�   �   �=��=�d=��= Z>9��c���jE��@о��&�W�eю�Vb����ڿ�L��[��b�e$&��B)��D&�����'������ٿjk������g_U��$��%˾��w�����02��u^<�N=Ì�=���=G��=���=�s=�1=�(�<Pm<�}ݻз��*����^��(�̼8�u� ���@<X<��<F.2=nc=�   �   \�A=<i[=ּN=��=P�;*7���>�e�PA���� �D�R���u��d�ȿ������7�� ��Oh�A�����A���2�[�ȿ���������B�2C
��B��t�\�������t�<x,G=�Ƅ=Vƌ=�Հ=*�J=���<	<�}��|� v�2�`��0Z��/ ���C��ٛ���J����@o��h5�<�u=�   �   ���<��=8,=��	=��(<e��Ž2:A������U��	,�\f��h���d���п��,� �R���F
�z�/=����ѿ��o���*�e��M+�*0�j����:��̵������<�8=�_=l�R=�E=�s�< �9�Dh1��՝��ὟI�>�'��8���>��;��-�|���`��q����f�L!μ@�;�   �   0���\B�<��<8��<01t<\ԏ�JA����������ɾ�h�W�B�^zy����Ӈ���*˿8�ݿ� �fu�꿈߿Z�̿1Ӵ�������z�YPC��~��Dɾ����o��h���H�3��e�<��=f$=d0�<���;P�漡m��Z����%���U�3����ޑ��R���ɡ��ڞ�ה������6`�7�1�Hn��L��P '��   �   lH��0C�8J<�!�<D��<@}��8�9�26޽I��-��m��j���L���{�H������a���+ ÿ��ƿ��ÿ�湿x?��|���!~�� N�-4��⟾��H�@+۽�D.�  Q8�ܿ<�]�<��<`+�8.�Y4��7e��S����Î��Ѵ˾���۶�����g��G��)о�ݲ��ӑ���_�3�͛ƽ�   �   �ͽ"�C��o%�(�D<�Ǔ<�+�;#��ۤ��Z)���k��������U��wuF��l�񯆿oᓿTu��o�������	��n$���o�FI���!������Ų�,�o����{���Ҭ��<���<ງ< i���&�����!�m�q�<^��)�Ӿ�� ��$��m%�Z0��4�1�B='�%�����پ�����5|��Y+��   �   ��&�ힺ�VS���.��[x<x�<�E��K�h鰽vK ��Pz�g,���.���2���M��b�)�p��u���q�
�d��FP�Y�5�<��H򾭾��}���k�&�5���L�@q.��]x<��<���XU�L�?P �Wz��0���1�a3���M�"�b���p���u��q�4�d��JP���5� ��M�m¶�V����   �   ɰo�̓�����4۬�H<���< ć<�*��T�&����R�!�v�q��Y����Ӿ�� �E!�j%��0��4�G	1��9'�܏�'���پ�����/|��T+���ͽt�C��W%�@�D<\Ǔ< �;`0��-���:-�
�k�����*��2���xF��l�����㓿�w��ᥟ�������&��po�;II�?�!�����Ȳ��   �   w䟾2�H��/۽�I.� I8<޿<�d�<Ĥ�< *�� ��+���_��S�[��މ��R�˾��㾚�󾢼���`��f羟$оٲ��ϑ��z_���ƽ��G�PC���J<%�<0��<P�����9��;޽D
I��0��J������L�<�{�R���X¨�̬���ÿ�ƿ�ÿB鹿�A��f���$~��N�[6�f��   �   Gɾ6�����������3� f�<$�=R$=�?�<`P�;x���d��q��X�%��U�󃀾=ڑ��M���ġ�*֞��Ҕ�~���//`���1�(i��D����&�0���xN�<T�<��<�*t< ݏ�E����������ɾxj�ӳB�c}y���؉��-˿��ݿ��w����߿r�̿մ�o�:�z�|RC�����   �   Y2�����:�ϵ�`����<��8=��_=*S=�M=Ĉ�<�9��W1��˝�܇�XC�l�'��8���>���:��x-�[��U��4��x�f� 	μ`Y;`��<J�=|
,=�	=�(<�i��Ž=A�����pX�,��f�!j��Ef����п��I� �|��H
���=>�����ѿ'󲿢����e�3O+��   �   D
��C���\���������<�-G=	Ȅ=fȌ=�؀=� K=̥�<�C	<H�}�:m��v��坽�V��2P��g���:��Y�����I���㼰���F�<n|=�A=2l[=.�N=~�=0�;<�7�m!����e�C������D�Q���Kv����ȿ:��߇�,��!��Qi�8��������3뿄�ȿ�����*�B��   �   h%�y&˾��w�E���12�u^<�N=���=���=4��=-��=�s=��1=l:�<`�<�$ݻ���H�j|��F����̼��u�@��\X<0&�<�32=rc=��=��=��d=�= �<9��c�T��eF��oAо	��\�W�%Ҏ�<c��	�ڿ&N����c�&%&��C)�KE&�Q��L(������ٿl��C���4`U��   �   �!���׾i���ҭ���K�x�6<8�Q=�L�=���=䥷=���=���=�W�=�L=�a=��< d^<P3�; �O; Wp;@<`�{<@I�<��=G=f�s=�#�=���=� �=0�p=&'= �O�(���""����&�ݾ��#�G,d�Ȣ��B콿��{=����
�%�)/��`2�/�$�%��q������ꅼ����� a��   �   :$��Cܾȥ������gT��8(<��R=�ʜ=V�=J@�=4f�=!��=��=�yl=��8=&�	=���<,F�<�n<�Cs<$��<���<�=T6=D}a=r��=�r�=���=��=zEt=��= ��l��^�΍��e⾁5'�lh��R��4���������=�a�(�k42�A�5��12�G�(�������|����$����)e��   �   !���׾���������K�0�6<��Q=iM�=���=��=Ɩ�=���=
X�=��L=b=��<Pd^<�3�; �O; Xp;�@< �{<�I�<�=RG=��s=$�=똓=T�=H�p=�(=`�O������ �<�����ݾ��#�3+d����n뽿���<���N�%�a/��_2��/�m�%�Hq������� ���-���a��   �   �#�K$˾��w�-��P,2�8�^<`�N=t��=v��=���=`��=>s=��1=�:�<��<�$ݻ䟞�0�L|�4F��|�̼`�u����^X<x'�<n42=�rc='�=t�=̠d=�= �@9��c�"���D��-?о|��P�W��Ў��a��(�ڿ�K����Bb��#&�9B)��C&����'������ٿ�j�����:^U��   �   B
��@����\�د���D��<1G=$Ʉ=$Ɍ=6ـ=XK=���<�D	<��}�"m��v��坽�V��"P��L���:��!���4�I�,�㼐���H�<�}=��A=Vn[= �N=��=��;�z7�U��X�e��?������D�����t��2�ȿ<��/��R��+��Qg�D�����d��1���ȿ����k�B��   �   c-�Z
����:�ȵ����!�<�8=Z�_=�S=�N=��<�}9��W1��˝�ԇ�TC�j�'��8���>���:��x-�<�hU�����j�f�xμ�r;\��<��=,=��	=ț(<�_�FŽ�7A�你�ZS�\,�df��g��+c��d�п$��� �2���E
�V
�<���C�ѿ�����e��K+��   �   �AɾQ���0��}�����3��s�<��=P$=<C�<PY�; �漋d��J��N�%�
�U�񃀾<ڑ��M���ġ�"֞�|Ҕ�j���/`�1��h��C��8�&���� T�<�&�<ę�<8It<8Ǐ�>=�������p�ɾ�f�+�B��wy�m��������(˿��ݿ2���r�5��*߿#�̿2Ѵ������z��MC�}��   �   ߟ�^�H��$۽h:.� s8d�<(n�<Ī�< a*���/+��t_���S�W��݉��S�˾��㾛�󾡼���`��\羍$оٲ��ϑ��z_����ƽ��G��C���J<0�<ĳ�<�C����9��0޽JI�6+���~�3���	L�Y�{�\���󽨿�����¿
�ƿ�ÿ�乿8=��r��~���M��1�.��   �   ��o�Z����������5<x�<�̇<�����&�g��-�!�`�q��Y����Ӿ�� �E!�j%��0��4�F	1��9'�ԏ�����پ����:/|��T+��ͽ��C��H%�X�D<t֓<`g�;���Z����%���k�����N�󾲉�KrF�Dl�߭��.ߓ��r�����N��X��C"���o��BI���!�I��������   �   Y|&�p��� @���-���x<���<�A�rI��谽>K ��Pz�],����.���2���M��b�*�p��u���q��d��FP�Q�5�2��H򾊾��Q�����&������H�`#.��yx<X��<�+��A��ⰽ�F ��Jz��(��?�쾬+���2��M�ƶb��~p���u��q���d��BP���5�&��C�{���1����   �   .�ͽ��C��+%��D<Tؓ<�W�;��ģ��)�t�k��������U��wuF��l�򯆿nᓿUu��p�������	��l$���o�FI���!������Ų�̫o�������ɬ�@+<L�<�Ӈ<@ߊ�R�&���<�!��q��U���Ӿ�� ���f%��0�4�t1��5'�s���ɳپ~���^(|�QO+��   �   �G���B�p�J<�5�<��<�X��D�9�M5޽�I��-��e��h���L���{�H������c���, ÿ��ƿ��ÿ�湿v?��y���!~�� N� 4����៾\�H�*۽A.� �e8��<�r�<,��<��)���#��/Z�f�S�V��*����˾	��o��O����Z��e�оԲ�bˑ��s_��n�ƽ�   �   0;���a�<�/�<���<�Gt< ͏�@��L�������ɾ�h�W�B�]zy�	���և���*˿9�ݿ� �gu�꿈߿X�̿.Ӵ�������z�PPC��~��DɾZ���������x�3��q�<0�=6$=`P�< ��;���M\�����%���U�����Ց�,I���Mў��͔�+���s'`�@�1�{c�J;����&��   �   `�<�=4,=:�	= �(<Pb��Ž�9A�~����U��	,�\f��h���d���п��-� �S���F
�{�0=����ѿ��m���$�e��M+�0�I����:��˵�P��D�<��8=�_=�	S=�U=d��<8L9�0H1���	}�<=�þ'��
8�J�>�~�:��q-��x�?J����P�f�\�ͼ`;�   �   &�A=r[=^�N=T�=	�;&}7�����e�EA������D�R���u��c�ȿ������7��"��Ph�A�����A���2�Y�ȿ���������B�+C
��B��3�\��ཬ��8�<F1G=ʄ=�ʌ=�ۀ=2K=(��<p	<�O}� ^���u��ܝ�*M��1F��u��1��p�����I��㼰���,[�<
�=�   �   ��=��=@�d=��= \@9N�c����^E��@о��&�W�eю�Ub����ڿ�L��[��b�f$&��B)��D&�����'������ٿik������c_U��$��%˾��w�d��6/2�0~^<6�N=쎒=���=��=���=�#s=��1=K�<`�<��ܻ܈������o��-���l̼�zu� `��X<6�<h:2=�wc=�   �   ՙ�=�=:�p=()=�O�����.!�l���E�ݾ$�#��+d�U����뽿{��$=�Z����%��/�E`2�/�Ѷ%��q����T�俟������� a��!�i�׾1��������K��6<&�Q=�M�=`��=Ȧ�=Ɨ�=���=�Y�=֊L=~f= ��<�y^< b�; P;@�p;PW<P�{<dS�<2�=�G=��s=J%�=�   �   �u�=�O�=D�X=���<��¼��ƽ,}P�I����I�/N�Fɍ�钹�ǒ�fw��\$�}�:��YM��Z�!�^���Y��3M��@:�?�#�\��5��p���9苿��J�P
�^)��aqF�O��8�e��=��=�M�=d��=�ʠ=峍=Hg=��,=@��<�v<Pg�;`!�@q���d���kL:@n<�<�|
=�@=B�q=���=�   �   ��=/w�=@T= ��<�#��z���6yK�­���
�]7J�)E��g��ۮ��
��!�#N7�n�I���U��>Z���U��xI��	7��� ��V	�&������{���G�m��������A�u����!T�TR=�8~=�&�=d�=���=v��=^�G=�W=�ڎ<�qZ; ��Г�����0���{B� R���)<�5�<<.!=HX=���=�   �   �Xi=�m=d�D=���<�-��m⯽�=�����m�E?�8����/���fٿ�Q��m���-���>�WJ�"N��4J�r�>���-�a<�G��',ؿͫ�y����q<���������~74�e7��@Q"��2=��l=�W�=щ=T�n=�B2=�:�<P�;0s����@���g��x��
p���P����γ��>\��8�<2�	=��D=�   �   4�=`�8=�(=賻<�r^�<���&��H����Ƶ-��
q�����ǿ����]�Dd.��q8�i<���8���.�����>�^���Mǿ�����9o���+�n��f����U�tφ�@��� =�M=(�_=oC=L\=��$<<���&4����B�Ľ�콴��W6	�I
�
W���yнf��>nV�D�μ ��9�V�<�   �   �#<̖�<|�<$�<P�n3n���3}���˾��}�S�p]���_��n�ֿ���(������N#�f}&�9�#�d� h��8��"�׿j���D4��_!S�	���|ɾd�w��K���T������u�<D�=�R=�%�<�0ֻP!��������j���C��`���s�${�$,v��We��SJ�v�'�� �ح��"�G��i���   �   �� `���Pw<"t< �J��P,��Pٽ��L��o������3�8�n��ڗ��ϸ��Fؿ�)��1�.|�1�L��A�����N�ٿ�	��雘��o��3�y#���5��סI��Gѽ�b���;0�<|w�<p��;웥��Or�#b۽�7%��_��r��	2���ͺ�WȾ�};۽ɾxs��/ҩ���h��.�;��䊽�   �   /��B:��Ļ ��; xɹ��ۼ7#��]���烾V�ʾ3���(C�Xz�.���鳿5�˿'Q޿*�꿬��p뿁�߿�vͿ ��������@|�V�D�"��Z3˾�Ճ�b�)ʗ���ü�4`;xl,<�v	���������kH�ZL��BS��Vsܾ�< �ў�@	�S������4�/\�~LΆY���-��Q���
��   �   �����T��� ����I�8rd��7F�-ٽ��A����v߾8]��<E�Lws�揣����E(��u������z��SL�����Йv� �G�+<���ᾕǚ�E~C���ڽx�D���O� �:P3���p�UG����	�_�Z�G>��δҾ&K�� �F�8��)L��X��]���Y�&N��Z;��J#�����׾z����
b��   �   �]�w�N{��H�Ѽ�u�� �����ż���B��HX�p(���ᾂC���8�a\���{��l��I��������3��՜����~��_���;�E��F"��n����\��s��v���Ѽ o�������ż���T���X�C,���ᾐF�x�8�Ne\�6�{�Go��厒�b���D6��L���F�~���_�T�;� ���&�Nr���   �   cʚ�*�C���ڽ
�D���O��F�:�	��4^�x@����	��Z�:����ҾH�7| �@�8�K%L���X�j{]�q�Y��N��V;�9G#��
���׾�����b��
�(������ �I�8�d�x?F�e3ٽ��A�! ���߾�_�@E�T{s�P�r������+��S��������}���N��4�����v�D�G��>�ѣ��   �   N6˾�׃��d�J͗��ü @`;(|,< �����>|��F��BdH�'H��2N��umܾ�9 �=����������b1��X��F��T���)���xQ��
�(���0�`mĻ`��; �ɹ��ۼ�'��Ƣ�tꃾЕʾ���r+C��z�J��=쳿ܘ˿ T޿"�꿫￺s�F�߿yͿb��������C|��D�$���   �   `&���7����I��Jѽze���;���<���<�>�;@���F?r��W۽r1%��_�#n���,��Ⱥ��QȾ�w;�ɾ�m��.ͩ�������h���.�k��)݊���  +�`aw<'t< �J��U,�8Uٽ"�L�<r������3�(�n��ܗ�Ҹ�VIؿ-,��y2��}��2����� ������ٿv��|�����o��3��   �   Z���~ɾ��w�!M�r�T� ��hy�<v�=VY=�8�<��ջL@!��ｴ����C�ڳ`�J�s�q{��#v��Oe�kLJ��'��� �����z|G� S���>#<���<4�<��<����8n��d6}�!�˾Ȱ���S��^��Ea��^�ֿ��g����VP#��~&���#�Le�Fi��:��Ӭ׿Җ��g5��%#S��   �   ��+����f���!W��І���>� =�M=�_=�uC=e=x�$<ܛ���4�����vĽ������^0	�q��K���oн[����^V���μ ��9�f�<�=9=��(=���< |^�m>��
�&�?J����:�-��q�Ğ�R�ǿ���x��^�xe.�;s8��<���8��.�����?����Oǿ����<;o��   �   �r<�����X���D84�(8��(R"��3=��l=&Y�=HӉ=�n=J2=\L�<pi�;��r������@�Ȼg� x�,�o��P� ��������[��H�<��	=��D=P\i=�m=L�D= ��<�1��^䯽�=�2����n�b?������0��
hٿyR��n���-���>�SJ�#N��5J�G�>�a�-��<�����,ؿ�ͫ�򐂿�   �   bG����ن����A������ T��R=�9~=Y'�=�	�=+��=L=��G=�\=��<��Z;Н�����̃��T����`B������)<�>�<2!=BX=���=R �=�w�=dT=���<�&������8zK������
�8J��E���g��z��P
���!��N7���I��U�>?Z��U�NyI�9
7��� ��V	�~��#��������   �   ]�J��O
� )��qF��
���e�X =��=+N�=���=�ʠ=��=^Hg=�,=���<�v< i�;�� � q�� e�� iL:�m<��<`|
=��@=��q=���=gu�=�O�=��X=X��<X�¼/�ƽ�}P�����J�bN�dɍ�
�����ww��\$���:��YM��Z�#�^���Y��3M��@:�/�#�L����S���苿�   �   rG���ㅫ�w�A�㥭��T�zT=�:~=�'�=�	�=E��=[=ԣG=�\=��<��Z;�����������<���x`B����h�)< ?�<F2!=�X=��=� �=x�=�T=0��<�!�������xK������
�7J��D���f��~�俸
�Έ!��M7� �I�s�U�+>Z��U�_xI�j	7�J� �0V	����`�������   �   �p<����������54��4���@"�v6=��l=�Y�=�Ӊ=x�n=jJ2=�L�<�i�; �r������@�Ȼg�x��o�ЊP����춳�@�[��I�<D�	=l�D=\]i=l!m=p�D=\��<4(���௽�=�P���Xm��?����.��,fٿZQ�Um�.�-�¦>�hJ�!N��3J���>���-��;����#+ؿ?̫�ȏ���   �   3�+�R��ߒ���S�̆��׷�4� =p�M=��_=�vC=�e= �$<l����4�����vĽ������\0	�j��K���oн.���F^V�4�μ *�9�h�<p�=,9=��(=l��<�a^��9��x�&��G��S�뾬�-�*	q�������ǿ�����\�%c.��p8�"<�y�8���.�����=�Ć�Lǿv����7o��   �   c��Gzɾ��w�I�v�T� ����<��=F[=�:�< �ջ�?!��흽�ｴ����C�޳`�M�s�p{��#v��Oe�WLJ�Ա'�b� �A����{G�lP���E#<���<x!�<���<�h�-n���20}���˾�����S�F\��0^����ֿ��� ��t���M#��{&�ν#��b��f��6��>�׿͓���2��<S��   �   ���3���I�BѽxY��;<�<|��<@O�;�����>r�lW۽b1%�
�_�"n���,��Ⱥ��QȾ�w;�ɾ�m��!ͩ�q���^�h�x�.����q܊�$�� ���qw<8>t<�oJ�$I,�Lٽw�L�|m������ 3���n�hٗ�θ��Dؿ'���/��z��/�������|�����ٿ���(���,�o�K3��   �   �/˾�҃�(^�>ė���ü��`;��,< ��|�漞{����+dH�"H��2N��wmܾ�9 �>����������_1��X��F��T���)���xQ���
�'���-�PMĻ��; �Ź`�ۼ<�����僾C�ʾ%���%C�z�<���糿��˿jN޿B�꿲��m뿩�߿�sͿ���������<|�i�D�Ҍ��   �   AĚ�IyC�+�ڽ��D�ȟO��@�: ᐻ�W�y?����	���Z�:����Ҿ	H�:| �B�8�L%L���X�k{]�q�Y��N��V;�1G#��
���׾{���Pb�
��}��@������ wG�HPd��-F��&ٽ��A�����߾�Z��9E��ss��쏿x���O��z%�������(x���I������Õv���G�c9�����   �   ��\�o��o���pѼ�������|�ż~�����X�a(���ᾂC���8�!a\���{��l��J��������3��Ԝ����~��_���;�:��)"澶n���\�s�+u���|Ѽ�1��0���p�ż�y��F���X��$����ᾪ@�h�8�#]\��{�Xj���������1��R����~���_�0�;�-��D��j���   �   U�-w����������%G�8Yd��3F��+ٽ��A����h߾5]��<E�Nws�菣����F(��u������z��QL�� ���șv��G�<�۟�jǚ��}C�*�ڽ��D���O� L�:��H�s9��*�	��Z�56����ҾE��x �]�8�!L��X��v]���Y�~N��R;��C#����׾U�����a��   �   k��(#��Ļ  �; uŹ0�ۼ�!������烾E�ʾ/��(C�Xz�.���鳿7�˿)Q޿*�꿭��p뿀�߿�vͿ��������@|�L�D���83˾QՃ�ja�Hȗ���ü`�`;@�,< F��漌t��H���]H�-D��dI���gܾ_6 ���������+���-��U��@ᾺO���%���qQ���
��   �   ��  5`�w< Ht<�tJ�nL,�kOٽB�L��o������3�9�n��ڗ��ϸ��Fؿ�)��1�/|�1�L��A�����L�ٿ�	��囘��o��3�^#��x5��Z�I�8Fѽ
^��
;p�<p��<`��;�j��z/r��M۽=+%���_��i���'���º��KȾ�q;<�ɾhh�� ȩ�㲐���h���.�c��WԊ��   �   j#<t��<P)�<��<�k�80n�l��2}���˾��}�S�p]���_��n�ֿ���)������N#�g}&�9�#�d�!h��8�� �׿h���B4��X!S�����|ɾ
�w�K�"�T�@V��x��<��=�`=�K�<`mջ81!��䝽���B��A�C��`�۱s��{�v��Ge��DJ��'��� ������kG�,8���   �   �=�	9=p�(=���<�d^��:����&��H����ŵ-��
q�����ǿ����]�Fd.��q8�i<���8���.�����>�^���Mǿ�����9o���+�Z��G����U�;Ά��添V� =n�M=t�_=�|C=�m=H�$<����~�3�����lĽ������j*	�����@��*eн�NV��μ ��9Tz�<�   �   �ai=l$m=R�D=���<�(���᯽�=������m�E?�8����/���fٿ�Q��m���-���>�YJ�	"N��4J�r�>���-�`<�G��&,ؿͫ�w����q<���������?74��6���G"�86=��l=�Z�=sՉ=��n=�P2=�\�< ��;X�r�`��u@�d�g�J�w�j�o��|P����������Z��Z�<h�	=�D=�   �   �!�=�x�=�T=���<�!��"���yK������
�[7J�*E��g��ڮ��
��!�#N7�o�I���U��>Z���U��xI��	7��� ��V	�&��ߍ��z���G�j������i�A�����T��S=,;~=)(�=�
�=l��=�À=��G=Xa=�<�6[;���w���u��,����EB����@*<I�<�6!=(X=t��=�   �   ���="az=��5=�L5<�y5�_h�́���ھF�(�v�s�u��R�ؿo���#��A��E]�$�u�� �������\u��\��6@�C�"�
8�\Nֿ@d���Mp���%�?�վ
E{�����B����<�P=�̊=�:�=o�=fl=j�1=���<�j:<��C�ؙm�j����μ ����Ì� �޻��;���<8�=��Q=�{=�   �   �D|=�o=��/=�H4<6�/�@
���}��a־��%��co�㒣�y�ԿV+� !�ϔ=���X�=�p�\]���F��;c��2yp��X��<��( �����ҿৡ��l��"�Z�Ѿ�u�ۙ�B����<ށJ=��=���=��=��N=�k=85�<�o&��N��̱�$�:�&����@�(��P����:<\�<\t4=��d=�   �   �ZH=aL=�z=��-<��1��*m�Cuɾ�B���b�1���lʿ
@��*
�.�3���L�jb��2q��v��mq�Q�b���L�.Y3��}�\����ȿF����_�����\ž��e�rs�.c����<j'7=@�f=��b=�%9=���<pj�;��y��K�H�l�~c���)��F����H���Y��`�}�T�.�L��� _�: [�<��=�   �   l��<V�=���<��<T&�!�ѽ�mS��k������N�	���繿���ߧ�̎$���:�{�M��iZ�� _��Z��CN��m;���$�b��z[�������/�L�[��Q"���WM��Ž��༈�s<�c=f�(=�=@^{< � �a"��|����ҽ���d7,��
2�F�-�Sj �گ
�j�ݽ(ޞ�vz<��g��8<�   �   P���(�U<�3�<P�;|ۼ��R|3��B�����$5���z�+ؤ��3Ͽ�d���*��O%��5�ƻ?��C�OK@�C�5��>&�����6���qϿ����`�y���3�e.��H百O�.�=��������1<\��<��< �:���\5��)9ὴ��s�M�[kw��O���3��OR���@���H��p�|�`;T�2�&�f�@Օ�t���   �   ��L�PÎ� �X� �!��F�����!j�qG���?;�V���T�⌿N�� �׿���g!�O5���#��('��~$�<3�u<�����!ٿ�ٲ��A���T����̾�}��7�*~���F���ui;��;�7I�� 5�%����"�FT�Z&���Y��.˾��W��n��N��~t�Hsξ���a��N\��>���ý�   �   �ݽ~zk�G˼`�9��q��.lJ�ދڽ|G��Ѣ�{8��7,-�vg�(L���n��,ҿG?�Pl�*���*� 	� ]��q�/-Կ���|����h�_�-�<���ʾ��^oF�~!׽rhA��;���L�D���8�X�yҽ�C,�TS}�C(���۾�;�/�ٴ*�b�5���9��e6��F,�C&�$��(o�dd��~i���2��   �   9�}?ݽAh�t�ݼt柼����B���.�3-t����ڝ�6���i����������d��ѿ��ܿ���ݿG�ҿZ��s窿�8����l�M�7�)��z?��j�u�y��G��������@�˼�B\�g{ս�!4���������6��` ���?��[�
�q��%��fՂ�#�����s��1^��VB�Y�"�a��c�ľ�6���   �   ���E-���Ľ��E��)ɼ�dƼ�bA�x���Z]*��c���ƾ^d�)b1�Y�[�PI��7Z�������竿/[������r����3���!�^���3�9b
�isɾ�|���@-���Ľ*�E��'ɼ�jƼjA�� ��b*��f��Q�ƾ;g��e1���[��K���\�������꫿4^������F�3������� �^��3��d
�qwɾ�   �   �B����u�l�������� ����˼08\��sս4�1�������0���
 ���?�b�[��q��"���҂�������s�-^��RB��"������ľp3��9��8ݽ�8h�H�ݼ�柼��aG��j2��2t��Ļ�[��D6���i�ً��H����g��?"ѿ�ܿZ��+�ݿY�ҿ�\���骿�:��W�l�6�7�e���   �   ����4����rF�&%׽rkA�l:��;�����z�X�xҽ�=,�~K}�`#��5�۾88�]���*��5�!�9��a6��B,��"���~i྽_���e��q�2��
ݽnok��9˼`�9� t��NqJ�͐ڽ�G�hԢ��<���.-�}yg�7N��q���ҿSB��m����,��	��^��t��/ԿY���~����h���-��   �   M�F ̾D�}��9�����F����i;�4�;�I��5��������wT��!��]T��$(˾Y�⾑���g�����n�pmξ������\�G9�>�ýހL�0��� �S� \!��J��䌈��l�xI���B;�X�9�T��㌿X����׿�����"��6���#��*'���$��4��=�W���3#ٿU۲�IC��^�T��   �   V�3��0���虾�.�􏤽� ����1<���<��< �:4q�M,���-������M��bw��J���.��AM���;���C����|��3T���&����̕�p���`��p�U<�:�<�!�;8ۼ���~3��D�����5�>�z��٤��5Ͽg��=,�[Q%�Y5���?���C�M@���5�@&�����8��sϿ󫤿o�y��   �   j�L�:��|#��*YM���Ž��@�s<�f=��(=,=P�{<�t �HQ"�hs��Ԅҽ�	����0,��2�z�-��c ��
��ݽ2՞��k<��O���3<���<��= ��<(�<�(�׃ѽ�oS��m��/��7�N���鹿F��ר��$��:� �M��kZ��"_���Z�FEN�0o;���$�0���\��	��Q���   �   ��_�+���]ž��e�Ut�~c�x��<�)7=��f=��b=,9=���<@��;��y�>�<�l�a[��#!������a@��R���z}�N�.�脫� ��:j�<V�=�^H=�cL=�{=�-<Z��g���m��vɾ�C�͐b��1���mʿCA���
��3���L�8kb��3q�S�v�oq�c�b�~�L��Y3�H~�A�����ȿҬ���   �   �l�<�"���ѾJ�u�
��fB�$��<4�J=��=ɪ�=4�=�N=�p=�@�< �$�@������&������@���@ͱ��:<�d�<�w4=J�d=|F|=�o=��/=�E4<�/� ���}�|b־3�%��do�a����Կ�+�� !�T�=���X��p��]���F���c���yp�\�X�m�<�!) ����ҿ����   �   �Mp���%���վ�D{�<���^��,�<v�P=͊=5;�=9o�=�l=ʀ1=0��<l:<@�C�ؘm��i����μ@����Ì�0�޻е�;���<�=��Q=��{=���=�`z=�5=�I5<�z5��h�Ḱ��ھv�(���s�/u��x�ؿ&o��#��A�F]�5�u�� �����
��
\u���\��6@�0�"��7�8Nֿd���   �   �l�q�"���Ѿ��u����?����<F�J=��=��=j�=F�N=�p=�@�< �$�,@�������&���������̱�`:<0e�<x4=��d=�F|=�o=�/=(M4<"�/��	�a�}�Ua־b�%�xco�����(�Կ!+��!�r�=���X���p�]��'F���b���xp�S�X���<�t( �8�%�ҿh����   �   ��_�����[ž��e��p὆^��<�+7=�f=��b=�,9=x��<0��;p�y�>�J�l�d[��-!������^@���Q���z}��.�L���@��: k�<�=�_H=@eL=�}=Х-<��t���m�ltɾ[B���b��0��>lʿ?���	�q�3���L��hb�r1q���v��lq�%�b���L�TX3�}�1���&�ȿ}����   �   ��L�#��� ��1UM�A�ŽL� �s<�i=��(=J= �{<ps �Q"�as��΄ҽ�	����0,��2�x�-��c ��
�ͪݽ ՞�k<�|N���7<���<��=X��<`�<�!�[~ѽ�kS��j����F�N�0���湿M����ȍ$���:��M�PhZ�F_�~�Z�^BN��l;���$�s���Y迢��t���   �   ��3��+��9噾P�.�����4����1<|��<�!�<��:�o�,���-������M��bw��J���.��DM���;���C����|��3T���&�c�R̕�:���R����U<PB�<�O�;�ۼ�����y3�DA��ƃ���5���z��֤�/2Ͽ�b���)�{N%�5��?��C��I@���5�3=&�����4���oϿ�����y��   �   ���̾��}��4�
y���4�� j;PR�;�I��5�Z������wT��!��_T��&(˾]�⾕���g�����n�gmξ�������\�
9���ý�~L����� �O�����7��Ѕ��vg��E��O=;U�:�T�����}�����׿������3�)�#��&'�}$��1��:�����ٿ�ײ�*@��p�T��   �   '���û���jF��׽�]A�(��0#�,���*�X��ҽ�=,�fK}�\#��5�۾:8�`���*��5�"�9��a6��B,�"���niྦ_���e���2��	ݽ�lk�H1˼�h9��`���bJ�8�ڽVxG��΢��4���)-�sg�JJ��ul���ҿc<�j�z��)�g	�z[��n�o*Կ����z����h���-��   �   �;����u�5������`����,�˼�4\�vrս�4��������0���
 ���?�e�[��q��"���҂�������s�-^��RB�۷"�{����ľI3���9�M7ݽ�4h��ݼԟ�d��O=��"+�/(t��������&6� �i�b���+��a��ѿ��ܿ��࿮�ݿ$�ҿ*W���䪿P6��ȇl��7�����   �   Ky���;-���Ľ��E��ɼpTƼ|]A������\*�oc��сƾ[d�)b1�[�[�RI��9Z�������竿0[������s����2����^���3�,b
�Hsɾ�|��^@-�ڻĽ��E��ɼ�QƼ�WA������X*�{`���}ƾ�a��^1�g�[�G���W������嫿.X�������죿����������^�7�3�R_
��nɾ�   �   *9��/ݽX*h�ܽݼџ�����@��&.��,t����՝�6���i����������d�� ѿ«ܿ���ݿF�ҿZ��q窿�8����l�B�7���R?���u����ڵ��,����x�˼�+\�}kս�4����R���+��X ���?��[�(�q�i ��Ђ�므���s�m(^��NB�;�"�v����ľ�/���   �   � ݽ`k�!˼@X9��_��DfJ��ڽ�{G�_Ѣ�k8��4,-�vg�)L���n��0ҿJ?�Ql�,���*� 	� ]��q�--Կ���|����h�T�-���������nF�x׽LbA��)��8�`�����X��ҽ�7,�D}������۾�4�����*�Ƃ5���9�<]6��>,���]|��c྾Z���a���2��   �   qL���� �I� �P8������ji�=G���?;�V���T�⌿P��"�׿���i!�Q5���#��('��~$�=3�t<�����!ٿ�ٲ��A���T����̾��}�7��{���7��@!j;@{�;��H��5�������pT�v��HO��a"˾�����`�����g�ogξC��Y��R
\��2�+�ý�   �   p��� �U<dK�<P_�;Tۼ\ ���{3��B�����#5���z�+ؤ��3Ͽ�d���*��O%��5�ƻ?��C�OK@�C�5��>&�����6���qϿ����\�y���3�J.��百��.�`���h����1<���<�.�<�D	:�U뼦#��L#ὔ��0�M�#Zw�(F���)��:H���6��-?���|��+T��~&�*�EÕ����   �   ���<�=���<��<P"��ѽ,mS��k������N�
���繿�����̎$���:�~�M��iZ�� _��Z��CN��m;���$�b��y[����~��*�L�R��3"��TWM���Ž̃༐�s<�k=��(=�=p�{<PD �dB"��j��{zҽ�5��),���1���-�T] �ޣ
��ݽ�˞�`[<��4���_<�   �   �dH=�hL=$�=H�-<|��j���m�8uɾ�B���b�1���lʿ
@��)
�.�3���L�jb��2q�	�v��mq�Q�b���L�.Y3��}�\����ȿE����_�����\žb�e��rὊ`�@��<�,7=��f=��b=B29=,��<��;X�y�@1�Ƭl��S�����+����7���I���k}���.��l�� Ӳ:�{�<��=�   �   �I|=�o=l�/=0P4<�/�
���}��a־��%��co�䒣�x�ԿV+� !�ϔ=���X�=�p�]]���F��;c��1yp��X��<��( �����ҿৡ��l��"�R�Ѿ��u�y��PA�l��<��J=k�=뫋=�=��N=@u=4K�<�F#��2��H�� ���&��������奼 ����3:<o�<4|4=��d=�   �   gs=Rd^=��=�rȺ�����"�T%��İ��׾A�&؊�.�����������+:�4W]�u&��Ef���ޙ�\����ٙ��F��G���U\�g�8������p��(��Z?�Oo������#��p���@;:H#=�o=�=�=�%q=B=�=f<@Ya��ߜ����`m#��r0���'�2�	�4���P�ڻ8l*<�;�<�U1=�/`=�   �   �`=��Q=�2= BԺ}���䕾����!>�b��pM���s�c_���6�Y�@�z�u>���h��S��>o���3��"�z�?X���5��6��?�Lb��3̆��;�������������i�`v6;��=��b=��q=L�W= a!=X#�<`c;�쉼
��@?D�:Di�B~w��m��QL����`�� ��h��<0�=��F=�   �   У&=��*=�>�<���8k��L������"��3�;������t�俛���X-���L� �k��`�����c���ʌ�و���k���L�:�,��$���wx��!���w1�ۏ澲���'3���X�@�;�f=��;=p�7=�c	=Pu<��,��j�n�lڤ�k8ɽo�L�mg㽡�ͽ���LD}�,-��K�ȯ/<�E�<�   �    _�<�c�<H�<`�w��Q����E3|���ӾI#��l�3d���9ҿCr�f����:�&�U�?�l�\�|�HN���;}���m��gV�9?;����$�Vѿ�l��J=j��!���оQ?w�'��֤@� ��8��<<��<PJ�< ��9x⼚5y�/pŽu�.�&��)@���P�R/W�aTR���B��'*���
�ܐν�酽x]� y���   �   ���  : D�;`����4�_J�@WX��J�������O�-Ŏ��ʺ��	�fT�`%���;���N�I�[���`�HU\��O�x�<��(&�%���I�p����Z���N�����F����T��%ٽ��&�P�����<���;@*����G��R������C���w��-���ƥ��뱾�l���Ѳ�tq��Di����|��JI��Q��FĽF�Y��   �   NM��2�	���l�P�u�t�A���z1�JΗ�����j/��5s��#���|ɿ����/�� ���/�>$:�	�=���:�} 1�k�!�v8����`Yʿ<����Ls��/�w������x.��C��f]��F�@x8� ���چ��=7�Մ����xY˾������������������V�ξ[6���҂�ъ<�=����   �   Bx
����},��޼�]�zI���	�rno�s���b�U�F�����S��M˿�W�����"�c7��>�3���#�3�\}�v�̿ɂ���Ԅ�$�G�H�8��n��R��d	�A˼�=!��;��L�\R�rÖ�J ʾF���<.���1��.D�dDP�#�T��Q��E�r|3�)=������;�ڙ��(W��   �   ��^���
���t�7�\���\�7eʽ
u2�� ��U۾����P�����t,��^x���pؿ5쿄������������qڿm���դ��ˆ��R�����ܾBȑ�L�2���ɽ��Y��&�Zx1��U������Z��a��&�ᾶ���b8�`�[�({�]剿�푿㔿�z���⊿��}�6Q^�L�:�^��k��b���   �   2���Q����� ��V�-�z�,�Gm��Z���O;O�U��[��Q��)�K��H{��i�������_��t�¿<wƿ�fÿ
���A"�����N:~�V5N�����:������Q����������-���,�_q��_����@O��X��[�羉���K�pM{��l�������b��Ƭ¿�zƿ@jÿ/���&%��Q���>~�9N����w?��   �   ��ܾ�ʑ���2���ɽt�Y��$��q1�P��[����Z��]�����R���^8���[���z��≿�ꑿ����w��/����}��L^�j�:�'��P����Q�^���
������7�T��|�\� jʽy2��#��@Y۾¤�Z Q�㉅�/��L{��/tؿ�8�.��^���_������tڿ�o��?ؤ��͆�K�R����   �   �I��ﾾ��n��T�k�Hc	�\7˼\4!��4��G��R�����ʾ����c*�T�1�*D��?P�6�T�Q�Q�E�;x3�k9����s�;s֙�b"W��s
�s���u,�l޼�^�RL��ܪ	��ro�� ����P�F�h��GV���˿�Z���k$�_9��@�*���%���B����̿܄���ք�ūG��   �   h /�,��l���{.��E���]� �E�(\8������҆�3�6�P|���~S˾��Q��ق��� �i��5�ﾁ�ξf1��u΂�a�<�i���)F����	�x�l�P�u�4v�p���\1��З���<m/��8s��%��ɿ;��k1�ҷ ���/�^&:�3�=���:�g1��!��9���b[ʿބ��UOs��   �   ��N�ڊ�mH����T��'ٽ(�&�����h�<�̍;����~G��H��^�N�C���w� )��"���O汾"g��"̲�(l��ld��Y�|��CI��K�=Ľ��Y�`祿 �:�b�;���4�4��M�ZX��L��,����O��Ǝ��̺��꿪U��a%���;���N�y�[�Ȋ`�jW\���O��<�Z*&�B���K�㞺��[���   �   �>j� �!��о�@w������@� x�8(��<	�< [�< G�9���$y��eŽ�n�h�&�?"@�.�P��'W��LR�c�B�� *���
�ɆνGᅽ*P� '���m�<�m�<�< �w��Q����5|���ӾnJ#��l�ge��f;ҿ-s�����:���U�!�l�g�|�RO���=}�Q�m�,iV�g@;�����$�DWѿ�m���   �   ��mx1����9����3�*�X���;fi=��;=�7=�j	=�5u<�x� ��Nrn��Ѥ�L/ɽ��ཧ�^㽨�ͽ�����5}�� �`�J� �/<�R�<j�&=�+=<A�< (�.;k��M�����6$�1�3��;���������M���Y-���L�M�k��a��ߨ��4��oˌ�������k�եL��,�X%�~�y���   �   ă�*�;������������i� �6;�=�b=��q=��W=�e!=L.�<`�; މ�ؿ�v6D�;i�uw�
m�XIL�������X��,��<
�=��F="�`=�Q=3= XԺ��}���\啾���B">��b���M��Lt��_�H�6��Y��z��>��#i������o��4����z��?X�C�5��6�P@b���   �   �'��&?��n���������p�@A;�H#=V�o=�=�=:&q=dB=J�=0f< Ua� ߜ�p��<m#��r0���'�:�	�x�����ڻXk*<`;�<bU1=�/`=�fs=�c^=�=@�Ⱥo��
�"��%������A�F؊�T����������+:�MW]��&��Of��ߙ�]����ٙ��F��2���U\�O�8������_p���   �   �ˆ�F�;�Ö��E�������i� �6;H�=��b=�q=@�W=�e!=�.�<��;$މ���z6D�;i�uw�m�`IL���|�� U��|��<N�=�F=��`=��Q=H4=�Ժ��}���|䕾ƪ��V!>��a��.M��Gs�%_�q�6��Y���z�>��Dh������n��C3��f�z�z>X�x�5� 6�V?��a���   �   ����v1�W�澛����1���X�`;�k=��;=­7=Tk	=�6u<�w� ��Xrn�Ҥ�P/ɽ��཮��]㽩�ͽ�����5}�f ���J���/<T�<~�&=.+=F�<���r5k��K������!�q�3��:��1��������X-���L���k�=`��K�������Ɍ����<�k��L�g�,�+$��㿗w���   �   w;j���!�ƾоw<w�����@� T�8`��<��<|]�< ��90���#y��eŽ�n�l�&�H"@�7�P��'W��LR�a�B�� *���
���νᅽ�O�����p�<�q�<��<��w���P���31|�1�ӾH#�bl�Cc���8ҿ�q�r����:���U�|�l�b�|�?M���9}���m�fV��=;����5#��Tѿsk���   �   ˑN�	��{D��d�T�� ٽ��&��y��P�<Pߍ;���~G�wH��Q�M�C� �w�)��)���V汾(g��&̲�)l��hd��I�|�nCI��K��<Ľ��Y��뤼 m:0��;������4�dFརTX��H��L��˘O�Ď�wɺ���FS��^%��;���N�+�[�X�`�S\��O���<��'&�����G꿼���|Y���   �   8/���,���Su.�A>���S�h�E��K8�����҆��2�6�D|��񥾂S˾��T��܂����j��1��z�ξY1��c΂�*�<�����:E����	���l�(�u��k�����~�0�@̗�ӿ��h/�Z3s�"���zɿ!��n.�_� ���/�,":���=�i�:���0���!��6���$Wʿd����Is��   �   �E��龾$�n�0O��鋽"Y	�T*˼B0!�x3���F�\R������ʾ����f*�X�1�*D��?P�9�T�Q�R�E�8x3�h9����a�;X֙�"W�6s
���q,��޼TT�oD����	�>jo�����b���F�����Q���˿�T�^��� �s5��<�:���!�y�Jz���̿�����҄�'�G��   �   ��ܾő���2�}�ɽ��Y����k1�*N�����N�Z��]�����P���^8���[���z��≿�ꑿ����w��/����}��L^�c�:���9��Z���^�D�
�统�F�7�L��j�\��^ʽ�p2����4Q۾h����P�����*���u���mؿ�1������������^nڿj��>Ӥ�yɆ�m�R�����   �   �����Q�J�������ֶ-���,�wj�������:O��T��K��N��)�K��H{��i�������_��v�¿?wƿ�fÿ���A"�����I:~�N5N�����:꾰���Q�.�������޹-��,�Jg������.6O��Q�����Z��y�K�TD{�Og�������\��0�¿�sƿ�cÿج��D�����5~�U1N�P���5��   �   ��^���
�1�����7����,�\��bʽOt2�z ���T۾����P�����v,��`x���pؿ5쿈������������qڿm���դ��ˆ���R����ɣܾȑ���2�=�ɽ�Y����f1�GI�������Z��Y���}�#���Z8�?�[���z��߉�葿ݔ��t��`݊�pz}��G^�O�:�������#����   �   /n
����� h,�p�ݼ�S�EF���	��mo�J���Z�P�F�����S��N˿�W����"�e7��>�4���#�2�[}�t�̿ł���Ԅ��G��G��p�n��Q�^싽Z	��#˼�(!�7-��B��Q�ݺ���ʾV����&�,�1��%D��:P�O�T�1	Q���E��s3��5�:��ղ;�љ�AW��   �   b=����	� �l�8�u�&l������ 1�Η�����j/��5s��#���|ɿ����/�� ���/�A$:��=���:�} 1�j�!�v8����]Yʿ:����Ls�v/�R��c��� x.�DA��`U���E�X58������ʆ��(�<�6�9t��쥾�M˾�������:��/����t��x�ξ/,��ʂ�M}<�3����   �   lԤ� }:���;������4�qHཫVX��J�������O�.Ŏ��ʺ��	�gT�`%���;���N�L�[���`�JU\��O�w�<��(&�$���I�o����Z���N�����F�� �T��#ٽb�&�ps�� �<�;�����oG�?��a��C���w�:$��뻥��౾xa���Ʋ��f��u_��|�|��;I�WE��2Ľ��Y��   �   ���<�}�<���< �w���P�����2|���ӾI#��l�5d���9ҿDr�g����:�'�U�A�l�\�|�HN���;}���m��gV�8?;����$�Vѿ�l��F=j���!���о�>w������@� t�8P��<��<0l�< ��9���py��[Ž+i��~&�@���P��W�ER�	�B�*���
�'|νG؅�:A� ���   �   �&=+=�J�<`���5k�L������"��3�;������s�俜���X-���L��k��`�����c���ʌ�و���k���L�:�,��$���wx�����w1�ˏ澑����2���X��;�l=��;=P�7=�q	=�Wu< O�����cn��ɤ�w&ɽ����齂T㽔�ͽE���t&}�>���J�@�/<lb�<�   �   z�`=��Q=�5=��Ӻf�}����䕾����!>�b��qM���s�c_���6�Y�@�z�u>���h��S��>o���3��!�z�?X���5��6��?�Kb��2̆��;�����啒�d����i���6;��=��b=
�q=�W=�i!=8�<@';�Љ�B��:.D�L2i�lw�
vm��@L��������@���|��<��=��F=�   �   ��\=,F=���<��D��b��*�;��=�����U������Kοw����'��^M��v����������-���w��&(��*ݡ�~����u�z3L�ae&�H����̿;����S��]� �����7��������T��<(�P=6Wg=��R=�=\��<�oT;/~��j�: ;� �^���k��a��k@�����s�� }k:�D�<��=h(H=�   �   {H=&�8=v�<ȥF��۞�Į7�����iQ
�.R��ݕ���ʿ]f���$�ŋI�Nuq��Ό��I��W,���b���2���>��J����p�ɌH��#��l�y.ɿ\���\�O�����0��0�3��(���s��W�<xC=��R=�
7=$U�<ȁ=<�l� >��vG�����]��o���8ٖ������N�|$�xA�x�<�8�<�,=�   �   ��	=��=�ҫ<�CP�����K�+�����h���F�~#��F��������o�z�>�.Gc�K��'ד�pȞ�����C���������c��&>�i������z��H��*�D��� �@���P(�B����P#��<�=$�=�/�< +�;�R��ֶE�������ʽ����Hr
�Ԝ��=���=ϽoΞ���P���¼�M�:�_�<�   �   P��;h]�<I6<�$n��ن��<��ʎ�`G쾢�4��	�������G��My.�3gN���m�~�����!\���%���؄��Wn�D�N��o.����d4�~4��dE���3���1U�mD���D��^<��<8E <�A�@�,�0.��CJｂu�DHA�1]�|o���u��#p���^���C�:�!�߳��=���n�8�@@o��   �   ����!��p��Ч���No�����v��n;�d��:e��ꜿޟ̿y �D��d�5�6�O�߉e�Y�t�Vz��Nu�2f��|P�f~6�^,�6 �/y̿_���bd�Ћ���˾h�s�q1��e��!��@l�@g�4��B��
x�6(�:�a��+�����ú���Ǿ�̾n�Ⱦ
���@�� ����e���+��n������   �   3���f@��ּ̇ۼ�3V�//ܽ5�K�
�����IB����]Я��ܿbK�]��@�0�H�A��M��Q��N���B�?�1������jݿ�"��N��tB�f��	2����I��tؽڧN��˼L$żw6��-�������S�x���WK��� �VY���eR�!�����7���}�1��jʽ��ғ�O�W�$m��   �   �\!���Ľ�f���#�fuI������� �8��$־��� \��}������ҁ޿������( ��%)�4|,��)��!�������߿߲�� ����\�Z)��־ʇ�>���S��ZD����"�^��̿�;]�"6q�������⾋��-r+���D�Y��!f���j�8�f�LZ�:xF��-�4t�$��1��Qu��   �   �R}���!�$wý��s���N� $������M�M���T����,��g����<����ѿ �?�D�a�
�ɱ��������ӿ(���)��4�h���-�K`��Z���"N��N�r'����K�t3o�h\�����vWz��K��vn��z�$�MiL���r�zb���ŗ��k�����{㠿�����n���t��mN�O&�<!��"U���   �   �H���So�$v� |��x�i���h�_��fh���m�紾e}�wG/�f�a�����9@��� ���!ʿ�6տEBٿ��տ�D˿�c�������̋�v�c�$�0�����D���No��r��x����i�f�h��c��4l�D�m�"봾 ���J/���a�4���!C����%ʿy:տ�EٿR�տ$H˿g��X���ϋ��c�c�0����   �   [d��/����N��R��(��x�K��,o� V��¾��Pz�JG��~h��Ɩ$��dL�m�r��_�����h��苣�W࠿����4l��(�t��iN��K&�����P��`L}�q�!��qý��s���N�z&�������M�����Y����,��g�����>����ѿ��A�F�i�
�Ƴ����^����ӿǪ��5+��h�I�-��   �   {+��־�ˇ�����U���D����&�^�>ſ��W��.q�˧��z������m+�.�D��Y�Ff�+�j���f�GZ��sF��-��p�f�徥��i�t��W!�څĽ�f�V�#��vI�ΰ���� �����'־ ��U\���������޿0������* ��')�x~,�H�)��!�������F� ������p�\��   �   �B���4��R�I��vؽ�N�ܢ˼0żk6�d%����(�S�Ѐ���E���侪U�$��:N���e��H��\z�Ҟ��Ľ�ZΓ�E�W��g�p���P\@���ּ�ۼ�5V��2ܽX�K������sLB����dү���ܿ�L���B�0���A��M���Q��N��B�&�1�0��n��?lݿ�$������   �   �cd�)����˾��s��2���e�$��@��򻨘� :���l�X(���a�'��Z�������z�Ǿի̾Q�Ⱦ<	���;��R����e�2�+�bd�~����!� O��T����Qo�j�� �v�Cq;vf��<e�K윿��̿� �����5�B�O�<�e��t��Xz�Qu�s�f��~P��6��-�4  ��z̿�����   �   $F���3�B�@��D��آD���^<��<hi <��@�҂,��$���>��n��@A�$�\�
o��u�ep���^���C��y!����,�����8��o����;�g�<xS6<�$n�;ۆ�J>�&̎�{I�#�4��
��������G���z.��hN���m�8��#��[]���&���ل��Yn���N��p.�T���5�~5���   �   �����D�E ��@���Q(�|��� L#�D�<�=�=T?�<�y�;�:����E�E���q�ʽ����m
�����3���4Ͻxƞ��P�4�¼�o�:�m�<��	=��=�ի<�EP�%�����+�π��yi��F�C$��A�������p�t�>�nHc���
ؓ�cɞ�����)����������!c�W'>�������V{���   �   ������O�ƴ�1��Q�3��(��hp��Z�<�C=��R=�7=�^�<��=<�P�.���G�R����X��i���TԖ�D{���N�����@��<TA�<:�,=H}H=h�8=�v�<��F��ܞ���7�^����Q
��R��ݕ���ʿ�f�
�$�[�I�vq��Ό�WJ���,��c��	3��@?������h�p�$�H�&�#�(m��.ɿ�   �   ����S��]�ᢩ�J�7�������|��<��P=�Wg=�R=|�=(��<�tT;�-~�Rj��;��^�|�k��a�l@�Ƭ��s�� pk:D�<.�=(H=��\=�+F=���<��D�Zc����;�>��B���U�ޅ��Lο�����'��^M�-�v���������-���w�� (�� ݡ�q����u�^3L�He&�3��m�̿�   �   燔���O���0���3��&��`h�`]�<tC=Z�R=�7=l_�< �=<�P�.���G�W����X��t���[Ԗ�J{���N���h�@�`<�A�<��,=�}H=L�8=dy�<H�F��ڞ�j�7�l���;Q
��R�Nݕ���ʿ+f�R�$�f�I��tq�/Ό�hI���+���a��
2��X>��ڙ��2�p�8�H�t�#��l��-ɿ�   �   �
���D��� ��>��;O(�z����<#�(�<N=��=t@�<@|�;h:����E�I���z�ʽ����
m
�����3���4Ͻpƞ��P���¼�|�: o�<��	=L�=�ګ<�5P����>�+���$h�:�F��"����������3o���>�#Fc����Y֓��Ǟ�ȸ��R������#��� c��%>����Ճ���y���   �   gD����3��	꾢쌾��@����D�(�^<�!�<�n <��@�X�,��$���>��n��@A�0�\�o��u�np���^���C��y!�˨������Z�8�o����;|l�<�a6<�n��ֆ�;��Ɏ��E쾄�4����������s��:x.��eN���m�}������Z��v$��oׄ��Un���N��n.�����2�<3���   �   �_d���s�˾Ŵs��.���e�\���9�򻨕�9���l�O(���a�'��b��������Ǿݫ̾X�ȾB	���;��O����e��+�d�{}��h�@�!�`-������Go�����v��l;Xc��8e��霿D�̿y �����5�O�O���e�ٰt�dSz�Lu��|f��zP��|6��*� �Ww̿㏜��   �   �	B����\/��	�I��nؽH�N��˼hżbh6��$�����	�S�ˀ���E���侬U�(��=N���g��I��\z�Ξ��Ľ�KΓ��W�yg�����nY@��xּ�uۼ�*V�4*ܽ��K����F��GB�����ί��ܿJ����]�0��A�-}M���Q�"N���B�@�1�������gݿ� ������   �   �&�־OǇ�7���M����C������^��ÿ�XW�~.q�����w������m+�3�D� Y�Lf�0�j���f�
GZ��sF��-��p�X�徎�� �t�VW!�c�Ľ8{f��#�lkI�O���!� ����� ־z��3�[�|��H���!޿���J���& �T#)��y,�ެ)��!���V����߿g������T�\��   �   �[��ڔ���N��F�� ���K��%o�T��#��GPz�2G��th��Ė$��dL�o�r��_�����h��닣�Y࠿����3l��&�t��iN��K&�����P���K}���!��oý��s��N�h�����M�>���P����,�Og�P��r9����ѿ����=�B�\�
�ɯ����f��Õӿ]����&��M�h�r�-��   �   �@��dHo�6n�#q���ui�b�h� \��zg���m��派\}�sG/�h�a�����;@��� ���!ʿ�6տHBٿ��տ�D˿�c�������̋�n�c��0�����D��No��q��u��Jyi���h��X��Bd��m�J㴾�z�8D/�d�a�B���v=������HʿS3տ�>ٿ%�տFA˿�`������ʋ�c���0�΁��   �   "E}���!�tiýМs��N��������M����T����,��g����<����ѿ �?�D�b�
�ʱ��������ӿ&����(��,�h�~�-�'`�����QN��K�@#����K�� o��N���� Jz��B���b��K�$��`L���r��\�����se������/ݠ�����^i��
�t�.eN��G&����$L���   �   �Q!��|ĽZqf��#��jI�O���t� �����#־��� \��}������Ӂ޿������( ��%)�6|,��)��!�������߿޲�������\�K)��־�ɇ�"���P����C�����^� ���_R��'q�;������y���i+���D�Y�f���j���f��AZ��nF�d-�m�I�徶�����t��   �   �ﰽtM@��iּ�nۼ+V�v,ܽ`�K�������IB����]Я� �ܿdK�]��B�0�L�A��M��Q��N���B�?�1������jݿ�"��K��lB�T���1���I��qؽT�N���˼T ż�]6��������S�a|��[@����R�B��J����=��O���v�>��O����ɓ���W��a��   �   ���x�!�0��`���hHo����R�v��n;�d��:e��ꜿߟ̿z �E��f�5�8�O��e�Z�t�Vz��Nu�3f��|P�f~6�^,�6 �.y̿^���bd�ŋ���˾ķs�f0���e����@��P���~�1��yb��(��a�z"��#���K���n�Ǿ��̾1�Ⱦd��B6����6�e�4�+��X��t���   �   �2�;,y�< q6<Pn�h׆��;��ʎ�HG쾞�4��	�������H��My.�4gN���m�~����� \���%���؄��Wn�D�N��o.����e4�~4��cE����3����팾��B��P�D��_<8,�<�� <��@�t,�����3ｔh��9A�U�\��o���u�p���^�"�C�*s!�^���k}��ܷ8���n��   �   ��	=v�=�߫<P1P�M�����+�����h���F�~#��F��������o�z�>�.Gc�K��'ד�oȞ�����B���������c��&>�i������z��G��(�D��� ��?���P(�¸��x>#��!�<n=ޘ=0N�<�Ã;$���E�x�����ʽ%��ѷ��g
�����)���+Ͻ;�����P���¼���:p~�<�   �   րH=��8=h|�<�F��ڞ���7�����fQ
�.R��ݕ���ʿ^f���$�ŋI�Nuq��Ό��I��V,���b���2���>��J����p�ɌH��#��l�z.ɿ[���Z�O�����0����3��'��0k�^�<� C=��R=7=�g�<��=<�7�x��RG�ְ���S������qϖ��v��F�N����@��<�K�<��,=�   �   61M=�Y5=���<�o��������L��U����]�c��ӡ��hڿ
p���1��M[�p���.��������Ӽ��g��м�0���c���.;���~Z�d1�\��s;ٿ�砿NVb����Y����dJ�[���t"��t��<��:=\�R=��<=��=0�}<����Hļ�5*��+c���������˄�h.f�I.� μІ����g<U=�t7=�   �   ��7= '=��<�d��Iٴ�`�H���������_������ֿ.���.�|W�HŁ�G9����������c��� ���j��老�IlV�`.�dq
�>�տ�.��RK^����S���-F�D���O��x��<ȩ,=�X==�
 =d��<�i�;����f$!�,�p��͗�'&��Ov�����2e��t�t��0&�x��@*@;�.�<�j=�   �   H#�<l��<8�}<ē��f}���><��ت������S�t�@̿3R�	�%�8BK�~�s��U�����(���q���@���5��x\����s�3�J�v%����f˿�>��@�R���
��z���:��립�"��DG�<D� =\��< q�<`�s��O����p���������R�B��&T���ZB�F*�T洽*�v��k�� �����<�   �   �p:7<p/�;@���C���)��F���B��N�@�	C��󿻿��(p���9���\�i��������P��Ǳ���M���	��O�\���9��A��6��ŉ�&@�g����&��˰'��}��,���_�;(�M< 3;�䦼�V�bI���h� a/�T��Fq�6���t��h���wr�m�U��-1��G������]�`����   �   �&��e��Xg4��2ؼ����4��s����ܾ�K)�� t�,���&�ؿ����[$���A��^��v�����`ʆ�1��(<w��^��4B�/�$������ؿ�o��=�s���(��۾4Ԅ��i�M��L�ͼ�z��&������✽"D ���9���v�P_��0���ɾ�K׾O5ܾջ׾�Nʾc=��拚��Iy��<�~L�-x���   �   $Ƚ��e��D����T7}����)^��y�����(]O����������j��%�a<���N���[��{`�3\��O���<�:-&�G��	��l线h����7O�4e��뷾]�O����x��
��f��J`���Ľa��h����*_ʾ)����"�ou�Z'�>�*�b�'�����/0����˾�}���j��& ��   �   �1��ܽ�:���[H�xp��iɽ�1�����C�_	)���j�WК��ÿ�!�2�	�r���>*���3��j7�$D4���*��l�
���+�ÿ�6���k��.)��>��Q���o0�QȽ�l�8�D�{��d6ڽ�T/�윃�ѿ��c��S]�g�7��|R�6�g�&Zu�3z��u�}{h��{S�?�8��_�'���3�����   �   `@��q�1�ܽ�m���v���HD���`��W��b��:9�܈v�����)����޿�~�� 	����.1������	�ū��~�߿4o��WI���{w�4�9���驱��a��.�����6Gt�7#���Gڽ��0�+X���ƾ���@d0��Z�胁��g���u��A}������˪���U���8����[�=z1����OǾ�   �   k9ľ������"�[ǽ�r��1>��d�ƽ0 "�1l��l[þ���;�!�p�8���������Ŀ��ֿ�#�H�P�⿳M׿�xſX���q���r��<�q���5ľB�V�"�~Wǽ�q��@��
�ƽ4$"�;o���_þ����;���p�祓�	����Ŀ��ֿ�'��K���IQ׿
|ſK����s���r�T�<����   �   ��ꬱ��a�1�'���"Et�����@ڽ̋0��T���ƾi��T`0�f}Z�9����d���r���y������jȪ�����n��Z6����[��v1���]KǾ=����1�rܽ�j���v��!��G�R�`�/[�����v9���v� ������U�޿���� 	�ȇ�Z3������	�c�����߿�q���K��\w��9��   �   +1)�.B��S��$r0�kȽh�l�лD�D��A.ڽ�N/����������\��|Y���7��wR�ޭg��Tu�j-z���u�6vh��vS��8��[�!�� /��7���<1���ܽi6���WH��p�&mɽ�1�����QG��)��j�|Қ��ÿ�$���	�{���@*�b�3�2m7��F4���*��n���
�x"��ÿ�8���k��   �   �9O��f����]����N�x�&�
��^�f>`��ĽI��h����3Yʾ;�����8q��U'���*���'����%��s)����˾y��v�j�K! ��Ƚ��e�b>�����9}��!��T,^�?|������_O�J���/���n꿢k���%��<�N�N���[��~`��5\�O�O���<��.&����Y��K麿঎��   �   ;�s�`�(���۾_Մ��j����d�ͼhc���(���ٜ�J> ���9��v�7Z��`*���zɾ#E׾�.ܾZ�׾gHʾ�7��񆚾>Ay�<��F��o���	&�DU���U4��0ؼ���
�����v�ܾ�M)�B#t�����#�ؿ��|]$�ԶA��^���v�����ˆ�����>w�&�^�r6B���$����o�ؿ/q���   �   �ŉ�,'@������'��Ʊ'�1~��������;ȡM<`�;0˦���V�M?���b� Z/�)T�>q����:p���c��\or���U��&1��A�x뼽~w]�짳��1r:(!7<�E�;D���Ы��x�)�rH��&E����@�D��M���˝�8q��9�d�\����
��_���aQ������N���
����\��9��B�|�7���   �   ?���R�7�
�{���:��립� ���L�<�� =���<L��<@Us�`6���{p������彛M�����N�a�-=�� ��ݴ�ʬv��_��Ԫ�0��<�-�< ��<�}<Д���~���?<��٪����ϫS�B���A̿�R���%�JCK���s�eV�����)���r���A��k6��4]��ԡs�	�J��v%�O���f˿�   �   �.���K^� ������-F�(��,N�����<,�,=�[==� =���<���;�}���!�ʚp��ȗ�� ��q������H`����t��(&��q��@�@;T7�<n=�7=�	'=о�<f��Tڴ�R�H�t������X�_�����ֿ��M�.�!W��Ł��9��~�������}��猸��������0����lV��.��q
���տ�   �   �砿Vb�Ƹ����NdJ�˝��� �����<��:=ηR=:�<=��=��}<�}���~ļh5*��+c����������˄�r.f�6I.�|μ������g<�T=*t7=�0M=6Y5=L��<Lq�������L�,V��K����c��ӡ��hڿ"p���1��M[�����=�������Լ��g��м�$���S���;���~Z�L1�E��J;ٿ�   �   .���J^�F������,F����I��p��< �,=l\==< =$��<���;�}���!�ؚp��ȗ�� ��q������R`��~�t��(&��q�� �@;�7�<Vn=��7=f
'=x��<�a���ش��H�u������M�_�T����ֿ����.�W��ā��8��z���~���c��ҋ��������������kV��.�q
���տ�   �   �=���R�Ӯ
�<y��$:��覽����Q�<8� =���<|��< Ps�6���{p�����形M�ǎ��N�i�2=�� ��ݴ���v��_�@Ѫ����<�/�<\��<��}<�����{��x=<��ת���ҩS���W?̿�Q�g�%�^AK�V�s��T��3���'��}p���?���4���[��W�s�(�J�Ku%�7��e˿�   �   �É�r$@���� %��\�'��y���������;��M<��;�ɦ�N�V�0?���b�!Z/�2T�>q����@p���c��for���U��&1��A�K뼽�v]�8�����r:h*7<�b�;�v��\����)��E��CA���@�<B��⾻����Do���9�"�\�v����������N��p����L�������\�g�9��@�v�D5���   �   ͔s��(�g�۾G҄��f�����ͼ�R�������Jٜ�,> �{�9��v�;Z��f*���zɾ-E׾�.ܾc�׾nHʾ�7��񆚾3Ay��<��F�Ao���&��O��`D4�$#ؼ�����������صܾhJ)��t�ڧ��y�ؿ����Z$�D�A�~^���v�.����Ȇ�����9w���^��2B���$�]����ؿNn���   �   �4O�?c��跾�]������x��}
�\Z��;`��Ľ��h����2Yʾ>�����=q��U'���*��'����&��r)����˾y��J�j�! ��Ƚ��e��9�p��.}�����%^�Iw�����ZO����.����	꿪h�d�%�Q
<�j�N�D�[�'y`�[0\�i�O���<�b+&����x��R庿�����   �   H,)�;�O��yk0��Ƚ��l�h�D�����,ڽPN/�ݘ�������\��}Y���7��wR��g��Tu�p-z���u�:vh��vS��8��[�� ��/������1�W�ܽ4��ZPH�

p�Edɽ�0�����2@�)���j�hΚ��ÿ�쿆�	����z<*���3�Kh7��A4�u�*��j�H}
����ÿ�4��k��   �   �8�����`��*�����":t����>ڽ%�0�]T���ƾd��S`0�f}Z�;����d���r���y������lȪ�����o��Z6����[��v1���?KǾ�<��A�1�:ܽlg���v�/���@���`�zT��,��J 9��v�3���j|����޿h{��	����/�f����	����"�߿El���F��~ww��9��   �   1ľ����Z�"��Oǽ�j��99��@�ƽ:"��k��F[þ���;�!�p�9���������Ŀ�ֿ�#�H�R�⿶M׿�xſX���q���r�ߑ<�d��b5ľ��X�"�HTǽ�l��Y8����ƽ�"�>i��kWþQ�z�;���p��������a�Ŀt�ֿ �8D濄��J׿ZuſF���Sn��!r�,�<�����   �   J9��/�1��	ܽ�c���	v�����B���`�}W��T��29�؈v�����(����޿�~��	����01������	�ƫ��~�߿4o��UI���{w�*�9������&a�p-�C����9t�W��)9ڽ��0�Q��Jƾt���\0��xZ��~���a���o���v��Z���Ū�����t���3����[��r1����[FǾ�   �   �1�3�ܽ�.���JH�f	p�[fɽ� 1�����fC�V	)���j�VК��ÿ�!�2�	�t���>*���3��j7�&D4���*��l�
���*�ÿ�6��|k��.)��>澇Q���n0��
Ƚ�l���D������%ڽI/�=���ܵ���V���U���7�/sR���g�Ou��'z���u��ph��qS�}�8� X�����)��#����   �   �ȽF�e��1����n.}���)(^�ey�����#]O����������j��%�b<���N���[��{`�3\��O���<�9-&�G��	��k线g����7O�$e��뷾 ]�n���x��{
� T��0`��Ľn�nh�����Sʾ������m�TQ'�V�*���'����B���"����˾t��]{j�� ��   �   b�%�=��(-4�Lؼ1���!��!���ŷܾ�K)�� t�.���)�ؿ����[$���A��^��v�����bʆ�2��(<w��^��4B�2�$������ؿ�o��:�s���(���۾�ӄ�~h����D�ͼ�@�p��v���М��8 ���9���v�SU���$���tɾ�>׾#(ܾ�׾7Bʾ2��ف��p8y��<��@�2f���   �    �t: E7<@��;�s��ԧ���)��F���B��I�@�
C��󿻿��'p���9���\�i��������P��ȱ���M���	��P�\���9��A�!�6��ŉ� &@�J���m&��
�'�T{���������;��M< h;|���"vV��5��]�jS/��T��5q�Z���k��:_���fr��U��1��;�<Ἵ�f]������   �   4<�<��<X�}<D����{��><�xت������S�u�@̿3R�
�%�9BK�~�s��U�����(���q���@���5��x\����s�3�J�v%����f˿�>��=�R���
�_z���:�(ꦽ����T�<�� =��<ܐ�<��r����fmp�����彈H�b��I��
��7� �=մ���v� S��~�����<�   �   ��7=�'=�ĭ<�_���ش�'�H���������_������ֿ.���.�~W�GŁ�F9����������c��� ���i��老�IlV�_.�cq
�>�տ�.��QK^����D���-F����dK����<N�,=�^==� =ģ�<ȍ;�p��<!��p��×�����k������Y[��B�t�V &�0c��@�@;B�<xr=�   �   ��F=�H.=lڪ<��qG½�nT��1���$���i�T�����߿�����6�B�a����yr���2�������v������,��d������+�a��t6����8�߿b¥���i����ʾ���S��K������ҭ<�/=� H=<�1=��<��E<�����\�<��v��卽�[��{���uw���=�����(�V@<�D�<0k0=�   �   ��0=�= ��<T���u����P�zb���4���e��+��Z*ܿX���|3���]�&*��͝�j
���h��D��oj������Ý�#���e]�LL3��l���ۿ�򢿤ee�L�������vO�;���Ĺ���v�<�!=^$2=�+=��< �&:,����4�����ِ������A��zR���������\5��j�� W�9|,�<v�=�   �   (8�<�,�< �V< p�����RC�tf����w�Y����uѿİ��b*��HQ���{��|���"��欲���������*��p����{��/Q�(C*����=ѿ��<EY�${����.�B����lW����\<���<��<��d< ���������������I���Na �F��v��x�˾��ʃ� p�����^<�   �   �Q�h�< #;��ͼ�椽�j0�;z��o��F����ϭ�����������>���c�M���S��G���,��DS���e���\��p�c���>�n|��������&獿�MF�S�m2����/�5��8$˼ -9;�=<����Оʼ��k�d�Ž�����7��X]��"{�b'���}���<���r{�G�]�5=8��D���ƽʛm���ͼ�   �   �5��� �e���������L�m��I��xU.��	{�44����޿�]��)�4�G��ke�!��`��P����o��Q� �e�$�G��)�nd�<�޿�&��}�z�84.���㾷7��2��|���R��r`��)��Di3�~ƨ�y����B����j���㺾;�о�޾؏㾦�޾��о+��������2IC�[������   �   Prҽ�v����L���k��<� ��f�}�������U����߿�!��_d��c*�Y�A���U���b��g� c�0�U��	B��*������￿߱���{U��	����Hff�r� �i䆽������(u���ѽt0&�LEr��Y����ѾPB������"��,�V"0��,��"�� �k���sFҾ鸤�h�r���&��   �   C58����3B����X�-߀�D_Խ��8�Eߘ�"��KR.�ζq��N��6�ȿ�����@ �\B/��09�ڵ<��J9��m/��q ������ȿl��l�q��^.����՘�9b8��Խ}����W�����E��7�����������&�=��#Y��n�+�|����
�|�� o�hY���=����z����!��b���   �   ���#9��e��ꗽ(+��h������i������'���>��~��<��Z
Ŀ6C�nT����ʇ�y,�����|}���LĿ�m��<S~�1
?�
@�F˷��i�����F��������潛�8�u֍�(S;e�(96�{za������ӗ��)��SP���{���e���O�����t����a�'�6����U�;�   �   ��ʾ����)��ҽz2���"��lUҽ��)�v���Afʾ���аA��Nx����8˲�<ʿM�ܿk[�q�,y迩�ܿ�{ʿ�
���T��ܧx���A�j����ʾ[�����)�3�ҽ�1���$��*Zҽҷ)������jʾ�����A�RSx����]β�?ʿ�ܿS_�u�
}�T�ܿ�~ʿ���xW��9�x�8�A����   �   BB�^η��i����HH�����X������i�8��ҍ�"N;�a�!56��ua�灅��З��&���L���x��<b��}L������β��u�a�\�6������;���9�`�藽
+���j�������i����
*��>�2~�@?��\Ŀ�F�[V��������.���� �W�Q���NĿ-p��W~�.?��   �   a.�?��ט��d8��Խ�|��x�W�^����<��7����V������Ў���=��Y���n�q�|�7���^�|�t�n�cY���=�,��>������\^���/8�~�罺=�� �X��߀��bԽ׆8��ᘾ����T.�L�q�,Q��߫ȿ2�����0B ��D/�839�k�<� M9�<p/��s ������ȿn����q��   �   �}U�R�-����hf��� ��䆽޸�̴��u���ѽ2*&�*=r�oT��b�Ѿ1;�������"�y�,��0�`�,�ҹ"�������@Ҿ�����r��&��iҽ��v���$��m��� �t�f�(�����:�U�ů��/῿ƃ��e��e*���A�L�U���b���g��c���U��B�ؒ*�a��F���b����   �   ��z��5.�����8��i������M�([`����v[3�0���z���B������d�� ޺�ԥо_�޾����޾U�оF%��󳟾_��BC������(�4�d�����e����9����N��n�����RW.�V{��5����޿3_�l	)�$�G�Kne��#�Gb��ۋ��uq���S�X�e���G�%)��e���޿(���   �   �獿&OF��S�j3����/����� ˼�p9;�X<�Ķ���ʼ�k��Ž���~�7��P]��{��"���x��o8���i{�e�]�=68��>���ƽ �m���ͼ�:�0�<@?#;��ͼ9褽Ql0��{�������F� ��1���F���͈�8�>���c�0N��U��lH��n.���T���f���]��
�c���>�X}����#����   �   ;Ú�FY��{�m����B����,U���\<��<@%�<X�d<����������������PD�;���[ ����&��Zn��¾�&Ã��c������^<�B�<h3�<��V<q��i�����C��g��Ǵ���Y����vѿn���c*�JQ��{��}���#���������ô���+��7���(�{��0Q��C*����X>ѿ�   �   ���ee�|�������vO�#��������y�<!=�'2=,0=L�<��(:���24�*���������|<��,M����@���S5��\�� 9�9�5�<��=
�0=��=���<���������P�<c��W5�f�e�0,���*ܿ���*}3�;�]��*���͝��
���i������j��;	���Ý�p��Wf]��L3��l�"�ۿ�   �   ?¥�c�i�����ʾ�"�S�SK�����\ӭ<d�/=H=��1=��<x�E<0�����<�Ʋv��卽x[��~��vw�"�=�,�鼘)�8U@< D�<�j0=F�F=(H.=8٪<����H½QoT��1���$���i�{����߿�����6�b�a�����r���2�������v������,��	d�������a��t6�p���߿�   �   5��de��������VuO�l��������|�<�!=4(2=z0=��<��(:����,4�2�������"���<��9M����D���S5��\�� I�9�5�<<�=��0=d�=p��<h���̂��iP�7b���4�V�e�z+��*ܿ"��^|3�$�]��)���̝��	��th������i��0��Ý����Be]��K3�:l�5�ۿ�   �   �����CY�<z�|��I�B�����L����\< 
�<<'�<��d<P������������� ��TD�F���[ ����-��cn��¾�Ã��c���� �^< E�<�6�<��V<�h��)���1~C��e��W����Y�l� uѿJ��*b*�HQ�e�{�|���!��᫲���������)���~����{��.Q�RB*�e���<ѿ�   �   捿VLF��Q��0��Z�/�0��h˼`�9;�a<�����ʼ��k���Ž���~�7��P]�{��"���x��v8���i{�k�]�>68��>���ƽ��m���ͼ��@�<�y#;�ͼ�㤽�h0�	y���~�̂F�������&���̆���>��c�L��R���E���+���Q��sd��p[����c�!�>�Z{����������   �   ��z�W2.��㾿5��<������?��I`�,���Y3�����X���B������d��޺�ݥоh�޾���޾^�оM%������Z��BC���������4���(�e����ײ��{J�k��"���S.��{��2����޿�\�|)�o�G��ie�e�L_��ƈ��zn��DN�ęe�6�G�6)�0c�>�޿%%���   �   �xU������	bf�*� ��ކ�^�����u���ѽ�)&�=r�gT��_�Ѿ1;�������"��,��0�e�,�չ"�������@Ҿ	�����r���&��hҽʌv�Z�����:g���� ���f�����A�U�����ݿ��~��b�!b*�2�A�-�U��b�0�g�B�b���U��B�$�*�S��D���#����   �   \.����Ҙ��]8��Խ�v����W�����F;罤�7����G������ώ���=��Y���n�x�|�:���c�|�x�n�cY���=�*��5������;^��b/8���^;��v�X��ـ�vYԽ�8��ܘ�����O.���q� M��Ǧȿ ��>��> �@/�>.9�N�<�H9��k/�ro �(����w�ȿ�i����q��   �   ~=�|Ƿ���i�T���?��`ꃽÍ����潸�8��ҍ�N;�a�56��ua�灅��З��&���L���x��?b��~L������ϲ��t�a�W�6������;��i9��]�䗽o%��b��=��4�i�:���F%���>�&~�V:���Ŀ�?志R�������@*�������{����	IĿBk��O~��?��   �   $�ʾ����y�)�8|ҽ�*�����.Rҽ��)�+���fʾ���˰A��Nx����8˲�<ʿR�ܿp[�!q�/y迬�ܿ�{ʿ�
���T��ڧx���A�^����ʾ�����)���ҽ~,�����zNҽ@�)�n���$bʾ���L�A�NJx�T��8Ȳ��8ʿ��ܿ�W�0m�Iu���ܿxʿ���R��2�x���A�i���   �   ���69�W�����]$���c��|��.�i�O���{'���>��~��<��[
Ŀ6C�oT����̇�|,�����~}�	��LĿ�m��8S~�(
?��?�˷�F�i�+��HB��Gꃽ�������"�8�4ύ�nI;�^�W16�%qa�F���͗�a#���I��u���^��:I�����������a�S|6�d����;�   �   n)8����6����X��ـ��[Խ|�8��ޘ����@R.�ȶq��N��6�ȿ�����@ �\B/��09�ݵ<��J9��m/��q ������ȿl��g�q��^.����2՘�a8��Խiw�� �W������3�>�7���\��������6�=��Y�B�n�Й|�X�����|� �n�^Y��=�9���������0Z���   �   �_ҽ�v�:�����dg���� �.�f�=�������U����߿�"��_d��c*�[�A���U���b��g� c�2�U��	B��*������￿ޱ���{U��	�Ď��gef� � ��߆�>�����~u�@�ѽ)$&�m5r��O����ѾT4�����~�"��,�40��,���"�	�g���p:Ҿ�����r�e�&��   �   ��4��ݤ��{e����H����K��l����mU.��	{�44����޿�]��)�4�G��ke�!��`��Q����o��Q��e�$�G��)�nd�>�޿�&��z�z�/4.�\��d7����	��(>��7`�� ��jM3�+��������B�4����_��Mغ���оˢ޾S��Y�޾��оl�����������:C���W����   �   ��庐�<�#;��ͼ,䤽�i0�z��b���F����Э�����������>���c�M���S��G��-��ES���e���\��q�c���>�n|��������'獿�MF�S�52���/����`˼ �9;�x< ���\kʼ�k�0�Ž�����7��H]�z{�I��Tt���3��3a{�a�]�/8��8���ƽ�zm��ͼ�   �   �Q�<�?�<��V<�f��m����~C�Rf��޳�v�Y����uѿŰ��b*��HQ���{��|���"��笲���������*��q����{��/Q�(C*����=ѿ��:EY�{������B����M��X�\<��<�1�<he< 5�����s���u������?�����U ����|�yd�
���j����V�@Y�@_<�   �   ��0=��=���<���������P�jb���4���e��+��Y*ܿX���|3���]�'*��	͝�k
���h��F��nj������Ý�$���e]�LL3��l���ۿ�򢿢ee�J������HvO�w��� ���<}�<L!=�*2=�3=��< *:\���D4�����ˆ�����-7���G������bK5��M�� m�9t@�<h�=�   �   [J=�,2=(��<x׫�d�����Q�oD������h������/޿��LO5��/`�����o-��Ҵ��a���
���d��Iߴ��L��/����`�!�5�UP���޿x7��G�h�@T�z���
S�:����i����<��/=��G=��1=�0�<�xG<�}��`���:��t�B���c���݋���r���8��߼����Q<�k�<$?4=�   �   ��4=�#=�l�<,���KѺ�frM����������c�L��ڿ��X02�o�[�#������춰����ʞ����A�������I��QO\�M�2�@���&ۿFe���d��f��O��ʭN�ü�k�����<2� =�1=�=�g�< �I:,����2��t������F��,���۴�iT���i���0�pZ���F�:�ʰ<��=�   �   (��<�|�<��h<즲��p��	A����t�[�W��̙�B п����@)���O�C+z��r�������e������,Y��5��"p��Hz�hP���)��
��wп8/��nqX�����\��(B�,?��hʸ�`�]<�!�<�:�<X�e<p�������6���꼽�J�M��~�����>��������q�����	� ߻�p<�   �    ���� < �l;x�ü����,.��松�c���D� ���l���i�������=�bwb��|���^���/��:������=���`���]b���=�ٷ����������M���uE�\��Y��v"/��2���+ɼ�B;��<��� ɼ��j�n Ž#���6��1\��y��F��,y��Z��cy��h[���5��7��5ý�Dg���¼�   �   �8/��ᚼ�}R�X������S�I������-� by�B-��҈ݿl�
�r5(���F��?d���}���������i��IX}���c�dhF��(�*�
���ݿ3O��z�y��[-�pe�=���\�	������\��C���=2�����>�Q�A�1����������Ͼdeݾq�N,ݾ�/Ͼ�|���#���3��@�f�5=���   �   ��ν��p�|��F��j���s����md�@+����T1T��ޑ�쾿�n�_���)�7A�ĆT�ޢa�N2f��ha��'T�C�@��_)�2���.￫Ҿ��ݑ��JT��7��z���e����������0�@os��|н�x%��Qq�����Ѿ�<���L���!���+�	/�i�+���!����p��Hо���>p�{$��   �   G�5����Vv����S�d�|���ѽ��6�?���KV��P-�zp�񕞿6�ǿ����M�j��F�.�%J8�T�;�H8�>5.��K�f���l�ʂǿAc���Ip�DB-��`�$З�7�l=ҽ�Q~��U�W���j����6�*~��b���o"�������<�NBX�ιm�`{�����&{�IRm�T�W��X<�py��>��E���퇾�   �   ���07�4N�m���ꁽa���z��!h�P����j���=���|����� \ÿ���� ��o����^����,�H� ����A�¿pD��R�|��=��B��i��xh�����]���\��5
��R*�o�7��"���m̾/����5�:�`�
���@��x���{��Ƅ���R���/��;斿Ҭ��k`��4�ai�8�˾�   �   l�Ⱦ<����,(��Ͻ,#���7���Aн�q(�ƅ�W\ɾU&�8�@�bw������/��z�ɿ�ۿ�M翉2�2�jWۿ�
ɿ'����+����v��m@�w��v�Ⱦ����$)(�\�Ͻ@"���9��~Fн�u(�*Ʌ��`ɾI)��@��fw�I����2���ɿӿۿnQ�w6�
�[ۿ�ɿ$���[.���v�q@�)���   �   #E��l��yh�Ӎ�<_���[������#�D�7�;���h̾����5�q�`�^���=��;u���x��W����O��],��I㖿0�����_�Z�4�^f���˾�����7�xH�@j���ꁽ���\}�Y&h�֐��8m���=���|����_ÿ$���� �r�0��A`�:���.�� �����¿�F��&�|��=��   �   �D-��c�Mҗ��7��?ҽ2Q~���U�}����
�6�#z��$���������,�<�<=X�X�m�cZ{����� {��Lm�f�W�pT<��u��8��7@���釾��5�#���q����S���|�ɋѽ*�6�ӳ��Z쾀S-��}p� �����ǿ���O������.��L8�ߤ;��8�7.��M����o�8�ǿ:e���Lp��   �   �LT�b9��|��H	e����8������'�`bs��sн�r%��Iq������Ѿ�5���H�C�!�,�+�w/��+�Q�!�����i��8Bо� ���p�Ju$�A�ν��p��������������pd��-�����3T�\���D�q������)�zA�[�T���a�.5f��ka�L*T�i�@��a)�����0ￖԾ�iߑ��   �   ��y�]-�lg�t������	����}\��0��02�Q�E����A��,��b���������Ͼ�^ݾ�⾱%ݾ�)Ͼ7w�����+���@�����4��,/��К��kR����m����T����|�Ὰ-�~dy��.��Ԋݿ��
��6(���F��Ad�K�}�,�������k���Z}���c�(jF�=(�B�
���ݿ�P���   �   lN���vE�+��W���~#/�s3��x(ɼ�XB;H< ֦��ȼ��j�!�Ľ��z�6��)\�*�y�SB���t������y��`[��5��1�7,ý05g���¼�|�@� <��l;T�ü�����..�M蝾e��E�	��Vn��Rk������=�(yb�~��`��1���������P>���a��W_b���=�¸���������   �   �/��9rX���p]���(B�s?��0ȸ�x�]<�*�<lG�<��e<�.������.���Ἵ�@�FH�By���\9�p���w�����V�	���޻�q<��<��<�h<ܧ��<r��|
A�6����t���W�Z͙�Lп5���A)���O��,z�gs�������f������2Z��"���p��@Iz�KP�E�)�s�hxп�   �   ~e��\�d��f��O����N��¼�Ti�����<�� =X�1=�=(r�<�bK:����v2��o�����_A�����pִ�hO��e���0��L��@��:�Ӱ<8�=�4=R�#=�m�<����TҺ�YsM�K���&��Q�c�����ڿo���02��[�x#��>���~���l��[���������������I���O\���2�u��''ۿ�   �   T7��
�h�T�3��R
S�����Xh��l��<�/=R�G=��1=x1�<pzG<0|��_会�:�Rt��A���c���݋���r��8�`�߼���Q<4k�<�>4=�ZJ=R,2=���<٫�����T�Q��D����h�ķ���/޿+��hO5�0`�����-��Ҵ��a���
���d��>ߴ�xL��/��h�`��5�=P���޿�   �   �d��K�d�f��N����N�G����d�����<�� =��1=6 =�r�< mK:�����v2��o�����hA�����wִ�rO��e���0��L����:�Ӱ<��=��4=&�#=xp�<H򬼤к�rM�I���g��D�c����ڿؒ�02��[��"��W���t���R��<��������������#I���N\�͔2����9&ۿ�   �   g.��2pX�����[��/&B�3<��Կ���]<$.�<�I�<x�e<�+��r���.���Ἵ�@�KH�Ly���c9�w���w�����6�	���޻Xq<��<��<��h<����o���A�I����s���W��˙���Ͽ��*@)���O�*z��q������d������X��2��@o���Fz�NP�ʃ)�P
��vп�   �   �L���sE�0���}���/��.���ɼ`�B;x< ���<�ȼx�j���Ľ��z�6��)\�3�y�ZB���t������y��`[��5��1�,ý�4g�L�¼�$�8� < #m;�yü���++.��坾c���D�/���k��:h������=��ub��{���]��S.������#���;���_���[b�)�=�ö����"����   �   ��y��Y-��b�F���h������l\�0+��P.2��什����A��,��a���������Ͼ�^ݾ�⾹%ݾ�)Ͼ<w�����+���@����-4��t*/��˚�`ZR�Ф�����P�������e-��_y��+���ݿX�
�4(�ߨF�X=d���}�9�������h���U}�o�c�zfF�P(��
���ݿ�M���   �   HT��5��w��te����a���n��(#�\_s��rнWr%�qIq������Ѿ�5���H�F�!�1�+�~/���+�V�!�����i��4Bо� ��p�u$�d�νخp�>���������"���jd��(��"�/T�"ݑ�6꾿�l����K�)�A�F�T��a�o/f�
fa�8%T��@��])�����+ￅо�,ܑ��   �   �?-��\�>͗��7��6ҽ`E~��U��z����彘�6� z�����������,�<�>=X�Z�m�hZ{����� {��Lm�k�W�rT<��u��8��&@���釾s�5��但o��F�S�Ҽ|�ɂѽX�6�Ȯ���R쾂N-�wp�������ǿ
��7L�k���.��G8�Ο;��8��2.��I�����i�'�ǿa��"Fp��   �   e@� f���h�\���V���U�����Z!彑�7����h̾����5�p�`�^���=��=u���x��Z����O��`,��K㖿2�����_�W�4�Yf���˾�����7�GF佹f��$偽f
���v��h����{h���=���|�3���RYÿt|�&� ��m�����[����*�`� � ��G�¿�A��$}|���=��   �   ��Ⱦ���$(�l�Ͻ]���2���>н�p(��Ņ�)\ɾJ&�1�@�bw������/��{�ɿ�ۿ�M翍2�6�nWۿ�
ɿ*����+����v��m@�o��O�Ⱦ8���,((�)�Ͻ4���1���:нm(�Å�:Xɾ�#���@��]w�󒗿�,��"�ɿw�ۿ�I翢.�V翸Sۿɿ���
)����v��i@�~���   �   Ӫ���7��?��b��䁽���%y�� h�����j�w�=���|�����\ÿ���� ��o����	^����,�I� ����B�¿qD��P�|��=��B��i���h�2��AY���U��( �����7����d̾���*�5��`�����:��r��+u���}��=L��")��F���x���!�_�Y�4�"c���˾�   �   ��5�hw�2j����S��|��ѽָ6�鰗�V��P-�zp��6�ǿ����M�j��F�.�(J8�W�;�K8�>5.��K�h���l�̂ǿAc���Ip�:B-�^`��ϗ��	7��9ҽ�F~�X�U�8v��M��7�6�Jv��+�����������<�S8X��m��T{�>��E{��Gm�^�W��O<��q�2���:���凾�   �   9�ν��p�,�����规������ld� +����M1T��ޑ�쾿�n�_���)�8A�ĆT��a�O2f��ha��'T�D�@��_)�4���.￬Ҿ��ݑ��JT��7�jz���e���������V����0Ts�[jн�l%��Aq�����$Ѿ�.���D��!���+��/�x�+�!�����b��!<о����pp��n$��   �   �/�h����BR���鼇����Q��������-��ay�A-��Ԉݿl�
�s5(���F��?d���}���������i��JX}���c�fhF��(�,�
���ݿ5O��{�y��[-�Ge�섉�F������(Z\�����!2�N秽�����A�K(��Z������r�Ͼ)Xݾ��ݾP#Ͼhq�����*"���@���� +���   �   ���8� <�em;�vü����+,.��松�c���D�����l���i�������=�`wb��|���^���/��:������=���`���]b���=�ڷ����������M���uE�O��"���!/�0���ɼ �B;�"<������ȼ�~j�D�Ľ����6��!\���y��=���o��N��/y��X[���5��+��!ý0$g�t�¼�   �   `��<��<8�h<`���Ho���A�죮�t�V�W��̙�C п����@)���O�B+z��r�������e������.Y��4��$p��Hz�hP���)��
��wп7/��nqX�����\���'B��=��������]<�4�<T�<��e<���n���'��ټ�7�C��s�b���3�%��:��Jn��w���f�	� m޻1q<�   �   Ȟ4=~�#=�s�<�𬼈к�*rM�{��������c�L��ڿ��Z02�n�[�#�����������˞����B�������I��RO\�O�2�@���&ۿGe���d��f�|O����N�O¼�|f��\��<�� =>�1=�#=x{�<��L:t~���n2�?k�����;<��y	��.Ѵ�hJ��V`��.�/��=��@ɼ:<ް<��=�   �   �xX=.A=,H�<xy�؉���E��������":^�:%���տQi
�p.�ojV�>����%��s���˵��:=�� ���_ɫ�Rh��=��dW��/�[H��׿�F����_�P����h'H��w���:��TI�<�:=�Q=�<=��=pd�<��z� ��p�$���[�Z~~�ℽ�|�~X�B������@�H�<ʒ=� C=�   �   BbC=J�2=�_�<�v{�5 ���@�`&��!�f@Z�6w��>,ҿ.�+�*xR���}��Д�#̧������������֧�����ym~�,MS�:�+�
���ӿƆ��c�[�HD�4����C�|Ϯ��(��0��<��+=Vi<="o=t��<@Z�;�3��j���Yj�����ܦ�	 ���Υ�����	e����<{�Щ�;���<Zt&=�   �   �=�l=��<����@��	5�L���^����N�R����ȿs��g�"�{CG���n��e�������}��P����a������2_��$"o���G�jK#�NK�sɿ�����P�	��s����7�j���<:��1�<�b =�$�<<�< _`�,"�4l��ɮ�TD��z�|��0�Bs��U��/޽�6����d��ἀaͺt��<�   �   l�;��l<��
< q��m򑽹 #�0��������<�Lb��� ���3����o6���X�{��V��3l�����29��F���z���X��y6���h�ￊ˸�F���z�=��������ZU%��ܢ�P��;��P< �,;,��j`S��ö����,���P�xm���H����H~���k���N�n�*��F��B��&�J�,<���   �   j��0�Z�����P	���Ђ���:����H׾[�%�`To�����yfտ}��6�!���>�n�Z��r��J��m���
��k�q���Y�(U>��!�����տ�����p�sI&�8�ؾ�͂����2��H�Ƽ�^�xjv���\���'[��,�7���s��`�������Zƾ��Ӿ��׾%Ӿ�bž�^��.���O�p�S�4�Le��OG���   �   ���b�T��/���= �\m��7�[�W���������K�G@��X跿U��T����#���9��L��8X��W\�n�W�,4K�$�8�4�"��#�Q�(����;��a�K��IǴ�%Y���pr�\��p��[�{���(��[e�C��RȾ���eC��,�Τ$���'��F$�R���e���%ƾ����njb�����   �   
�*���ҽ�~���9�ʀa�a��*�+�������&�g�*���k���i}��`����!"(�M1�uW4���0�f'��(�4���Q�d뿿?8��2�f���%���ᾋZ����,���½�ae�B>����/ֽR�,�jꁾٍ��i�񾚡��y5���O�4�d�4�q�<�u�Gq��c�0�N��34��k��{�mδ�.����   �   9��l�+��ӽ� ����h�5J��VA��[����V���S6�_Vs�	Ú�Nu�� �ܿ3������K������5����n���:ۿ�X���,9r�a�5��;�Y����[��d�����)k�w����<սLj-��N��{nþ?�_c.�1X���������h������ᪿ#���j����ᐿ�|~�ŏV�t-��������   �   �W��
�|�!�����r������g����z�O)~��S���/	�K9��n�3��0֫��i¿��ӿ"߿��⿶�޿;ӿ�R��:������	�l��-8�Dk��S����|������r��Q������w~�G/~��W��X2	��N9�Ln����:٫�-m¿p�ӿ�߿m��l�޿�ӿ6V��ª���:�l�718��m��   �    >�V����[��f�U���'k�𯈽86սPe-�$K���iþ ��_.��X���������e���	��sު�⫧�Q���ߐ�lw~�d�V��-��	�/����5����+�<ӽ5��<�h��L��D�h�[�P�����,W6�jZs��Ś�5x��Q�ܿ�������g������7�����q���=ۿ�[����<r�B�5��   �   ��%���ᾡ\���,���½^ae��<>�䩁�'ֽ��,��恾ǈ����̝�*u5���O��d���q���u��q��c�o�N�w/4�h��uﾴɴ�����Ґ*���ҽ�}�8�9�Ёa�s!��6�+����H�ᾃ&�wg�F�������p�鿱b����Y$(�cO1��Y4� �0�)h'��*�۠��T���):��2�f��   �   ��K���aɴ��Y���pr�������t[�����"��Se�:>��l�Ǿ���?��(�t�$�X�'�^B$�?}��a�j��pƾP���cb���ꗽ�h�T��"��`; ��m�*;콏�W�I�����6�K��A��n귿���٩�ȋ#�Ǯ9�b	L��;X��Z\��W��6K�*�8���"�5%�XS����/=���   �   �p��J&�$�ؾ�΂�P��3����Ƽ�G�hEv����i����O����7��s��[��󞱾�Tƾ�Ӿ5�׾��Ҿ�\ž?Y��S
�p���4�yZ��?��^���iZ�@d��t���т�g!�˾��KK׾�%��Vo����dhտ�����!���>���Z�p�r�L�������ܸq���Y��V>�>�!����b�տ(����   �    ����=�&������[V%�r�٢�P��;0Q<�e-;� ��>PS�������*�,�'�P�	m�)	��{��6@~�R�k�[�N�*�A�{9���J� %����;�m<��
<�p����\#���������p�<�Sc���!���5����fp6�|�X�${��W���m�����w:��i��ϐz�y�X��z6�����ￚ̸��   �   ����P��	�"t��u�7�����8���6�<<g =81�<x�<��_���%l�E����:ὦu��1+��m��P��&޽S.����d���� 5̺�ĝ<"�=(p=���<�������a5�g���5��ɲN�����ȿ��/�"�DG��n�}f�������~��T����b��r����_��E#o���G�
L#��K�,ɿ�   �   ������[�vD�g���C�jϮ��&��T��<��+=�l<=Bs=���<��;�$�����Pj�����צ�����ɥ�/���� e�X~�8"{����;p�<�w&=�dC=��2=�`�<�y{�/����@�'���� AZ��w���,ҿz.�|+��xR���}�є��̧�!���+������)ק�5���
n~��MS���+�?��@�ӿ�   �   cF����_�"�ۼ��'H��v��d9���J�<V:=��Q=N<=�=<e�<��z�x��*�$�.�[�(~~�ℽ�|�~X�^�����@D���<x�=� C=`xX=�A=�F�<�y�i���^E�>³����`:^�`%���տji
��.��jV�M����%��~���ҵ��:=�����Uɫ�Bh��.���cW��/�EH��׿�   �   L�����[��C�k����C��ͮ��"����<��+=
m<=�s=<��<`��;�$������Pj�����צ�����ɥ�6���� e�T~�"{�@��;��<�w&=,eC=��2=pc�<0q{�������@�&����@Z�w���+ҿ�-��+��wR�8�}�/Д��˧����������+֧�Z����l~��LS���+����Y�ӿ�   �   ͆���P�<	�Br���7������/���;�<�h =H3�<��< �_�l�%l�E����:Ὠu��:+��m��P��&޽[.����d�D���+̺�ŝ<�=�q=��<����v���5��������۰N�̧���ȿ���͵"��BG���n��d��̾���|��L����`������_^��� o���G��J#��J�sɿ�   �   <����=�P�������R%�약�͢����;�Q<�|-;����OS�v�����%�,�(�P�	m�2	��{��@@~�[�k�b�N�Ɲ*�A�[9����J��#��`��;Hm<��
<�e����"����������<��a������2�����m6�^�X�8
{�yU���j��A���7����׌z�N�X�zx6������6ʸ��   �   =p��G&��}ؾ�˂�A���-�� �Ƽ�6�`:v����ߡ��CO��ߒ7��s��[�������Tƾ�Ӿ?�׾��Ҿ�\žDY��U
�p�v�4�CZ���>������_Z��B��4����̂�i�û���F׾�%�jRo�?����dտu����!�7�>�d�Z�w}r�YI����Q	��߳q���Y�YS>�u�!����ƇտJ����   �   ɻK�+��~Ĵ�Y����$er�h�����q[��������Se�,>��e�Ǿ���?��(�v�$�]�'�bB$�B}��a�m��oƾJ����bb���������T����24 �Hm��2��W�r����u�K��>���淿����H�#���9��L�V6X�GU\�ҵW��1K��8�e�"�I"��N����:���   �   �%���᾽W��q�,���½�Ue�t5>������%ֽ!�,�b恾������ǝ�)u5���O��d���q���u��q��c�t�N�z/4�h��uﾦɴ�|���j�*�b�ҽ��}���9��va������+����M�ᾳ&�g�B�������z�G_����(��J1�U4�U�0��c'��&�v���N��迿"6��Җf��   �   �9�������[��`������k�g����3ս�d-��J���iþ�x_.��X���������e���	��uު�嫧�U���	ߐ�pw~�f�V��-��	�����5��W�+�!ӽ���r�h�fD���=�=�[�����'��Q6��Rs������r��ڍܿ�����~�9��k��u3����dj��Z7ۿ�U��G홿"5r�.�5��   �   gO��;�|�޻�?濽_k������8����y��(~��S��s/	�K9��n�2��0֫��i¿��ӿ$߿��⿻�޿@ӿ�R��=������
�l��-8�<k��S��4�|�Ϳ��꿽+m��Ҧ������;v�z#~��O���,	��G9��n����Lӫ��f¿O�ӿm߿ۤ���޿�ӿ�O��;��������l�1*8�eh��   �   !2��Z�+���ҽ-��`�h��E���?�
�[����C���S6�XVs�Ú�Lu����ܿ2������L������5����n���:ۿ�X���,9r�]�5��;�#���<�[�dc�����k������.ս:`-��G�� eþ0
��[.�+X�\��׬���b��c��'۪�����1���ܐ�.r~�ІV��-���L����   �   ��*�e�ҽD�}���9��ua����	�+����m���&�g�'���j���g}��`����""(�M1�vW4���0�f'��(�6���Q�f뿿?8��1�f���%�r��<Z����,��½We��1>�G���~ֽ�,��⁾������*���p5���O���d�A�q�"�u�[q���c���N�+4�Nd�{oﾡĴ������   �   G���HT�8
���0 ��m��4�y�W�}�������K�D@��W跿R��T����#���9��L��8X��W\�q�W�/4K�%�8�5�"��#�Q�*����;��^�K��Ǵ�PY�O��^gr�`�����f[�����J�KLe��9����Ǿ ���;��$�)�$���'�>$� y�^����ƾq���:[b����   �   ����:Z�P��\���9͂���缁��H׾O�%�]To�����xfտ|��6�!���>�n�Z��r��J��m���
��l�q���Y�)U>��!�����տ�����p�lI&��ؾ~͂���J/��h�ƼP%��v�������yD���7���s��V��u����Nƾ�{Ӿ��׾j�Ҿ�Vž�S��Yꕾv�p�W�4��N���5���   �   ��;H6m<��
<�b�����"�����q����<�Kb��� ���3����o6���X�{��V��2l�����29��F���z���X��y6���j�ￌ˸�G���x�=�|���]���T%��핽�͢���;01Q<�.;D袼�@S����8���,���P�� m�� �gw��~7~��k���N��*�0;��/����J��
���   �   �=�u=D��<��������5�+���W����N�P����ȿr��f�"�{CG���n��e�������}��P����a������2_��%"o���G�kK#�PK�vɿ�����P�	�bs��[�7�璤��0��x>�<*l =�=�<"�< _�0��l����t1὜p����%��h�yK�<޽�%���ud��t���ʺ�՝<�   �   >hC=��2=�f�<�m{�n�����@�O&���d@Z�4w��=,ҿ.�+�*xR���}��Д�#̧������������֧�����wm~�+MS�<�+�����ӿƆ��c�[�DD�%����C��ή� $��ċ�<�+=Xo<=�v=���<p��;���^�� Hj�Y����Ҧ�����ĥ�X�����d�8v��{�@�;��<�{&=�   �   .p=6Z=T�	= 6������/�ݍ������qM�@ے��ǿS	���!�y5F�ħm����+���ާ�������4���	��N�n�irG� #�0���ȿuh��u�O� ���y��B:4�嚘�(��0?�<��M=��c=��O=�=0\�<�x;�mj�P���r�/�xP�f�Y���L���)�t1輀lB���;T��<�+*=��[=�   �   v0\=$�L=�y=pL��ht��x�+��3��tN��I��Y��w�ÿ4���x5���B��i�D͇�Ğ��<�����f��)��������i�S�C��U �& ��ſϑ�G	L�H����c?0��'��hz�pX�<�H@=x�O=��4=���<`!@<���L7���=�~�v�I$��F���rv��TTp�D%5�L�ռ�Q��0dp<�=��@=�   �   !=،#=$��<�ϻ.L��� �ԉ��Z���>�>���2N���������8�I
\�b%��َ�E������"��������qU\��]9��R���󿬸���@����@�[���{����$��~��p�����<NF=��=5�<��;Xt����?���3DĽaC齪G ����¤������c���K��P3�����`q�;���<�   �   �FT<,4�<���<h��Vzn�"��h����S��.�&{��h���)߿���v�)���H���f�Vt���K��3X��X��:��"Df��_H�u�)��	���Q����|�_�/����L�����<W{�h�8�H�a<4�<��!<��9��(�ק�����r���<�_tV�kg�Knl���e��CT��*9��,���<h��\��0���   �   �Dм��|� �:p#Q���R�4���6j���ľ����]��@��Nǿ^���W��x1�bkJ��n_�څm�DHr���l�Jp^�.jI���0���mZ���<ǿ����a�^����B�ƾ�fm�g���]��
|�����pRܻ���F?���޽ȿ$�]�R�����jϵ��¾Z�ž�<���c��.���r뇾�X��� ���ֽ@v��   �   *,���t$��Z��x竼�R<���̽�~A��9��(� �*K<��K���g���׿�|�\����,��P=�Q#H�P�K�PG��B<���+�<��d��[�ֿO���D��E�<�� �*D��]�C���н�E��2��4^���/��æ�H�
�~�O�5�������Y߾�^�D�"����V��$O�� �F�ܾ}ϴ����\K����   �   ��Zi���1L����@52�4�������
Ͼ�U�CV����Bγ��2ڿ����������!%�*�'�[�$�g��I������g�ؿ����&q��t�U���!Ͼ:&������D��v8�����T��¹�Ph���k��6���r޾"�(���@��T�O:`��&d��_�ŽR��?�S3&�WU
��\۾������g��   �   ��p�"��t#���|\���9��]��|�1�E��ޞ����m�(�h�a�)���᯿�οV��;J���'�N;�y�����t�濭N̿x]��T���*a`���'��r�W��0�E��o�|����z=��a�񜸽,����s��*��(1��_!���H��"n�o����w��͈�����B������z����k��TF���)B��t��   �   ����>dd�Κ�?ͣ�ơV��_W���������@f�N#��O���+�+�]�����>��R|����ſBGп��ӿn�Ͽ�Ŀ� ��3���,���f�Z���)�֮��'���J_d�����ɣ��V�cW��������Ff�?'��������+�P]������A��}��)�ſ�JпB�ӿ�Ͽ[�Ŀ���������V�Z��)������   �   �v��Y��уE�t����4y=�n�a�ꖸ����6�s�u&��R+��d[!�<~H��n������t���������2��4����w��
�k�|PF�����<��M�}�p��}�6���w\�\�9�`����h�E��ើ*��f�(�1�a�z!��b䯿�ο̡��M���)�I=�g��������濟Q̿`��z����d`�<�'��   �    �$Ͼ0(������F���u8����l�T�,����b�M�k�/2���l޾����'��@��T� 5`��!d��{_��R�??�_/&��Q
�&W۾D���F�g��
��b���)L�8��$62��������Ă� Ͼ�W�9FV�����г�{5ڿ$���������6#%�Z�'�y�$�_���������ؿؼ���r��G�U��   �   X�<��� � F����C���н"E��+���O��f�/�Y�����
�,�O�����}���`S߾G[�1@�	����M��TK�5 ��ܾ<ʴ�����K����$���j$�tN��H㫼�T<�Շ̽ɁA�V<��� ��M<�M���i��i�׿�}�����,�S=��%H���K���G��D<�W�+�ˠ������ֿ���E���   �   A�^����ƾ-im�����]��|�@����ܻ����6��F�޽	�$��]���������ɵ�����D�ž�6��^������懾X�X�,} �w�ֽ�0v�.м`|�@��:�Q�v�R�W7���9j���ľ¬���]�ZB��ǿ�������z1�SmJ�8q_�L�m��Jr�J�l�pr^�lI�(�0���e\��x>ǿ4����   �   F�|�w�/�k��6���	��:X{���8�8�a<�#�<P"<�9���(�w��������R<�zlV�'g��el���e�<T��#9��&�=��f_��<��x��8fT<�>�<ࠈ<��}n���������U�m.��'{�:j��_+߿�����)��H�a�f�bu��M��_Y��v��9���Ef��`H���)�d
��R���   �   A��r�@�U�����L�$�@������¿<ZJ=b�=hD�<�h�;�\����?����.;Ľ�9齐B ��������*��([��D���B3�p���p��;l��<&=�#=���<�ϻdM��S� �ڊ�����X�>����!O����񿜑�q�8�p\��&��ڎ��E������#������@�pV\��^9��S����\����   �   Bϑ��	L�u�����?0��'��8w�T[�<�J@=z�O=��4=L��<�8@< ��x'�&�=��v�d��`����q��6Kp��5��qռ ��8yp<B�=��@=�2\=l�L=z=Q��Nu��L�+��4���N���I�PZ���ÿ�����5�
�B��i��͇�?������=�����������T�i���C��U �X �h�ſ�   �   Th��>�O�����y���94�c���@��D@�<�M=J�c=��O=$=�\�< x;�lj������/�<P�V�Y���L���)�t1��lB� ��; ��<�+*=��[=�p=�Z=�	=�;������`�/����%��rM�bے�"ǿh	���!��5F��m����5���ާ�������4���	��2�n�PrG� #��/���ȿ�   �   �Α��L������S>0��%��o� ^�<�K@=
�O=�4=���<x9@<���d'�$�=��v�h��b����q��NKp��5��qռ ��hyp<n�=�@=<3\=>�L=P{=�A���s���+��3��GN���I��Y��2�ÿ����85�)�B�ti��̇�`������@���
������^�� �i���C�1U �� ���ſ�   �   �?����@�����Q����$�=|������ǿ<L=p�=�E�<Pl�;\��l�?����(;Ľ�9齕B ��������0��3[��D���B3�������;|��<�&=|�#=���<0�λuJ��� �"���\�����>�����M�����Y����8�T	\�%$�<َ�1D������!��"�����AT\��\9�0R���󿻷���   �   ��|��/����ƽ���}��O{��8�Hb<8(�< "<H�9�$�(�=���z����P<�|lV�+g��el���e�<T��#9��&�7��H_�������8kT<�B�<h��<}��tn����T���R��.��${�h���(߿ֻ�t�)�?�H���f�Zs���J��W��2��+��OBf�^H�B�)���8��O���   �   �^�ݜ�̺ƾicm�����]���{� y��0�ۻ<��N6����޽�$��]���������ɵ�����K�ž�6��^������懾Z�X�$} �A�ֽ�/v�@+м��{� 	�:�Q��R��/��(4j���ľé���]��?���ǿr���&��w1��iJ��l_�x�m��Er�u�l�n^�;hI��0����2X��;ǿ����   �   ג<�8� ��A����C���нR�D����|F��l�/�d���X�
���O�����r���[S߾F[�3@�	����Q��XK�8 ��ܾ;ʴ����hK�Z��#��
h$�F���ի��I<��̽�{A��7��� �I<�+J���e���׿>{�Θ� �,��N=�!H��K��|G�n@<���+���������ֿX���B���   �   ��uϾ�#������>���j8������T�����{b� �k�2���l޾����'��@��T�#5`��!d��{_��R�B?�b/&��Q
�"W۾8����g�t
�]a��L%L�X��z+2�㉤�ú�C����ϾnS�F@V����̳�0ڿ�����������%���'�9�$�f��u��������ؿ:���*o��H�U��   �   Dn�S��.{E�<h�~���n=���a����������s�Q&��:+��[[!�6~H��n������t���������4��6����w���k�~PF�����<��:�'�p�^}�6��Tq\�0�9�AX������E��۞����(���a���߯��ο �还F���%�W9����?����濘K̿�Z�����_]`���'��   �   ���1Yd����£�d�V�`VW�������_@f�#��1���!�+�]�
����>��Q|����ſEGп��ӿr�Ͽ�Ŀ� ��6���.���g�Z���)�Ȯ������^d�����ƣ�ʖV��TW�:�����{;f����\�����+�"]�����<��Dy��u�ſ�Cп&�ӿ�Ͽ��Ŀ����a�������5�Z���)�x����   �   ��p��x����j\�2�9��Y����^�E�fޞ����b�(�_�a�%���᯿�οV��<J���'�P;�{������v�濯N̿z]��U���)a`���'��r��V��pE�am�z����n=��|a����������s�3"���%���W!�zH�n������q���������!��C���Au���k�2LF���6���谾�   �   ��Y���L�R���*2�ŋ�����*��
ϾU�CV����?γ��2ڿ����������!%�+�'�\�$�h��K������i�ؿ����(q��q�U���� Ͼ�%��x���A���k8�H����T�����]�N�k��-��g޾+���'���@��T�0`�Yd��v_��R��?�P+&�sN
�GQ۾����ڰg��   �   ���l\$�H7���Ϋ�BJ<��̽�}A��9��� � K<��K���g��
�׿�|�Z����,��P=�T#H�R�K�RG��B<���+�>��e��]�ֿP���D��B�<��� ��C����C���нd�D����:��J�/�۲��&�
�#}O�>���/���-M߾�W�`<�����D�zG�� �ɋܾ�Ĵ���+�J�� ��   �   �м�k{����:��P���R�2��D6j�n�ľ��y�]��@��Nǿ]���W��x1�akJ��n_�ۅm�FHr���l�Kp^�/jI���0���pZ���<ǿ����`�^�����ƾafm�m��]���{� �����ۻ��鼖.����޽��$�-]�������ĵ�����;�ž�0��nX��֞��F⇾X�X��v ���ֽ.v��   �    �T<�N�<�<(w��un�j��1���zS��.�&{��h���)߿���u�)���H���f�Vt���K��3X��X��:��#Df��_H�v�)��	���	Q����|�\�/�������d��R{�0�8�`b<d2�<P-"<X�9�z(�v���ҿ齲��G<��dV�
g��]l�o�e�H4T��9�D �8��V���s�0c��   �   �,=~�#=���<@�λ�J���� �����I���;�>���2N���������8�G
\�b%��َ�E������"��������pU\��]9��R���󿮸���@����@�O���]��B�$��}��ذ�8ʿ<O=D�= S�<���;0F��6�?�3���}2Ľ10齚= �v���������XR��+<���43� l��`�;t��<�   �   $6\=^�L=�|=�:���s��@�+��3��qN��I��Y��u�ÿ4���v5���B��i�D͇�Ş��=�����g��)��������i�T�C��U �' ��ſϑ�F	L�E����/?0��&���q��^�<
M@=*�O=�4=���<�M@< ����=�F�v���������l��:Bp��5�|bռ�齻��p<�=��@=�   �   j߇=�{=2�1=9�;�T������&�d7����r��F�����1�F!S�s,t�d|��{^��Z���c��������t�^T�� 3��`�ڶ�ڏ�������9� ��ؾ���,�k�`�#;�X=��g=F�{=.Ji=��;=�~�<�hf< ������̇�f
�^�Nu��׼HGf�@Ϡ:�<�<�=~*O=X�|=�   �   Re}=�+o=z+=���;��N��o��	���}�&�3�Y{���~��o�忂��^�.��LO�#]o������,������&��������o��P���/����u���t��&��nc6�M�������J�d��O;D=�Z[=v�i=�P=$+=Xn�<@|3;�]}��a�x�4�ƦT� �]���O�d�+�d��P3@��;�;���<ƌ/=<0d=�   �   7E=69I=4r=���;�r>�A���X����۾��)�>�u�᧿T�ڿ���_8&��hD�P�a��{��,���1������z�Z�a��D��&�ܾ	��]ܿln���ex��@,���߾���. �N�R� ��:� =��5=�1=��=`!k<�����Od�����m^��L5ӽ!}ٽ��н u��&+���S�X�⼀�V�l,�<�^=�   �   @��<r�=���< �;�)'�^���i�� ǾJ��0�`��L���ɿ����;�_ 4�ʚM��Kc���q�E�v�fqq�e�b��L���3�
 ��e���ʿ{L���b��s�#ʾ�Fo�ɣ��9� X�9(v�<�x�<�Š< �J9�jݼ�r�xc��%���) ���7���F��gK�cGE��
5��A��q���T����]��#���$�;�   �   �1���<0�`<�:ڋ�pȽ`�H������Y�z F��Ԉ�N���H��R�������5��bG�h,S��W�Z�R�}fF�v�4��6�f2�^�Ύݳ�E���5G�y�a����L�+Vн�'� +Z�(6<�ޓ;�j}�\SB�5{��!+�?>���o�>���u���c��)ӭ�Wq��ޱ������*�j�+w8��k��{����-��   �   �q��ȼ@�λ��黸 �������#����L���'���i��k��Y�¿|9�[
���1O*��3�,�6�q�2��=)����	���)¿���k�i�(��$�xY����&�����8m���*�l"�X/��8���F罭�1��ox��7��"6ž3��H��a�(�	�pm�����0����Ɲ��q�}�+�G�ܽ�   �   ������i	��៼HL�`l|�\����a�������]�?� O�,/��OTſs���2�x���#��v�ǎ�����_���ÿd���,�}��>����A���b� � �'� (���������%@��;��e�K��f���kľʯ�����,���=�c�H��L���G��<�:$*����|������O���F��   �   �iN��@�������� ���d�@��P���S(�Z~��ѨҾ��^@J�[���r���DQ��Ǆҿ�L�M񿒼��𿾟� �п�Y�������I��<vH�����QѾ�҉���'�$պ��D��=���� �<⑽/��p�R�d#����ھ����63�xU���s�����\݌�O.��ZN������Wq���R�	�0�%s�-2׾Y���   �   o����C��z�$�{�tw�����.�U����E�SE��-�߾�����E��Nt��X��5ƣ�]Ҳ�S6���)���w��M���#������Nq��pC����h"ݾ�k���C��t���{��u�֌��6����F��H����߾����E�FSt��[��ɣ�yղ��9��-��{��Q����&�����fRq�tC�c���&ݾ�   �   QUѾ0Չ��'��غ�VD��:���� ��ܑ����m�R�S��c�ھ=���23��sU���s�����ڌ�r+���K�����uq�V�R�N�0�p�B-׾XU��5dN��8�����Ј�l���z�@�<U���W(�5���լҾ@!��CJ�x���񦞿T���ҿ�O���&�����
���п>\������K��gyH�K���   �   }�������b�� �����@'���촼���W9��_��͉K��b���fľX���0���,�(�=���H�L���G�|<�/ *�j��_y������O���F��	������|a	�۟��M异q|�0a����a������!�9�?��R�^1���Vſk�濐4�G���%��x�������]�+��S�ÿl��{�}���>��   �   �(�s'�A[��Я&������m���*�hQ"�8�:1��<��1��gx��2��R0ž�,��A����i�	��i������*�x���M�����q�J�+�ǜܽ�q��ȼ�lλ��������v�#����l���'�Z�i��m����¿	<��	
����Q*��3�8�6�j�2��?)�H��h	�`��$¿v���i��   �   �7G�Oz�����L�;Xнj(�@Z��I<��;=}� DB�\q��%��7>��o�s���p��D^���ͭ��k��Ƭ������wj�(p8�
f��r��d�-��0��<��`< N:��sȽ��H�����p[��"F��Ո�󬳿G�ῃ��j��0�5��dG�s.S��W�Z�R�LhF�
�4��7�}3�*��߳�=F���   �   N�b��t�zʾNHo�������9� ��9�|�<T��<�ՠ< �U9�Nݼyr�LY��?��"# ���7�9�F�]`K��?E��5�[;�Zf���J��̼]��	�� u�;ܟ�<J�=���< �;,'���p�i��Ǿ�����`��M��y�ɿ����C��4�K�M��Mc���q�5�v�Asq��b���L���3�� �g��5�ʿgM���   �   �fx�:A,���߾����� ���R����:J#=X�5=b�1=��=�Dk<��D��
Ad�t�U��,ӽ�sٽ��нUl��7#����S��⼠�U��<�<�d=�;E=2<I=�s=P��;u>�_���Y����۾��)���u��᧿_�ڿd��(9&��iD�~�a�{�v-��p2�����_�z�j�a��D���&�_�	�g^ܿo���   �   V���c6����$�����6�d�`Z;�=�\[=:�i=v�P=�/=y�< �3;�@}��Y�޽4�ڝT��]���O��+�<��`@� j�;L��<��/=*3d=~g}=$-o=�+=���;��N�\p�*
���~�¸3��{��C��������.�oMO��]o� ���-��}���B'�����R�o�kP�<�/�������Bu���   �   쀅�_�9�ө򾞾��{,�2k���#;,Y=t�g=��{=�Ji=��;=��<jf<��� ��� ��,
��]�Hu��׼PGf� Π:�<�<�=@*O=$�|=I߇=��{=Ȑ1=@4�;�T�V��:���&7����r��,F����1�\!S��,t�n|��^��Z���c��|�����t�FT�� 3��`���뿹����   �   ����b6�`��M���ʉ�N�d�@y;�=V][=��i=؃P=�/=xy�<`�3;�@}��Y�ڽ4�ԝT��]��O��+�@��h@�`j�;l��<��/=b3d=�g}=�-o= +=��;��N�Do�[	��`}��3�-{���~����K���.�xLO��\o�H���H,������r&��Z����o�hP�q�/�6�����zt���   �   {dx��?,�!�߾������B�R��f�:�%=��5=n�1=`�=�Fk<������@d�j�U��	,ӽ�sٽ��н\l��;#����S���� �U�4=�<@e=�<E=z=I=�u= �;�o>�R��4X����۾:�)�Z�u�m৿��ڿD���7&��gD�I�a�e{�,���0��%����z�$�a��D�2�&�2�	��\ܿ�m���   �   !�b��r�4	ʾ�Co������9� �9���<���<�ؠ< �V9�Mݼ|xr�"Y��0��# ���7�<�F�c`K�@E�5�^;�`f���J����]�P	��z�;$��<4�=���<P�;�$'�b��"�i�b�ƾO����`��K���ɿd���Y�B�3�l�M�!Jc�$�q�W�v��oq���b���L�G�3����c����ʿUK���   �   �3G��w�$�����L�@Qн0� �Y��Y<�3�;86}��BB��p���$��7>���o�p���p��E^���ͭ��k��ˬ��	����wj�'p8�f�wr����-���0��<��`<��:D��;lȽۉH�͍���X��F��ӈ�橳����A�������5��`G�l*S�rW�P�R��dF�΋4�&5�11�X�� ܳ��C���   �   �(�|!�W��&�&�I什�c�(y*�@"���N0���;���1�agx��2��G0ž|,徿A����l�	��i������*�{���O�����q�/�+�e�ܽ��q���Ǽ@Mλ �黴���f����#��������'��i�^j��h�¿%7��
����bM*�$�3�#�6�r�2��;)�����	�r���¿����i��   �   ^�����E�b�f� �[���Tߴ�n���7����~�K�mb��~fľH���)���,�(�=���H�L���G�<�2 *�l��`y������D���F�	�������]	�`Ο�8:弐b|��U��r�a��򵾲��?��K�&-���Qſ���P1�����!��t���<��#�l��T�ÿ1�����}�4�>��   �   �MѾ�ω�:�'�κ��D�L'���� ��ڑ�L�� �R�.��I�ھ3���23��sU���s�����ڌ�u+���K�����yq�Z�R�P�0�p�;-׾CU���cN��7��� ���������4�@��J���O(��{���Ҿ�.=J�c�������N����ҿAI��������d���п�V��L����G���rH����   �   &h����C��l潈�{�$j�$��$)�w��R�E�#E���߾�����E��Nt��X��4ƣ�]Ҳ�T6���)���w��O���#������Nq��pC����Z"ݾ�k����C�Ns�^�{�Dm���:#�߂���E��A����߾��\�E�_Jt�xV��hã�Uϲ�&3���&���t��;|��� ������Iq��lC�i���ݾ�   �   �]N�T/��H����|�������@�,N��.S(�~����Ҿ��S@J�V���n���AQ��Ǆҿ�L�P񿖼�����п�Y�������I��:vH�����QѾu҉��'��Һ�	D� '��� �֑������R�t��a�ھ���.3�(oU���s�Y����׌��(���H��R���xq�ۻR�h�0��l��'׾5Q���   �   R���갋��T	�$ş��8��e|� Z����a�k�����S�?�O�(/��LTſr���2�x���#��v�Ɏ�����b���ÿf���.�}��>��������b�� �����Hٴ�8���1�����n�K�p^��saľ#������z,���=� �H�XL�E�G�<�*����s��9�����F��   �   ��q���ǼPλ`�����P����#����&㾷�'�{�i��k��X�¿z9�Z
���1O*��3�.�6�s�2��=)����	���,¿���m�i�(��$�CY���&�M򧽆e�@r*��*"���s)��t2罡�1��_x�.���*ž&&��:�����	�f�����3$�����c���v�q���+�=�ܽ�   �   ��0��8<a<�E:��%nȽċH�^����Y�r F��Ԉ�M���H��Q�������5��bG�j,S��W�\�R�}fF�x�4��6�g2�`�΅ݳ�E���5G�y�>���b�L�OTн�!�`�Y�Ph<j�;P}��4B��g����0>���o����sk���X��1ȭ��f������O����oj��h8��_��h����-��   �   0��<��=���<`�;b%'���콬�i�� ǾB��,�`��L���ɿ����:�] 4�ʚM��Kc���q�D�v�fqq�f�b��L���3� ��e��	�ʿ}L���b��s�ʾHFo�z�����9� ~�9H��<��<�< �`9�3ݼ�hr�qO������ ���7��F��XK��8E���4��4��Z���@���]���pϧ;�   �   �AE=.AI= x=`�;"p>�Ԃ��X��s�۾��)�;�u�᧿R�ڿ���_8&��hD�P�a��{��,���1������z�Y�a�	�D��&�ܾ	��]ܿmn���ex��@,���߾ꎅ�����R��X�:�&=��5=Ԡ1=z�=�fk<������2d��朽�L��#ӽ�jٽm�н�c��5����S��� <U��N�<l=�   �   �j}=�/o=^+= ��;��N�go��	���}�"�3�Y{���~��p�忁��_�.��LO�!]o������,������&��������o��P���/����w���t��&��nc6�H��階�����d�`o;&=r^[=��i=��P=�3=���<�<4;p&}��R�ص4�d�T�`�]�X�O��+������?����;���<�/=�6d=�   �   ʚ=c��=�7a=��<8��������i��DɾH���d��i��4H̿� � �ݧ6��Q�&�g��w�G�|�b$w�(�g�O�Q�p{7�u1��-���οxr��y�g����3Rξ�r���x��E}< �A=CՁ=tڊ=2��=��\=�n&=���<(`:<���X9�����5��4퀼�����:;|�<l�=6�B=�D{=.L�=�   �   ���=�'�=6<[=(k�<�{꼉�ܽ��d��5ž ����_��ʙ���ȿ������N�3��DM��1c�' r�iw�r��Bc���M��64�9��.��˿�����Kc�����ʾ]Nm���������|<�=<=��x=Ҽ�=�o=��@=�=P��< �D�Њj�t�μ~����	��\���ӵ�0�#���;��<�5 =\�^=I2�=�   �   ,�r=�v= �H=�M�<�Qμp{˽ՙU��p��Pj��FT�q$��b��i&�z_�a�*�KxB���V�8d�~�h�b�c��JV�PhB���*������������fW�L��췽��Z]�ڽ&��p�v<F�*=B�W=��S=n�+=؂�< ��;tw�~���]�����坽碽+~��<q���NK�����p��`�W< a=�{J=�   �   �?=jk:=��&=�٥<`b��7J���F>�6#����w�A���;����ݿ#��	��42�F�C��RO�8ES�b�N��C���1����'�|&޿������"�C����2�����D�����ټ`�a<td=��= c�<x�[<�q/�? ��΍���ɽ�����#� ��$�b	� z����#����#��
�`,]� �<�   �   �;�;̯�<X~�<���<y�񓑽�5!���2��[*�*6m�泜�7�ſN��,��[��!-��6� �9��86��K,�}��c����ſ 䜿un��y+����ď���D&�D�������.<$�<t��< &����(B��!�ڽ��X�E��Bl��>����������}����-��f�f��>�)��"T˽(Nl�T���   �   �-�8����%<8@<�7�*{`�4>���l������u�I��D��,P��cϿ�򿾙�1�����&:�_)��������B𿥩Ϳԁ��Pꅿ*�I�	�8���o�ȷ�p�p"}��?�;�;`�>��:/�,ⰽ�L�,M������}��^v¾�^ؾM �e�?�侼�վ���W���悾�E�`��k����   �   �����7�h�j��K����*"��e½l�7�������羦�$��]�q5�� }��OEʿ�_�Q���Y��p���6�����F��Gȿ�ު�����[���#��I�����%9��$ƽ�),��4P�pK���d��`L�[ɽ��%�>�s�Yԥ�[�Ӿ.	 �@���#�=�,�;�/���+���!�^��hn����ξ�k���l�ڴ��   �   �R&����L�;��4����>�P.ݼ�B���De��򱾲N ��:.���`����|����;��(�ȿ,KӿȊֿjҿbXǿ�W��7Ҡ�5q���]��_,��$���n��d�c�b;�B���D��p'[��>����H���Ƚ �+��J���X���{����k58���R�ܐg���t��x��ms���e�J@P��i5�Q����I������   �   ��|��%��D�� �"�(F��$H���3'��L���1 �x���������:r*�vuS���z�����.��^��o���C�����������{w��gP���'�k� �`����|��!��?����"�C���L��\:'��R��E6 �����򩽾����u*��yS�.�z�D����	���`��V������WĚ�$��L�w��kP���'�� �B����   �   ,r��٫c�R>�����h�� "[�|4��h�H�)�Ƚޚ+�%G���S���u��S �f18��R��g���t�֑x��hs�@�e��;P��e5��M�x��E������M&�)���Ơ;�T,����>�`5ݼ�������Ie�n���Q ��=.�~�`�������>��,�ȿONӿ��ֿ0mҿO[ǿ{Z���Ԡ�Ks����]��b,�=)���   �   M�r���)9��(ƽ�,,��3P�P,��@U��TL���Ƚ8�%���s��ϥ���Ӿ� �����#��,��/���+���!�΢�h��{�ξ&g���l�y������7�phj�`�P��/"�-j½
8�a���m��(�$��]�g7��o���Gʿpb�x��� ����8�����I�oJȿ�િ�����[�=�#��   �   �
�o:���o�����p�($}��T�;��;�>�p-/�*ٰ��F��$M�w����x���p¾|Xؾ�澊^���侪�վ��p����Ⴞ�
E�������T!�0���؟%<pG<��7�(�`��@�`�l�<��ȱ���I�eF��R���Ͽ��4�����[���;�+�:����RE𿾫Ϳ�����녿h�I��   �   b{+�$��6����F&����P����.<�	�<���< ��p��u9��]zڽr�֗E�::l�	:��ְ����������5)��:�f���>�����I˽�=l�f��`��;\��<`��<���<�	y������7!�����4澶]*��8m�]�����ſd��b�V]��#-���6���9��:6�M,�U~�e����F�ſH圿|n��   �   ]�C����a����D�����ټ��a<tg=��=|q�<�[<�@/��/ ��ō�F�ɽh������� �h�$����s�ϻ��)���������t\� �<F=�o:=��&=ڥ<�f���L���H>��$�����A���=<���ݿ��
��52���C�:TO��FS���N�'C���1�����'��'޿�������   �   9W���������[]�ڽ���H�v<X�*=��W=j�S=��+=���< ��;�Fw�h����]����ܝ��ޢ�v���i���@K�о��@]���W<Vh=��J=J�r=bv=F�H=PM�<�Uμ]}˽l�U�*r��.k�HT�2%��mc���'�%`�,�*�<yB���V�cd���h���c��KV�,iB���*������Z��������   �   Lc����ʾ�Nm�Ț����P�|<�><=��x=��=�!o=��@=��=���< �>�hnj�4�μ�����	�M���ĵ��#��I�;��<(: =� _=�3�=���=t(�=�<[=Hj�<�~�ԿܽǺd�U6ž���7 `�˙�8�ȿ�������č3�SEM��2c�� r��iw��r�QCc��M��64�~�����h˿߮���   �   F�g�����Qξ��r�1󽮛�0G}<r�A=rՁ=�ڊ=a��=��\=o&=���<8a:< ���9�����`5��퀼��� �:;t�<\�=&�B=�D{=L�=�ɚ=C��=<7a=��<č��-��(�i��Dɾt���d��i��VH̿� �' ��6�Q�4�g��w�I�|�[$w��g�@�Q�^{7�d1��-���οYr���   �   	Kc� ���ʾ0Mm�ɘ�X��@�|<@<=h�x=T��=2"o=�@=�=���< l>�nj��μ�����	�M���ĵ�0�#��I�;�<2: =� _=�3�=Ê�=�(�=�=[=�m�<|y��ܽZ�d�E5ž���0�_�kʙ�b�ȿ����Z����3�^DM�m1c��r�khw�gr�*Bc��M�&64�ш��
���˿-����   �   /W�d�������X]�Rڽ�����v<��*=�W=��S=t�+=���<p��;@Ew�6��f�]����ܝ��ޢ�v���i���@K�Ծ���\��W<�h=�J=�r=�v=2�H=�S�<Lμ�y˽��U�$p���i�FT��#���a���%��^���*�xwB���V�d�P�h�6�c��IV�YgB�*�*�G��ڎ����X����   �   ��C��������,�D������ټXb<�j=��=ht�<@�[<�=/�\/ ��ō��ɽI������� �k�$����s�ջ��'��������@n\� �<G=�q:=��&=��<XY���G��,E>��!����F�A�Q���9��H�ݿ`����32���C�HQO��CS���N�mC�S�1����+&��$޿�������   �   x+�B��ˍ���A&�����t��@�.<,�<��< D�����9��zڽR���E�,:l�:��հ������Ę��8)��=�f���>�����I˽r=l��d�� ��;x��<��<��<�x�v���_3!�t���/�pZ*�24m�������ſq����Z�� -�t�6�T�9�A76��I,��{��b�{���ſ�✿n��   �   �/5����o����:p���|� ��;�3�;ؒ>��+/�~ذ�|F��$M�e����x���p¾xXؾ�澋^���侮�վ��r����Ⴞ�
E�̕�������P⿻�%< ^<(�7�s`��;�,�l���:��A�I�gC��pN��Q Ͽ��\�������t8��'���B��I@�^�Ϳ����腿��I��   �   �E�/����!9�mƽ ,��P������L��HQL���Ƚ�%�~�s��ϥ���Ӿ� �����#��,��/���+���!�Ѣ� h��z�ξ!g���l�N��Z����7��Yj����s��!"�A`½��7�4���A��a�$��]��3���z���Bʿ�\�B������Ȼ�=5������C�WEȿ�ܪ����ҟ[�j�#��   �   Vk���c�V7�� �弈�Z��(��n�H���Ƚk�+��F���S���u��J �`18��R��g���t�ؑx��hs�D�e��;P��e5��M�v��E������M&����X�;�D!��Џ>��ݼ�톽����?e��ﱾ�L ��7.�B�`�k������8��:�ȿHӿ��ֿ gҿhUǿU���Ϡ�o��Y�]��\,� ���   �   ��|�
�@8��|�"��-���7��F.'��J��J1 �F���������0r*�puS���z�����.��^��r���F�����������{w��gP���'�i� �R�����|�!�5>����"��3���5��)'�F��q- �|���ơ�����	o*��qS��z�2���}��<[������h���뾚�!��Mww��cP�(�'��� �����   �   ^H&��}��t�;�8��0�>� ݼ����|��?De��򱾢N ��:.���`�~��x����;��'�ȿ,KӿɊֿjҿdXǿ�W��9Ҡ�6q���]��_,��$���n���c��:����ȣ�H�Z�� ��R�H�T�Ƚ��+��C���O��Ap�� ���-8���R�N�g��}t�Ȍx��cs�}�e��7P��a5�cJ�����@������   �   ������7�P:j��}�hp��$"��c½��7�}�����羚�$��]�n5��}��LEʿ�_�P���Z��q���6�����F��Gȿ�ު�����[���#��I���l%9�#ƽ�#,�`P��帻D@���FL�+�Ƚ��%���s�'˥�?�Ӿ� �����#���,���/���+�ρ!�.���a����ξ~b��H�k�����   �   ������@�%<�i<��7�bv`�n=�.�l�Z��֯�k�I��D��)P��`Ͽ�򿽙�2�����(:�`)��������B𿦩Ϳց��Rꅿ*�I�	��7����o����p��}����;0Y�;Hr>�|/�:а�A��M�9����s��k¾fRؾd�X�d�侊�վk��m����݂�}E��������   �   @��;���<Ȕ�<���<8�x����5!�����1��[*�%6m�峜�6�ſM��+��[��!-��6��9��86��K,�}��c����ſ䜿xn��y+��辡���9D&����������.<��<��< ���8���0���oڽ,���E�2l��5��$���⍑�����$����f��>����6?˽8,l��I���   �   6N=�v:=��&=,�<xZ���H���F>�#��y�r�A����:����ݿ#��	��42�F�C��RO�9ES�c�N��C���1����'�}&޿������"�C�������M�D�\��,�ټ b<�l=��=���< �[<`/�J! �'���4�ɽ���v�� �ڥ$�j���m�t����~��;�������[�,)�<�   �   ��r=�v=@�H=4U�<�Lμ�z˽��U��p��Jj��FT�p$��~b��j&�z_�`�*�KxB���V�8d�~�h�d�c��JV�RhB���*������������fW�J��߷��mZ]�Xڽ���8�v<��*=��W=b�S=Խ+=ȡ�<��;�w�����]�/닽�ԝ��֢�n���a��r2K�\����0�pX<Rp=2�J=�   �   틒=�)�=�>[=�n�<,y�+�ܽ��d��5ž��~�_��ʙ���ȿ������M�3��DM��1c�& r�iw�r��Bc���M��64�9��1��˿�����Kc�����ʾENm�(������|<L@<=f�x=9��=�$o=2�@=*�=̦�< �8�8Tj��μ���	��=��@���|#��z�;�#�<�> =�_=?5�=�   �   ���=x˧=�Ɋ=��#=�»'����f4�졾�� �h�=��x��<���V�ٿa��gS��4/���@��-L��HP��2L�b�@��/�T��ؔ��zۿ�ݮ��H��A��������>?�C��������P�<@gc=e�=���=փ�=��z=4�L=�=<��<8t<0p�; �;��:@?�;�6<Ľ�<��	=:�A=��y=��=d8�=�   �   Xx�=�ڢ=J�=ֵ"=���������/�E������<W:�J5�����Wֿv������>,�i%=�)pH��fL�hH��0=�n},�JQ�m^�d�׿۫�e傿aw=��A��㣾?~:�P���$g��4}�<��^=Y�=G��=��=��b= /=@�<(�~<��x;�����+��=�H���|^��%<x��<4=�[=���=B|�=�   �   �F�=k��=�e=��=�A	��%��&B#����.H�0P0��6u�fȡ�1�˿�������#��o3���=��eA���=��@3�<�#�w��r���;Ϳ^����w�<�2��?��]����,�n֚���H��z�<��P=r�v=��r=�dP=Nf=��<�0;خv�x����,���I���P�*�@����ż0�什�C<��<��G=~Ā=�   �   ��W=��r=�sa=�= ��:�Nb����~#��ߤ׾]� �}r`������뻿���+R�F��B�$���-���0�,�-�lE$�~O�����e��&g��=9b��|"�~۾i��ζ�n^�������<��6=�E= �)=@��<�\�;4Ӗ�>4�q���K4���۽��4���3�v�ҽ����x�X�(��\O�<�=�   �   lA�<�%=�3=0�=�h�;�-�7Wc���f����E��ă�%G��/t˿��h�=���`���������O���;�ʿ���+�F�������i�����MI���غ`\�<�=�<�u<p�zX&��ʛ�A�罁���89��R��Tb�M�f���_��M��Q2��*��jԽ$�W��@��:�   �   �D�P�i<���<�!�<@�<8O�kC���7�E������0�'���`������N����Ϳ�.�@���+��(�.��q������E̿?+��r؎�2`��v'�\t쾱뛾[e;�����W
��jH;L�<�פ<pS�;�e��j�o�ۘսP_��CV������]���ԯ�`���ܾ������U����>���ZL������&H��   �   ��v������;��<(v%<�	��!��+[�&�r�⫼�����8���l�>p���4��0���4Bӿ�6޿�ῄ`ݿ��ѿ=������x��оj���6���c����r����M톽�N��P��;�>< ��9LKۼⵋ�����"@�A����{�Ѿ]����@��NQ������f��0�̾jܦ����8c6�{���   �   ������~��櫼�);h�<���8��j���+`2�Y
����ѾB�-;�?~g�����F������l	��'ܵ�,L��J���b���7Q���{d���8�;9�vLϾvT��}g0�0?��<N!��U߻ 7�;��i���мj����(��O�"���3�Ⱦ���� ���f/�##A�?=L���O�08K�!??���,�����U���þ?��,�G��   �   &pE���x�_��S����; 5�:@����j�����J�m-���:־f���/���Q��_o��8��6m�����`Ή�����zl�ϖN���,�5S
��Ѿʕ�HkE�-轀�_��I����; ��:8K��Ρj����+�J��0��9?־H��|�/���Q��co�;���o�������Љ�H���~l���N��-��U
�l�ѾT͕��   �   0W��Rk0�9D��$T!��h߻@?�; uh�<�м$����$�ޓO�6���J�Ⱦ��������b/��A��8L�P�O��3K�;?�E�,�I��.P��q�þ�����G������~��׫�`A);h�< ��������`d2�Q����Ѿ��b";��g�����������#���޵��N��Ը������LS��hd���8��;�(PϾ�   �   B����r�l�������T�����;�>< 5�9 7ۼ���������@�=��L���Ѿ󾍙�����M�J����S����̾�צ����:]6�:����v�	��0�;���<�t%<P���$��8^���r��������8�.�l�<r��A7�������Dӿv9޿®�Lcݿ}�ѿ���؅��V����j���6����   �   6w쾵훾h;����Z
� bH;��<��<���;�N���o��ս%Y�*<V������X��zϯ��Z���־�U���������:��eSL������,H�p�C��j<���<%�<Њ<�W�`G��3�7��������U�'�o�`�X����P��5�ͿF1�������C*���������`̿-���َ��4`��x'��   �   ��������i�(����PI��	ٺ_�<t�=+�<6u<���I&�����;�����19�(�R��Lb��f���_�K�M��J2��$�V`ԽT憽|;�� �:�Q�<H%=>�3=�=�[�;>-��:Zc��ﺾ����E��Ń��H���u˿��3i����b�
����@��g������ʿ:��I���=�F��   �   �}"��۾l�����_��0뻠��<�6=&�E=B�)=��<���;`�����3�����b*��B�۽���Ԓ���'��ҽ@���R�w�JI��t�Pc�<�=XX=��r=�ua=6	= ^�:�Rb�h���$��Ȧ׾�� �4t`�����2�g��S�C��[�$���-�(�0�R�-�yF$�mP�R��%f��h���:b��   �   ��2��@�^����,�Tך�0�H��{�<V�P=:�v=��r=LjP=m=h-�<��;؁v�|�����,��I���P�L�@�~����ļ ����C<���<��G=�ƀ=�H�=���=�f=l�= [	�Q'���C#�$����I�2Q0�.8u�5ɡ�)�˿������޿#��p3���=��fA���=�|A3��#�
��c���Ϳ�����w��   �   �w=��A��㣾�~:�����,g��~�<��^=AZ�=S��=#�=*�b=D/=�I�<��~< Yy; K���+�xq=�x�� �\���%<���<�8=��[=��=l}�=:y�=ۢ=r�=��"= ���&���y�/�쀞������W:��5������ֿɧ�(��X?,��%=��pH�BgL��hH�1=��},��Q��^���׿U۫��傿�   �   �A�b��΅���>?�͜��x����Q�<�gc=��=%��=��=4�z=��L=H=���<pt<�r�; �;��:@�;�6<ܽ�<��	=<�A=��y=��=N8�=���=^˧=�Ɋ=�#=`�»����&g4�M졾�� ���=�y��Y���t�ٿq��vS��4/���@��-L��HP�|2L�Z�@��/�F��ɔ�ezۿ�ݮ��H���   �   �v=�FA��⣾A}:�����pb��T��<��^=�Z�=���=b�=��b=�/=\J�<P�~< [y;`J��Ȗ+�`q=�`�� �\���%<���<�8=��[=-��=�}�=ey�=lۢ=��=�"=��������A�/���������V:�5��D��ֿB������>,�%=��oH�IfL��gH�;0=��|,��P�^���׿�ګ� 傿�   �   3�2�5>�\��.�,�Ԛ��H�ā�<z�P=Ƴv=��r=(kP=�m=p.�<��;��v�����p�,�ĺI�n�P�D�@�p����ļЌ�p�C<$��<<�G=5ǀ=I�=*��=�h=(�=�	�)$��+A#�k���3GO0��5u��ǡ�x�˿���q��x�#�,o3���=�eA�ۧ=��?3�x�#����F���?Ϳ���n�w��   �   J{"�|۾�	�����2[�����(��<��6=H�E=ʘ)=
�< ��;ܷ��H�3�T���2*��%�۽���ʒ���'��ҽ:���D�w�,I��s� d�<X=`X=*�r=8xa== �:(Jb�*��n"��`�׾U� �q`�̧���껿���dQ�_��:�$���-���0��-�QD$�}N���4俲c��f��z7b��   �   ��}}���i�����EI��غti�<�=0�<h=u<����H&�#��������m19��R��Lb��f���_�L�M��J2��$�H`Խ@憽�:��@�:�S�<%=2�3=��=0��;�-�3��Tc��뺾����E��Ã��E���r˿���f���{_�Y��|�����&�����j�ʿK���탿r�F��   �   q�6雾�a;�a���N
���H;�!�<��< ��;�J����o�X�ս�X��;V�����X��sϯ��Z���־�T���������:��^SL���i��nH���C��j<��</�< �<�@��>���7�2������K�'�G�`�/����L���Ϳs,迬�����o'�ɝ����
��
̿G)���֎�N/`��t'��   �   ����r����熽(<��`�;��>< /�9d1ۼ��������f@��<��5��ұѾ	󾉙�����M�J����U����̾�צ����"]6���轺�v���07�;���<��%<���N��X�ۖr��������[8���l�cn���2��ɿ���?ӿ�3޿�Ό]ݿ.�ѿ���n���{��l�j�8�6�{��   �   YQ���b0�'8��,C!��
߻��;�g���мϜ��$���O����-�Ⱦ��������b/��A��8L�S�O��3K�;?�G�,�J��-P��n�þ���c�G�����~��ѫ���);8�<�������8���\2����"�Ѿ��,;��zg������������nٵ�}I����������O��xd�d�8��6�`HϾ�   �   �eE����~�_��4��@7; "�:�5����j�c��{�J�D-��z:־Y����/���Q�_o��8��6m�����aΉ�����zl�іN���,�5S
��Ѿ�ɕ�kE�S�ƭ_��@��@; >�:<-��H�j����šJ�
*��76־�����/�̪Q�8[o�b6���j�������ˉ����Svl�ޒN�&�,�VP
�t�Ѿ`ƕ��   �   ����$�~����� �);X�<�Ͱ��������_2�+
����Ѿ4�";�6~g�����C������k	��)ܵ�.L��L���c���9Q���{d���8�89�mLϾ_T��&g0�>��ZJ!�P&߻p�; Cf��мN��� ��O�s�����ȾN���a��_/��A��4L���O��/K��6?�}�,����SJ����þ���V�G��   �   �v�� n�;��<8�%<����D���Z���r���������8���l�:p���4��/���2Bӿ�6޿�Ὲ`ݿ��ѿ>������z��оj���6���Q����r�?���놽�D��`��;��>< ܟ9�ۼ������~@�99�����x�Ѿ��8��.��!J����@�$��P�̾Ӧ����V6����   �   x�C��=j<���<4�<(�<dF��A����7����m��%�'���`������N����Ϳ�.�@���,��(�/��t������G̿?+��r؎�2`��v'�Tt쾚뛾e;����|S
���H;T$�<x�<`�;D6����o�'�սS��4V�[���"T��Nʯ�U��]Ѿ��繾���Ր��L6��LL��
����
H��   �   de�<L%=�3=` 	=P��;�-��5�CWc�d�Z����E��ă�#G��.t˿��h�>���`�������	��P���=�ʿ���,�F��������i�%���|JI�@Wغ8j�<��=<:�<8\u<h���:&�����u�����*9���R��Db���f�{�_���M��C2�@�jUԽ%݆�4���z�:�   �   �X=��r=�za=.=��:xLb�N��\#��Ȥ׾T� �wr`������뻿���+R�F��B�$���-���0�.�-�lE$��O�����e��'g��?9b��|"��}۾U��|��Z]��P�����<��6=��E=&�)=��< �;؟����3�㋌�� ��Ħ۽��𽜇����`{ҽ����w�:��@��x�<�=�   �   K�=���=tj=�=@	��$���A#����!H�+P0��6u�dȡ�2�˿������ �#��o3���=��eA���=��@3�=�#�x��o���=Ϳ]����w�<�2��?��]����,��՚�P�H���<R�P=еv=s=�oP=�s=�=�<@e;�Vv�L�����,�4�I���P���@�\��d�ļp5仐D<\�<�G=�ɀ=�   �   lz�=)ܢ=o�=|�"=��������|�/�<������<W:�I5�����Vֿv������>,�j%=�)pH��fL�hH��0=�o},�JQ�m^�b�׿۫�f傿bw=��A��㣾(~:����e��P��<��^=[�=]��=m�=R�b=	/=�R�<��~<��y;`��X}+�PW=�Xo��T[���%<x��<:==��[=җ�=�~�=�   �   X{�=릾=�ť= Aj=,�<�_$�����&uu�K�ɾ�^��mT�b��п��[-ٿ�:������2�� &��)�x&��I�L�B���aڿ�.�����B�W�v~��%оaS����c�@X�:�W=�z=&�=�D�=���=2�=�ji=>�A=��=<��<�g�<�˫<��<��<��<0#=`?P=�ˀ=�M�=n�=��=�   �   .4�=�Y�=|`�=�Vi=D��<�!����%�o�a�žʄ���P�����ϯ��տ�&��qn�8��f/#�;+&�w)#�!��������ֿ�������S��z���˾|�|��	��>Y���(;��=�v=ex�=;��=pь=�y=��P=�c$=`m�<�֩<��f<��+<�)<p�a<h-�<(��<�-=Zoc=`}�=q��=ܗ�=�   �   N�=�-�=^�=�f=���<�����m�_��߹�n;��E�j����:���{˿J�?������|��������������̿ ���Ą�|�G�m��U+��(k�����M=����;��=�(l=tg�=Ɍ�=h]j=R�<=@ =\*�<��; �������#��lո�(����	)� N�:��<d=6�J=�S�= !�=�   �   B1�=�g�= ��=�^=@#�<(3¼����U�F�6Y��ʈ��BP4�GOq����� m����ۿ)A���k�h��f�v��������bۿy������r�J�5��Ɔ��eP�8�׽z��X�-<�G=��X=�c=�K=��=t[�< 9�9H���[$�,gk�YՐ��򠽊Z��x���`��j�E�0����ǻɆ<H�=��b=�   �   z_6=��i=6Qu=v]P=�f�<��X�����z�&�>ݏ�ލݾ 7�b U�ON���æ�y�ÿ�pݿ�}�7���2�Ψ����sܿ�	ÿ�E���'��xHU�P����߾����)�-�@(��p��芁<z�=�"9=x`)=�1�< ��;DF����@�NV��s�ٽ�1��t���'�n+�C�$��4��,��z�½E����@��0�<�   �   �yR<@[=��<=�F8=$�<`��X\��P�8�j�T��	(�[�4�h�h�
��ن��N྿Gп�;ۿ��޿8�ڿ�1Ͽԝ��"Z��\!����g�f%4��������m�����Ft�� ��~�<��= �
=X��<������A����潞���1K�t~q�����P萾@����K��w����zh��?������ɽ��d��h���   �   `���>�;8��<�=T��<�+<p�����8z4��ő��)־a�� �>�;�k�薋�|����O��`���L~��굿)0���2��o7��Q�i���<����1�Ծ=����4�1[��G� E;�)�<��<���<�����4"�>w����o�J���\ϣ�����_Ծ(������߾ Ѿ�x��8@����}��=�� �xC���   �   ����O���>�;��<d��<��<�(J�Bq��
 �c�X�釣����'��GZ:�{�]�Z�|�����5��n���i������HBz���Z�
�7�e0�>&�̞��^�T�����r�l�p�Q���e<���<<�<�P3��x�ɇ�����_Be��z��xȾ�M�z��t}��#��{&��"����s	����Y¾(���6�Y��Z��   �   ���啽@�ɼ %�;4}�<��<���;8��6�������]j�[���޾�V�A(���@��%T�k1`���c��"_�0R�7W>�d%�rx	�V�پ�����-b����ߕ� �ɼ�G�;��<�ݰ<י;(��E���"���cj��^����޾�Y�jD(�M�@��)T��5`��c�'_��3R��Z>�Cg%�({	�ғپ6���V3b��   �   ��T�`����l���Q���e<���< �<��2�jn���������;e��v���ȾKH�M��z�O�#�x&�V�"����pp	��쾴¾R����Y�<V�����l;���q�;��<���<�݃<P>J�6Kq�: �@Y�5��� ��Ή�u]:�'�]�o�|�����d7����������5���4Fz�*�Z��7��2�8*�ڡ���   �   ���W�4��_���L�@�D;L)�<��<���<�W���("�8o������J�(���ʣ�v��=ZԾH�����߾�Ѿ�s���;���}�ƺ=�� ��;��X�伀�;x��<X�=���<( <�������}4��ȑ�s-־�����>���k�Ә������R����������s쵿`2���4��@9��v�i�p�<�Х�j�Ծ�   �   1
���m����8Lt�(� �p}�<,�=�
=<��<@^��r������潃��l*K�yvq�d����㐾����~G��3���sh�$�?������ɽL�d�\P����R<�a=�<=$H8=��<����%\�2S��j��V���)���4�2�h��������e⾿WIп�=ۿ�޿��ڿ�3Ͽџ���[���"��4�g�v'4�"��   �   ��߾%���?�-��*���u�� ��<h�=�%9=Be)=|?�< ��;�-����@�8M����ٽ�+�Dn���'���*���$��.�+!��;�½q낽������<rf6=��i= Tu=T^P=Pd�<��X�������&�ߏ�_�ݾ�8�U��O��Ŧ�4�ÿ�rݿ���9���3������ouܿÿ G���(��XJU�����   �   �����P�c�׽���Ѕ-<|H=t�X=n�c=��K=��=�l�< ��9��$M$��Vk�q̐��頽Q��:y�����D�E�d���Jǻކ<��=Z�b=�3�=�i�=���=f�^=� �<�9¼����|�F��Z�������Q4�Qq�ǵ��Fn���ۿ�B���l�T��T��v���B���dۿ<z����3�r�y�5��   �   ��,,��8)k�!��jO=����;�=$*l=�h�=j��=�aj=�<=0=�:�<�0�;�w����������ؔ��`�(����:T1�<V!=�J=>V�='#�=��=�.�=��=xf=X��<�������_�ṾC<��E�����;���|˿2K�٪�5�m�-�������������̿� ��ań�K�G��   �   �z�S�˾�|��	�:?Y���(;�=Ƽv=y�=��=�Ҍ=��y=r�P=�g$=�v�<�<��f<Л+< 4)<@�a<@8�< ��<��-=<sc=�=Â�=㘶=�4�=�Y�=�`�=�Vi=\��<Z#�Q���3�o� �žN��/�P�`����ϯ�l�տ'���n�����/#��+&��)#�q��������L�ֿ���
��c�S��   �   R~�}%о6S����c��g�:TX=�z=L�=E�=���=W�=Nki=��A=֦=ؠ�<�h�<�̫<`�<��<P��<T#=n?P=�ˀ=�M�=d�=��=H{�=ئ�=~ť=�@j=�<D`$�����uu���ɾ�^�-nT�|��뿲�v-ٿ�:������2�� &��)�t&��I�D�+���aڿ�.��񤎿�W��   �   9z�6�˾Z�|��	�<<Y�� );��=ܽv=ky�=e��=�Ҍ=X�y=ڸP=,h$=Tw�<x�<��f<X�+<@4)<x�a<X8�<8��<��-=Nsc=�=Ԃ�=���=5�=;Z�=a�=�Wi=<� �E�����o��ž���8�P�ò���ί���տ&��0n���/#��*&�)#�Ŝ�k������`�ֿ+��g��a�S��   �   ���*��<&k�����I=�0�;��=@,l=_i�=
��=�bj=Ġ<=�=�;�<�4�;pt��T���D���������(����:p1�<x!=�J=`V�=[#�=6�=z/�=��=�	f=` �<v����A�_��޹��:�/�E�쯃�;:���z˿:I��������i��������{��̿/��*Ą�`�G��   �   ������P���׽���`�-<|L=d�X=��c=��K=�=8o�< �9�tL$�(Vk�?̐�頽�P��&y������E� �缰Iǻ�ކ<�=��b=/4�=?j�=���=��^=�*�<�*¼1�����F��W�����O4��Mq�ǳ���k��E�ۿ�?���j����{�"u�	����Aaۿ�w�����ӊr���5��   �   5�߾����V�-�$���b�����<F�=&)9=�g)=�C�<`��;+����@��L����ٽ�+�(n���'���*���$��.�!��,�½Y낽η����<~g6=0�i=�Vu=FbP=,p�<�X�=���:�&��ۏ���ݾ�5���T�.M���¦���ÿ$oݿ�{�5���1�������qܿ�ÿD��=&��PFU�����   �   ����m����B=t� � �@��<r�=�
=��< �����]���3�@��5*K�Pvq�V����㐾����zG��1���sh��?������ɽ��d��N���R<fc=��<=~L8=��<``��\�N���j��Q��v&�S�4��h��
�����X޾��Dп>9ۿ`�޿�ڿl/Ͽ����@X�����ԋg�#4����   �   }	��ڙ4�U���=� �E;h8�<н�<ԧ�< @��j&"�Qn��R����J����ʣ�`��.ZԾ?�����߾�Ѿ�s���;���}���=��� �p;������;<��<Љ=P��<�G<��+𽽞v4�{Ñ��&־M����>��k����u����M������{���絿�-���0���5����i���<�k����Ծ�   �   3�T�(�����l�p�Q�h�e<d��<���<`�2��k�p��V���;e��v��~Ⱦ4H�C���y�K�#�x&�U�"����op	��쾰¾L����Y�V�l����7�����;�<x�<$�<�J�j7q�G ���X�ӄ����㾨��CW:���]�m�|�k����2��$���$���刉�<>z�	�Z�ߡ7��-��!�j����   �   ��ؕ���ɼ���;T��<,�<� �;p��񶠽\��o]j��Z����޾�V�A(���@��%T�i1`���c��"_�0R�;W>�d%�rx	�S�پ�����-b���ߕ��ɼ�f�;؋�<d�<�<�;��鼢������&Xj�~W����޾�S��=(��@��!T�N-`���c��_�,R��S>��`%��u	���پɓ���'b��   �   Ⱡ�H"�����;p�<D�<t�<�J�?q�@
 ���X��������;Z:�r�]�T�|�����5��m���j������HBz���Z��7�d0�7&�����0�T�X���^�l��Q�@�e<��<���<`R2��b��x��ڼ��5e��r���Ⱦ�B�4���v�ß#�st&�į"� ��Lm	�z���¾H�����Y�Q��   �   |�� վ;���<��=���<@<��O����y4��ő��)־T���>�2�k�斋�{����O��b���L~��굿+0���2��p7��T�i���<����'�Ծ*����4�YZ��RD��cE;�6�<,��<\��< ���"��f�������J�N��Jƣ�f���TԾ{��.��<�߾�Ѿ�n��=7��:�}�4�=��� �<3���   �   �R<dj=@�<=�N8=��<����\�'P���j��S���'�Q�4�a�h���؆��N྿Gп�;ۿ��޿8�ڿ�1Ͽ֝��#Z��\!����g�e%4��������m�D��TDt�@� �X��<J =�
=8ï<�
��(��د�����{��n#K��nq����Eߐ�����B���{��1kh��?������ɽl�d�45���   �   �n6=~�i=�Yu=�cP=�o�<�X������&�ݏ�Ǎݾ�6�\ U�LN���æ�y�ÿ�pݿ�}�7���2�Ψ�� ��sܿ�	ÿ�E���'��wHU�P����߾������-�n'���j����<n�=B+9=l)=P�<0 <|��l�@�0D����ٽ�%��g�5�'���*���$�3(�|��ţ½S₽���@<��+�<�   �   �6�=#l�=,Î=��^=�)�<�.¼����F�Y������<P4�?Oq����� m����ۿ)A���k�i��g�v��������bۿy������r�I�5������>P���׽���(�-<BL=��X=h�c=��K=�=�< �9(٥��>$�~Fk��Ð�|࠽�G��p������E�q缐�ƻ��<��=��b=�   �   ��=�0�=p�=�
f=  �<���I��@�_��߹�i;��E�i����:���{˿J�@������}��������������̿ ���Ą�~�G�l��P+���'k�M���L=��	�;��=�,l=-j�=^��=�fj=��<==�J�<�y�;@&��ڈ����T����}��`�(����:�C�<�)=�J=6Y�=�%�=�   �   �5�=�Z�=�a�=ZXi=X<� ������o�X�žȄ���P�����ϯ��տ�&��qn�9��h/#�;+&�x)#�"��������ֿ�������S��z���˾q�|��	�">Y�@�(;(�=��v=�y�=���=�ӌ=��y=��P=�k$=L�<��<P�f<H�+<�I)<�a<�B�<��<�-=*wc=���=8��=��=�   �   n��=���=��=�a�=��*=`3ϻZ_����+��7��3�R=$���\��G���ˬ�1�ʿ���k���M����N����3�|�˿䥭��Z���p_�,'�}y쾙���t�<�����`�=x<�5=��{=�m�=*�=.Џ=Y�=�r=��W=v?=��*=L�=�y=<=�L/=�0I=�|k=	�=���=r�=��=}.�=�   �   m�=<J�=��=&ޖ=V0-= ;���Ȓ�sW'�������R0!��Y��݊�	쩿C�ǿ~�>���%�vm�
�$����:�H&ȿ�����Ջ��T[���#�y��>���8��5���༄��<Td6=
z=1�=��=��=�s|=�+_=�y@=��#=.T=d'�<�5�<�S�<P=Lq'=�L=f|w=#�=�8�=�¾=�%�=�   �   �9�=�=�b�=��=~�3= n��#�����2����XԾAQ�֛M��Ӄ�E���m����!׿���U���c����x���꿪׿�+������~����eO������پ�莾��)���������ޟ<��9=&t=�9�=U4�=r�o=��L=�u#=<G�<��<�:<pZ�;`�7; f;�v <��<|��<ě =~Z=��=��=¸=�   �   �|�=F��=�ϫ=^H�=|~<=@H�;�?S�d��ft�u����m
�~�;�̂q��Z��eƮ�#ƿ�Oؿ���A����G�׿�ſY����b��r�{�<�`��'�þ,~����%%��P�H��I�<�==0h=��n=��Y=��0=�!�<�fo< X��4k��x����*�/� F0��(�T[輀�l� i#;d�<޿#=
�k=�(�=�   �   �0�='
�= G�=c�=��D=��j<.����۽[ O�ə������$�{$U�4j���8��+������@�ʿOοہʿ1忿w���s����T��%���z���'V��X�`�G��[��p��<�^==�S=�ED=.Z=�J�< pZ������O=��O�������ҽ}��9�潌�ڽV%������b�S���ռ L�8�^�<�>=�   �   �=�^=ٻ�=�f~=,8I=���<�8���5���w%�2���ɾ��
���4�0`�7ք�< ���c���a��[N��Pϛ��2��*��^���3�>Z
��qɾ����(6)�߬���S�h32<LZ=�x7=�73=�=P�l<H�0��'�����!޽����H.�}E��R�v;V���N���<�03"�l7�tJ���@]�8���=<�   �   �L8;�^�<��B=B@]=�G=�,�< nI���V��u���S�Dd��cྙ�4u7��Z��fy�����V��FŒ��ۏ�懿@w�e=X��[5�$Q��;ݾ�w��i�Q�����@`������<Z�=�>(=*g=0 X<��x��2S�_<�������B���r��Ȏ�![��ꙩ�){����������+<��<�d�Ċ2����[ԛ�����   �   �� ��8t0�<F�/=j�;=�=`4F<�ּ�g���-��q��ƫ�Pl便��:,��BE���X�|Ee��/i��Qd��'W���B�_�)�����߾�g��(�i�cZ��v��4�Ǽ��;<�t=�#=�V= 9�<(@J��W��cҽ�L%�[�g�H7������Gվ�0���������N�����X�Ͼ�9��2��x�X�o��~���   �   ����J���];���<D�%=� =�D�< B2��?2��ǽ�J(�jx�t"����վF5�s��rI$�~�-�\�0�-���"��r�
�����Ͼ�� #l�w0�T��A� �];@��<��%=� =�=�<��2�NI2���ǽwO(�`x�3&���־�7�l���L$���-���0�e-��"��u�%����Ͼ]��(l��4��   �   ^��{����Ǽ0�;<�r=�#=<Y=�B�<� J�$W��[ҽ�G%��g�r3�����9վ]+�;��������������i�Ͼ45��x��RX�� ��v��j�� �8\;�<J�/=*�;=��=�#F<ּUm���1�q�&ʫ��p�J��0,�EFE�\�X�5Ie�T3i�6Ud�z+W���B�5�)�D
���߾k���i��   �   F�Q�&����G`�x����<�=(@(=�j=p9X< �x�&S�14��h����B�Z�r��Ď��V��:���lv������^��'8���d���2��	��7̛�އ� �8;�l�<h�B=�B]=�G=�(�< �I���V�b{����S�g�������w7�҂Z�*jy����W��<ǒ��ݏ��燿iCw�^@X�B^5�>S��>ݾ�z���   �   �����8)������]�@(2<ZY=ny7=�:3=а=(�l< v0�\�'�엽޽
��kB.��	E���R�4V�ƪN��<��,"��1��@���0]�d��@6=<�=l�^=���=h~=�7I=���<�B���9���z%�#4���ɾ��
���4��`��ׄ��!���e���c��GP��3𭿖����3�������^���3��[
�btɾ�   �   7��'*V�9\���G����� ��<F_==ȂS=ID=�_=�Y�< �3��ܺ��A=�+G��'쳽��ѽ��P��ہڽ'��b�����S��ռ ��8�r�<�>=�3�=/�=8H�=zc�=�D=��j<��d�۽3O�Ǜ�����J�$��&U�qk��7:���,��R����ʿ�Pο��ʿ�濿�x��C����	����T�~%�x���   �   ��þ.~�j��'����H��G�<�==fh=��n=��Y=��0=X/�<��o< ���S����r��|/��60����>輸�l� &$;�,�<��#="�k=o+�=�~�=���=�Ы=�H�=�}<=�4�;�CS����t�,���o
���;���q��[���Ǯ�uƿPQؿ]�㿼���㿥�׿D�ſo����c��r���<�V���   �   ��پD鎾��)�����	��<ݟ<��9=�t=d:�=�5�=�o=Z�L=z{#=`T�<��<��:<�; 88;�g;� <@�<`��<f� =Z=ؾ�=&�=�ø=;�=��=fc�=��=��3= u��ߟ��Ҩ�'����YԾ R��M�Tԃ����N ���"׿���j���w����y���꿉׿�,��D�������fO�����   �   ߡ羆��"8�T6��8��<dd6=�
z=��=��=��=0v|=�._=}@=��#=xX=�0�<T?�<x]�<#=�u'=�L=(�w=�$�=	:�=�þ=z&�=�m�=�J�=��=ޖ=�/-=0F���ɒ�KX'�����a���0!�kY� ފ�|쩿ìǿ�����o��m�Q�����O;⿨&ȿ����Ջ�PU[�<�#��   �   Hy�o���5�<�{���t��>x<�5=�{=�m�=L�=UЏ=��=n�r=�W=�?=�*=��=&z=N<=�L/=�0I=}k=�=���=z�=��=q.�=j��=���=��=�a�=`�*=�7ϻ�_���+��7��q�v=$��\�H���ˬ�E�ʿ��y���M����N����&�h�˿ϥ���Z���p_�'��   �   ��羠���8�~4����߼ȅ�<�e6=�z=��=��=��=�v|=F/_=�}@=*�#=�X= 1�<�?�<�]�<$#=�u'=�L=F�w=�$�=:�=�þ=�&�=�m�=�J�=F�=�ޖ=*1-=�3��PȒ�W'�����4��0!�kY��݊��멿�ǿ�������0m�������V:��%ȿB���FՋ�GT[�k�#��   �   F�پ�玾-�)�Y�������<��9=t=K;�=L6�=:�o=��L=x|#=4V�<d�<H�:<��;@>8;�g;�� <��<���<�� =JZ=���=@�=ĸ=[;�=b�=d�=��=��3= B��������������WԾ�P��M�(Ӄ���������!׿���U���U����w���꿱׿+������ρ���dO����   �   Y�þS)~���,"��x�H�R�<�==zh=��n=��Y=��0=�2�<8�o< ꃺxQ��T��Ľ��{/�v60�b�X>���l� )$;P-�<��#=��k=�+�=I�=X��=�ѫ=�I�=��<=�e�;;S����Yt�����l
�K�;�M�q��Y��ZŮ��ƿ�Nؿ{�����
����׿��ſ%����a���r���<�3���   �   `
���$V�#T�J�G� ������<d==x�S="LD=b=�]�< P,�Lٺ�@=��F���볽Y�ѽt��潷�ڽ��G�����S�8ռ 4�8\s�<X>= 4�=��=UI�=&e�=رD=x�j<l����۽��N��������$��"U�i���7���)�������ʿZMο�ʿ�㿿~u������1����T�;%�b���   �   �����2)�ާ��4D�(M2<2`=�~7=�>3="�=�l<xl0�F�'�6뗽C޽���'B.�f	E���R�4V���N��<��,"��1��@���0]�����8=<�=�^=ž�=�k~=D=I=��<t+���1���t%�0����ɾ�
���4��`��Ԅ����b���_��sL��l쭿����Y0���탿˜^�R�3�cX
��nɾ�   �   ��Q��~���5`�������<خ=nE(= o=�FX<�x��#S�)3�����"�B��r��Ď��V��+���av��򠧾X��!8���d���2��	��̛�@����8;�o�<؋B=NF]=�G=$9�< �H���V��o���S��a���߾���r7��|Z�acy����� T��TÒ��ُ�5䇿�<w�J:X��X5��N��7ݾu���   �   1V�.p��PqǼh<<�{=��#=T^=�J�<�J��W��ZҽNG%���g�D3��舷�վH+�.��������������e�Ͼ.5��r��?X�h ��v��n�� �8$@�<��/=��;=��=�QF<��ռb���)��q��ë�Fh�Q��f,��?E�O�X��Ae��+i��Md�r$W�~�B�k~)�I�G�߾dd����i��   �   ���@5��~^;Ԩ�<��%=>� =�M�<�2��<2���ǽdJ(��x�D"����վ75�h��iI$�x�-�Z�0�-���"��r�	�����Ͼ���"l�X0�����?� ^;���<��%=x� =S�< �1��42���ǽEF(��x������վ�2����IF$�)�-���0���,��}"��o�¥��-�Ͼ�顾�l��+��   �   .�� ��8XL�<��/=��;=��=�DF<|�ռ�f��B-��q��ƫ�'l侭��/,��BE���X�xEe��/i��Qd��'W���B�_�)�����߾�g���i�4Z�	v����Ǽ�<<,y=j�#=`=PS�<@�I�ZW��Sҽ�B%���g��/������Aվ�%쾆���/���ޯ��=~�_�Ͼ�0������xX�7��{n���   �   @�9;�~�<ʐB=
I]=@G=h6�<@6I�4�V��t��y�S�d��=ྌ�*u7��Z��fy�����V��FŒ��ۏ�懿@w�h=X��[5�"Q��;ݾ�w��I�Q�'����>`�h��D��<ڭ=xF(=<r=�\X<�|x�@S��+��0��J�B�"�r�����BR�������q��Q����z��4����d�`~2�6����Û��y��   �   � =��^=���=�m~=t=I=��<3���4��?w%��1����ɾ��
���4�)`�5ք�; ���c���a��\N��Rћ��2��,��^���3�<Z
��qɾ�����5)�N��� P�8?2<�^=�~7=�@3=N�=��l<�H0���'��㗽5޽a��<.��E���R��,V���N�<�<��&"�0,�7��6 ]��蝼c=<�   �   37�=(�=�J�=�e�=ȱD=��j<�����۽ O���������$�v$U�1j���8��+������B�ʿOο݁ʿ5忿w���s����T��%���q���'V�XX��G� ��(��<�c==އS=OD=�f=0k�< (	�,ú��2=��>���⳽��ѽu�q��%wڽ����x����S�bռ ��8���<l>=�   �   z��=쐲=�ҫ=lJ�=��<=�Y�;�=S���+t�]����m
�v�;�ǂq��Z��dƮ�%ƿ�Oؿ���C�翀��J�׿�ſY����b��r�z�<�_�� �þ�+~�٣��$����H��N�<^==6h=v�n=��Y=F�0=�>�<�o<�����;��t��2��2m/��'0��
�@"��zl���$;�A�<��#=��k=�.�=�   �   �<�=i�=�d�=��=z�3= �������N������XԾ<Q�ӛM��Ӄ�D���l����!׿���Y���f����x���꿪׿ ,������}����eO������پ�莾��)�E��������<L�9=rt=�;�=G7�=
�o=R�L=D�#=�a�<��<H�:<��;`�8;��g;�� <�<��<�� =�Z=���=��=�Ÿ=�   �   �n�=hK�=��=�ޖ=N1-=�5���Ȓ�^W'�������O0!��Y��݊�	쩿C�ǿ~�>���%�wm��&����:�J&ȿ�����Ջ��T[���#�w��<���8��5��� ���<re6=�z=H��=d�=��=|x|=h1_="�@=B�#=R\=�8�<H�<Xf�<v'=z'=�L=ȃw=D&�=k;�=�ľ=w'�=�   �   �]�=,��=u>�=�ٶ=�(�=t�<$��+[ӽ��L�9	��v��%%�^�U��샿����F��D¿��̿�nп�̿�¿0}��2g�������W�Kl'�^t�������_�dI�*�s�@;���<V�+=��\=Zt=��y=6�t=��i=�]=,WQ=LH=|C=�)D=�@K=DY=�Vn=�=�ĕ=�`�=̫�=6+�=*+�=���=�   �   P��=�i�=�Z�=�?�=��=�"�<�a㼁�̽K�G��������h"���Q�U���W���L���Ⱦ��Rɿ{�̿`Mɿ�̾�Zq�������.����S��2$� m�٨�PmZ����2�h��!����<�V.=�\=��q=8�t=�l=��^=��N=�?=(�3=�,=�r*=
�/=2H==V�R=�Oo=8�=
��=�=�}�=���=��=�   �   �b�=9��=���=�8�=S�=0�<t��A����f9�Jz��N#߾*��F�c�u�ʜ��E����Y���`��$�¿�H��*;����������f�v� �G��������ܝ�(WJ�x��X�G�@J��̻�<Z5=�\=D�i=H�d=�QT=��<=l2#=�
=���<��<x�<X��<���<���<�7=&�E=L?t=[Ӓ=�=*��=�8�=�   �   �N�=�N�=�L�=�%�=$H�=�=pS����H#��ć���ɾ :�xe5��`�6x���������ɯ�b岿���B@��ֹ���M��@a�z�5��@�;����B1�&}��p1��5�;@��<<
>=��Y=T�Z=��H=�A)=��=D��< 2<@��:��ɻ�%7��T�0m6�5����o;�-�<d]�<�<=R�{=k{�=�"�=�   �   ��=�5�=N�= '�=��=��=�V�F�m��e�s�g�����O��4�y9F���k�$���i����ۛ�`���s���+#���
��G�j���E�U�����zY��+n��t�,ȓ��r���Lp<"D=�YF=�R=� B=�=ԇ�<��%< Cӻ8����ȀS�4	z����@����q��MC��U���O��/<pI�<�hJ=���=�   �   �n=`��=�{�=I�=ϵ�=�6=�)<J
�ȍн.t;�]��|F˾�$���'�"�H�j^e���{�^%���|��Є���z���c���F��&��
�@�ɾ)����d=�)/۽��@���\��V�<��/=f�J=:5B=�#=T3�<`�T;8⡼8�6�(��Z��\���(��,��p��ƽ�ؑ���.�п_��ed<vW=�   �   ���<�_T=�s�=A��=�I�=6�H=�u�<@���*�������Rb��5���YؾkQ�O�#��;�ʩN��Z�\v^���Y�+?M�g�9��u!�*,��PԾ������\�	�
�W��������m<��=��D=�IH=,B'=4�< ;�l׼�dr��W½K��5}*���I�Eb�|p�d�s��=k�C�W�Z�:�L���@޽�Y��8c ��L;�   �   ��L�0d�<,�D=�s=؋y=\U=`�=@��:��(��Ľ>i&�0[u�I-��<eӾ�8�����I"��+���.��+�D� �9��#���qx;���2�i�8���ֲ���0��;� =�0@=PS=�j<=�Q�<�]�;d�ɼF���1O߽�3"�v]V��S������˫�np���Z���,���W��\���/x�C�N��]5���J*��   �   ��.� ��k�<l?=@]a=�X=��%=�.�<�3t�l�k�+>཮�-�\	q�ʀ���^���d۾>��� ����Ĕ���ﾏ�վٛ���̓���`����?����.���� w�<�!?=�^a=ԶX=��%=&�<Ot�d�k�E�(�-�
q�@����b���i۾:��� �P��������վҟ��3Г���`�����F���   �   jܲ�����s�;�� =H.@=�S=�k<=dX�<@��;��ɼ�����G߽./"��WV� P��%����ǫ��k��6V���(���S���
���(x�NC�w���-���>*��@L��q�<��D=Ʃs=�y=�U=�~= �:�)���Ľ m&�L`u��0��%iӾh=��b��L"� �+���.��+�� ��������:|;#��3�i����   �   �
�ߨ��������l<�}=��D="JH=�D'=��<@y;PZ׼�Xr��O½����w*��I�p�a��tp��s�g6k�t�W��:�����6޽�Q��BV ���;���<JeT=�u�=[��=�I�=��H=Do�<����z�������Vb��8��P]ؾ�S���#�̽;���N���Z�yy^���Y�BM�	�9�Ax!�).�0TԾP�����\��   �   �g=��3۽�@�@8]��P�<@�/=p�J=�6B=�&=L=�< �T;Xϡ�8�6�� �����lR꽯���D'�m����;�ƽ0Б���.���_���d<�_=L�n=���=T}�=�I�=е�=�6=��(<6�<�нUw;�@_��FI˾F&���'���H�"ae���{��&��~���ф���z�:�c�G�F�ނ&�X���ɾ- ���   �   �-n��v�˓�{���Ap<�B=�YF=pR=#B=��=l��<��%<�һ@�����:rS�T�y���������F�q��=C��F�пO�^< ]�<�pJ==u�=�7�=n�=~'�=���=��=����m��g�v�g������6�n;F���k�e�����ݛ�Ț��җ��x$�����c�j�r�E�������R[���   �   �����C1�����4�p#�;x��<�	>=,�Y=��Z=�H=<E)=��=	�<H:2<���:@sɻ��6�`PT� =6�Pִ� �p;�B�<\p�<�<=l�{=Q~�=�$�=]P�=P�=tM�=&�=�G�=`�=XS����J#��Ň�G�ɾ!;��f5���`�+y�� ������˯��沿2���WA��Ӻ���N���a���5��A��;�   �   �ݝ�IXJ��彦�G��W�����<�5=B�\=�i=��d=$TT=
==�6#=�
=X��<@(�<"�<�Ÿ<D
�<Н�<�>=��E=|Et=	֒=l�=��=x:�="d�=��=6��=�8�=	�=@�<8y��B���eh9�M{���$߾�*��F���u��������Z���a����¿�I���;��S���2���o�v���G��������   �   ]٨��mZ�����6�h��$�p��<�V.=(�\=��q= �t=X�l=x�^=�N=��?=F�3=:,=>v*=� 0=,L==0�R=.So=�9�=���=L��=�~�=���=���=���=�i�=�Z�=�?�=x�=� �<e���̽2�G�E���_���"�\�Q������W��;M���Ⱦ�mSɿ��̿�MɿI;��q��J����.���S�C3$�wm��   �   p�����_�<I���s�?;�H��<j�+=��\=rt=Ըy=��t=��i=]=�WQ=rLH=�|C=0*D=AK=dDY=�Vn=��=�ĕ=�`�=۫�=F+�=4+�=���=�]�=,��=l>�=�ٶ=�(�=��<p��[ӽ��L�k	������%%���U��샿$����F��P¿��̿�nп�̿�¿&}��%g�������W�.l'�.t���   �   eب�\lZ�����"�h�h�D��<&X.=t�\= �q=�t=V�l=T�^=��N=`�?=ܨ3=�,=�v*=B0=fL==b�R=\So=�9�=���=\��=�~�=���=���=��=0j�=E[�=@�=�=�$�<�_���̽ޛG�Z���&��#"�c�Q�����V��{L��)Ⱦ��Rɿ�̿�Lɿt̾��p������).���S�q2$�1l��   �   �۝��UJ��彴�G� 3�����<�5=��\=Z�i=�e=�UT=�==8#=<!
=���<,*�<�#�<�Ƹ<@�<���<>?=6�E=�Et=-֒=��=8��=�:�=dd�=c��=Ċ�=�9�=A�=P�<o�������e9��y��Q"߾x)�6�F�h�u�5��������X��`��R�¿�G��[:��ܕ��ẑ�&�v��G����p���   �   L����?1��y���,�@V�;|��<�>=��Y=��Z=ԸH=�G)=:�=@�<PA2<��:�hɻ��6��LT��:6�pҴ�`�p;�C�<�p�<&<=��{=�~�=%�=�P�=�P�=@N�=K'�=�I�=N�= �R���%G#�}Ç��ɾ9�Ld5���`�`w���������ȯ�;䲿瘯�$?��ʸ��M���a��5�c?�/;�   �   �'n�r�pē�g��`p<�H=x^F=�"R=�&B=�=x��<��%< �һ�������pS� �y�6���`�����q��=C��F���O��_<�]�<fqJ=;��=��=#8�=[�=�(�=���=��= ���}m��c���g�,�����}3��7F��k�����#���Sڛ���������!���	���j���E����߁�XW���   �   Ta=��)۽��@� �\��a�<��/=��J=L;B=+=�D�< .U;\ɡ���6��������Q�^�P�'�J�����ƽБ�.�.�0�_���d<f`=6�n=^��=X~�=dK�=��=�6=)<��нq;�[���C˾�"���'��}H��[e�-�{��#��
{���΄���z���c���F��~&���Z�ɾ�����   �   ��
�򞐽Ж���&m<��=X�D=�OH=@I'=#�< �;�S׼�Ur��N½��0w*��I��a��tp��s�F6k�^�W��:�����6޽`Q���U �@�;`��<�fT=�v�=�=L�=��H=|��<����/S��kNb�F3���VؾoO���#�u�;��N��Z�Gs^���Y�;<M���9�ys!�*�VMԾϱ��4�\��   �   �ϲ�����;�� =�6@=h	S=Vq<=�a�<@��;��ɼ����9F߽�."�WV��O�������ǫ��k��#V���(���S��
���(x�<C�a��W-��>*� 2L��t�<��D=جs=n�y=(U=��=���:��(���Ľ2e&�Vu�*��laӾf4��O�G"�1�+���.���*�|� ��������vt;���ȟi����   �   ��.�������<�(?=ea=�X=��%=�6�<@%t�@�k��<�
�-��q������^���d۾ ��� ���������ﾉ�վԛ���̓��`���{?���.�@���z�<�$?=ca=ּX=@�%=�=�<�t���k��6��-��q�V}���Z��t`۾P��t� �����������վ����@ɓ�{`�1��8���   �   ��K�0��<�D=�s=��y=�U==@
�:z�(���Ľ�h&��Zu�-��
eӾ�8�����I"��+���.��+�B� �7�����kx;��� �i���1ֲ������;~� =(4@=�S=>r<=�f�<`��;0�ɼ׳��Z?߽(*"��QV��L��E���~ë��g���Q��$��yO������!x�BC�`��4%��:1*��   �   ���<�lT=�x�=+��=�L�=��H=\}�<��������Rb��5���YؾXQ�A�#�	�;�ũN��Z�[v^���Y�+?M�f�9��u!�(,��PԾ������\���
�죐�����m<��=�D=�OH=&K'=p*�<�;C׼nJr�vG½����q*�"�I���a��mp���s�+/k���W���:���-޽.I��\H ���;�   �   ʪn=Ǽ�=��=ML�=H��=~6=()<����н�s;��\��TF˾w$���'��H�f^e���{�^%���|��Є���z���c���F��&��
�:�ɾ!����d=��.۽��@�@�\�t[�<R�/=��J=r<B=�-=@M�< �U;@�����6�������fH�J����!������H�ƽAǑ���.�xW_� �d<�h=�   �   a�= :�=��=�)�=��=��=�
�X�m�Je� �g�ٳ��4��4�q9F���k�#���i����ۛ�b���u���,#���
��H�j���E�S�����tY���*n�st��Ǔ�Xp�� Tp<�F=�]F=8#R=z(B=2�=���< &<��һ�＼��&cS�$�y�>���)x��Z�q��-C�8���O���<Xq�<�yJ=w��=�   �   �R�=�Q�=O�=�'�=�I�=R�=�S�����H#�{ć�l�ɾ�9�se5��`�6x���������ɯ�d岿���D@��ع���M��?a�z�5��@�;����B1��|���0��@�;D��<>=��Y=��Z=غH=�J)=��=l�<@]2<���:�ɻ(�6�� T��6�Pw�� kq;X�<���<H<=��{=k��=n'�=�   �   �e�=@��=O��=�9�=A�=�<�q��ͱ���f9�7z��?#߾*� �F�a�u�ʜ��G����Y���`��&�¿�H��-;����������f�v�!�G��������ܝ�WJ�L����G�`C��P��<.5=��\=��i=e=�WT=T==�;#=�%
=���<�5�<\0�<�Ը<d�<Ĭ�<F=��E=�Kt=�ؒ=�!�=��=$<�=�   �   ���=�j�=�[�=9@�=(�=L$�<�`�R�̽2�G��������g"���Q�U���W���L���Ⱦ��Rɿ{�̿`Mɿ�̾�[q�� ����.����S��2$� m�٨�GmZ�՞����h� ����<�W.=X�\=>�q=��t=�l=n�^=N�N=:�?=�3=L,=�y*=\0=�O==��R=�Vo=^;�=	��=���=��=���=���=�   �   R�=~X�=�,�=�'�=0�=,Q=PM<�D�w���FC[�32��������!@�#e�������0:��A���:��J���&����e��7A� ���2�١��cp�$��m_�����@�����<���<�9=�a=r=D�=jF=��=�)!=�+=�+:=^�L=v	c=�}=>M�=���=�`�=��=�l�=���=���=�h�=�   �   ؞�=W��=�r�=Lj�=rx�= �S=��$<�,;����0V������{�F����<�qa� ���Uo��
���M`��А���q���ˀ��a���=����N꾢Ϊ��Ij��Y��ɥ�D�� X7��)�<�U�<��=V=��=�7=l&=�=6�=�H=�^)=��9=��N=��g=䴂=�i�=5��=���=t�=J��=��=a��=�   �   �g�=�l�=6"�=f��=D�=d�[=(�e<�D ��eݽ��G�O����2ؾA��s2�e)U�6�s��"��F㍿-���ҍ�D��a�s��XU�R	3�G��zܾ���M[Y�*��勒���ἠ�);�n�<xi=�=�w=�=�	=���<���<D*�<�2�<Xp�<l =d�=jV'=��D=~�g=S�=�m�=;�=<��=�4�=�O�=�   �   TV�=B\�=O��=�N�=<A�=Ig=�<<��ཽ�0�c�����þ����"���B��_��du�Ձ��<�������t��^�6CB���"�'��ƾ|l���>�X_�_i����83<���<�=>{ = ~="�	=��<8�<�)�<0�H< �<� �; ��;0N< ]<p��<���<��)=Rr]=�ʉ=�8�=p5�=���=�   �   b��=���=?��=��=�#�=�s=�-�<�ȇ�A���BX���l�\���/	�i�M�*�lGD��:X�G�d��"i�	~d�XzW��\C��*����rS����
q�>f����� ��0!��<n=*�(=Vv(=^�=T��<�q�<Hq< M����4�Ȕ��ּ�����U���?ݼ<����f�`��;�i�<ZF=~a=��=`ج=�   �   nA�=9T�=ߖ�=qI�=6��=��}=�=`�I���V�K�齸�@�����S�����kF��&��57�B��E�k}A��6�p�$����H��,���{����?�L｜hv�(Ҍ��ZZ<��=�0=,;=b�+=	=�b�<�S�;P�!��Rܼd�2��\q�����ٔ��%����7������p���7��ż@Aʺ��<�/=��|=�   �   ~2^=�^�=v��=ጧ=��=�ځ=z�)=�A%<,���u䩽���غ]�l������p�\��f�����>� ��k�h��o~�9w������S��L��矽N����;ܹ�<p6=n�N=�H=L�'=tX�<��<��C��Y�t�{�.7���b�D���]����F�7"����I�߽����xgU�l���K�;l=�   �    "�<x�I=�ȃ=E�=�k�=Y�=D	?=L�<�?�p�[��Խ>@%�0�e�	��>T��H�о�F�M@��{f���A�e�{Y˾�^������fT�����,���q$��_����<®9=��a=��g=��N=�B=�>�<0�޻*a�1����ؽ���&�5�(�T�P�l�H�z��q}��Vt�E`��@B�������C����@*��   �   0g����<X�>=�
t=ө�=^�y=N�K=���<�â;�N弴ǉ��7彂7$�f<W��+��Mԙ������������l��⦥�[�����u��NA�����	��2�-��!��T��<H�>=Ht=㪃=8�y=��K=p��<0��;�[�h̉�)>彔;$�lAW��.���י�f���w�������o������������u��SA�@�����V�-��   �   �z$� G���<Ԫ9= �a=t�g=��N=JD=E�<P�޻xY��+��žؽ���*�5�|�T��l���z��j}�Pt���_�";B�o��"�q<��������L1�<J�I=�ʃ=��=\l�=6Y�=�?=8�<��?�8�[���Խ�C%�ԝe�����W���о�J羰D���j��)F��i�B]˾?b��d���kT�����2���   �   �쟽 ]��ן;p��<f6=��N=j�H=��'=�\�<��<��C��Q���{�m0���Z㽲���X�)��WA��������߽v����XU����� ��;�
=9^=�`�=<��= ��=X�=gځ=��)=`3%<�����詽��ξ]����
����s�h�����5���� �^�Em�i�����?z������$�S��O��   �   ��ov�\݌� JZ<f�= �0=;=d�+=\	=8h�<0w�;H{!�dBܼ��2�BPq���������Ί��V/��W���`���7��{ż@�Ⱥ��<�#/=Z�|=D�=6V�=H��=JJ�=|��=��}=�=`(J���V������@����������?H��&��77�YB�n�E��A��!6�l�$����K�:/���}����?��   �   ph�p����� p!��<�k=��(=�u(=��=���<�w�<ȃ< �����4������ռL����<���%ݼ�����5��R�;0~�<hO=B!a=��=�ڬ=l��=f��=P��=���=�#�=�s=`)�<�Ї�H���lZ��l�M����⾐j��*�WID��<X�p�d��$i�(�d�Z|W��^C��*����UΆ���q��   �   ��>�b�Nci�����-3<���<�~=�z =R~=6�	=��<�%�<l2�<P I<��<�]�;���;(r<�,]<�è<t�<��)=�y]=�͉=�;�=�7�=���=�W�=Y]�=
��=NO�=0A�=Hg=��<T��⽽��0�����V�þ��ݏ"��B�!_�wfu��Ձ��=��粁�Q�t���^��DB�ד"��ƾ�m���   �   �\Y���j���P�ἠ�);�k�<ph=z�=�w=�=:�	=���<4��<�1�<�;�<`z�<� =B�=n\'=��D=J�g=�=Jp�=7=�="��=46�=Q�=�h�=�m�=�"�=���=+�=|�[=�e<�G ��gݽ�G�L���:4ؾ��t2�{*U�h�s�J#���㍿ׇ���ҍ����x�s��YU�!
3�����ܾQ����   �   �Jj�Z��ʥ�x��`h7�,(�<�T�<6�=J=��=:8=�'=��=6�=bK=:a)=��9=ڿN=��g=t��=ok�=���=�=+u�=@��=���=
��=\��=���=�r�=Vj�=Tx�=|�S=��$<j.;����1V�.����|����C�<�a�v����o��e����`��&���,r��?̀���a��=����N�Ϫ��   �   9p�	��M_��Է�������<t��<�9=�a=�=x�=�F=2�=T*!=l�+=^,:=�L= 
c=}=qM�=���=�`�=2��=�l�=��=���=�h�=#R�=�X�=�,�=�'�=�/�=�Q=`K<��D������C[�^2��������!@�+#e�������7:��D���:��F���&����e��7A���s2ﾾ����   �   Ij��X��ȥ�����D7� ,�<X�<ּ=�=V�=�9=�(=��=H�=>L=�a)=��9=\�N=T�g=���=�k�=���=��=Bu�=U��=���=��=|��=ޣ�=s�=�j�=�x�=��S=P�$<�+;����@0V�C���q{���^�<�a�ⱀ�o�������_��y����q���ˀ���a�-�=�J��YM�Ϊ��   �   �YY�������ęἀ*;Hs�<�k=��=rz=L=ܣ	=l��<���<�5�<�>�<L}�<0 =8�=6]'=*�D=��g=7�=sp�=^=�=C��=[6�=3Q�=&i�=�m�=#�=B��=&�=L�[= �e<B ��cݽb�G������1ؾ���Qr2�~(U�.�s�"���⍿����]э����4�s��WU�`3�y��(ܾx����   �   ��>�\�Zi����(F3<<��<f�=�~ =j�=
�	=T��<@,�<�8�<8I<(�<�m�;���;xw<1]<XŨ<��<��)=8z]=Ή=�;�=8�=���=(X�=�]�=���=>P�=�B�=�Kg=��<���Nݽ�P�0�>���1�þ%���"�X�B� _�cu�2ԁ��;�������t�v�^��AB�k�"����žk���   �   �c�1�������� ��%�<6r=��(=${(=��=��<���<�< ����4�t|����ռ�����9��d#ݼ̆���2�W�; �<�O=�!a=�=J۬=���=���=��=���=z%�=Θs=�6�<𽇼Ӌ��V��l������⾼g���*��ED��8X�1�d�t i��{d�LxW��ZC�A*�9���P������q��   �   ���&`v��Č�PqZ<��=�0=P;= ,=�	=\r�<`��;�i!�\:ܼj�2�6Mq�8������������.�����`�H�7��zż��Ⱥ� �<�$/= �|={D�=�V�= ��=�K�=L��=&�}=� =��I���V�E�齅�@�򂌾�	����ﾭD��&��37��B���E�{A�I6�^�$�E��uE�*���y��$�?��   �   {⟽�<���<�;���<�6=��N=ƝH=��'=�g�< �<0�C�M���{��.��UY���qX����A��������߽6���DXU�����p��;T=�9^=�a�= ��=J��=3�=݁=.�)=X]%<<���%ߩ�����]��������wl�]��6������ ��	��h�W���z�t��f�����S�I��   �   �f$�@Q��� �<ƴ9=<�a=v�g=��N=�I=�O�<��޻�T��)��ܼؽ���t�5��T���l�U�z��j}��Ot���_��:B�O���~�5<��\����� 3�<��I=�˃=��=0n�=�[�=R?=t#�<��?���[���Խ-<%�?�e����P��x�оjB��;��b��a=�a㾕U˾k[������aT����&���   �   �ә�$��<��>="t=���=�y=�K=L�<��;�E弝ŉ��5彦6$��;W�V+��ԙ�����i��������k��Ӧ��L���߻u��NA�����	����-�������<��>=�t=���=��y=t�K= �<0�;\:�}���D0��2$�
7W��(���Й����������h�����ሒ���u�pIA�l��y�� �-��   �   �B�<j�I=΃=t �=o�=\�=b?=��<��?���[�D�Խj?%�v�e�����S���оkF�2@��if���A�e�oY˾�^��|���fT����l,���p$��A����<ʰ9=��a=�g=��N="K=U�<`\޻N��$����ؽ���Ј5���T���l���z��c}�VIt���_�35B� ���u꽝4����@���   �   n@^=d�=꣢=v��=��=݁=ض)=�Q%<�����⩽,��/�]�"�������o�J��W�����7� �	�k�f��g~�2w������S�{L��矽�L����;4��<�6=�N= �H=H�'=Pk�<��<�kC��E���{��(���Q�÷��S�����;�T�����߽�zIU��}��p��;�=�   �   "G�=�X�=���=lL�=���=��}=V=`�I���V����"�@�������ǉ�YF��&��57�B��E�j}A��6�o�$����H쾸,���{����?���gv�lЌ� `Z<��=�0=@
;=,=�	=�v�<��;�S!��+ܼ*�2��Aq�������������&������<P���7�P`ż@CǺ�4�<�,/=��|=�   �   ���=|��=(��=`��=�%�=@�s=�3�<�Ç�(����W���l�-���	�i�A�*�eGD��:X�G�d��"i�
~d�YzW��\C��*����mS�����	q�)f�٫�� �� !� �<8p=H�(=�z(=J�=���<���< �< l����4�l����ռ���H"��$ݼ�n����`��;@��<�X=R)a=N�=�ݬ=�   �   �Y�=�^�=q��=�P�=�B�=fKg=�<���<߽���0�<�����þ����"���B�}_��du�Ձ��<�������t��^�5CB���"�%�ƾyl�� �>�-_罜^i����h<3<���<H�=d~ =l�=��	=P��<(1�<�?�<XI<@�< ��;��;`�<pR]<<֨<<"�<:�)=R�]=*щ=p>�=K:�=���=�   �   j�=�n�=�#�=���=4�=��[=@�e<�C �"eݽW�G�8����2ؾ8��s2�b)U�4�s��"��G㍿.���ҍ�E��c�s��XU�S	3�F��wܾ~���B[Y���å����ἠ�);�p�<�j=�=Vz=�=��	=$��<���<�:�<�E�<(��<� =�=Zb'=l�D=��g=��=�r�=\?�=���=�7�=]R�=�   �   ��=4��=Zs�=�j�=�x�=��S=H�$<,;�o��0V������{�D����<�qa�!���Vo��
���O`��Ґ���q���ˀ�!�a���=����N꾠Ϊ��Ij��Y��ɥ����R7��*�<8W�<��=�=`�=�9=F)=~�=:�=�M=�c)=\�9=n�N=��g=ķ�=�l�=ͥ�=	��=0v�=��=���=���=�   �   i>��>���=�K�=^Q�=�j�=D1%=�/��9l���U8U��N���Ѿ�����8�nHK�l�W���[�#�W��ZK��P8�Y_ ���P^վ}U��\�j�-
 �9�˽Sm��@����O���z� -*� L4� !���f+� ��@��:�g�;�7^<�4�<��=�-=�DX=���=�&�=1�=���=���=���=]��=D� >��>�   �   ��>g�>�L�=T�=O�=��=�V(=�.��j�b�4�� gP�a����̾���m����4�׍G���S���W���S��G�)�4��C���"�о1���b�d�h����Ľf�a����+.����Ā:�=:��F��2�@z��@��:P5�;h�G<��<X��<X� =&VJ=�t=���=暤=L�=,�=Dk�=��=
��=��>�   �   "3 >���=0,�=D5�='�=�V�=�1=�35;�eH�w罂�B��Ď�����:����8�*���<��:H��%L��H�-�<�v�*�J>������þ(5���2T�`�:ǯ��0@����������T;P��;��;@�; �S9 �B� �'9�H;�!�;@�e<��<Ф�<f�=x�F=�0p=�r�=D�=Z��=��=�0�=��=R�=�   �   ̍�="��=�%�=�h�=2��=cʘ=g==�6<h) ��Cɽ�--�wh��v���m޾���b��+�\6���9��6��h+����.�2g޾Ư�[փ��%:����:+���u�h"���;`n9<P�O<��-<���;�2=; \�� ���� ��`g9;��;@�[<�T�<���<=��J=z=B�=5%�=cu�=w��=�z�=�   �   ��=8��=��=�O�=H�=Q�=ֺJ=�A�<<�޼Z��ݶ�]�S��������I���w�ε�K�"�lD���u��r�辷ÿ��8���*^�@�B��JK�l򏼀ay;@��<���<䡭<P�<hJ?<�1�;@�����ԻX%.���Z��m��c�`69���׻ ��9�<�@�<�
=D=Ԩ~=|��=1�=P�=�   �   Hf�=ҟ�=�S�=S�=-��=ɗ=��U=��<�ao��x�y��ɟ5�*o{�p졾Až<X�T����?������O����ྗ���/L��l�r��Q/�i)������ؼ���:(~�<���<�=�L�<U�<�߀<P�; z���fp��Ƽ�{�FK!�4��y;��W5�2[ ��d��������;���i<|.=��L= �=	�=�   �   �Y�=�B�=2ö=0��=oM�=�%�=��[=���<@�8��*�8U������G�)����7��d���w�˾_�׾@�۾6�վ�Ǿ&��	<��1s�O'7����Ę��u
�@ � �<��=ȏ.=t21=�:=���<�&�<�~;��=��a㼞4� �s����ά���������h���Ĩ�iS���M�H�뼀���hR�<0"=�l=�   �   xYO=r��=���=(%�=\ �=j��=nBZ=*8=��;<ʼ��{��ҽ���X�E��|r�����9�����fŧ�3���W�������x ^���-� ���o������j�,x�<��%=�WR=Ԯb=��Y=��:=F	=�u�<@Lغخ��r%?��]����½M𽎠������ �;7 �S���.߽g�����V�8*���~�;x��<�   �   ���<t�8=��p=���=ӌ�=6�{=�_O=0�=�Fc<�$7���#�_���Kؽ&"�tN0�M���b�A�o�~iq��h�X6T�v|7�Fi���۽� �� sƺ<�<B�8=v�p=h��=H��=>�{=aO=�=`@c< 27�v�#�X���Pؽ�%��R0�:M�+�b�ڌo�4oq�6h��;T�k�7��m���۽a����� �Ǻ�   �   `hk��k�<��%=tSR=p�b=&�Y=��:=pE	=w�<@غ����:?�lY���½�x𽙜�K��G� �i2 �:N�����%߽ƨ��ByV�|���ʳ;�<�_O=��=��=�&�=��=#��=�BZ=H7= �;#ʼT|���ҽ���C�E���r�r���
<������ȧ�]���[�������h%^�3�-�C����t��6��   �   �}
�`{ �hޫ<8�=�.=t/1=�8=d��<�&�<�+~;��=��X� 4�X�s�����Ȭ�e���q���a������K��ԟM����P@���e�<:*=ԉl=�\�=�D�=�Ķ=z��=TN�=.&�=v�[=`��<`	9��*�Y��z�-�G�N���&:��M�����˾� ؾ��۾��վS�Ǿ���>���5s�
+7�(���ɘ��   �   �Ã��(ؼ �:Du�<���<�~=�G�<|Q�<$ހ<P�;�l��0Zp�<ƼRu��B!�N4��n;��K5��N �L�������;���i<�7=��L=e#�=��=�h�=���=BU�=T�=΂�=6ɗ=��U=��<Ppo�>x���뽌�5��r{���ž3[侏���kA�R��͏�CR�����-���hN���r��T/�F.��   �   �E��	K���� y; ��<���<���<L�<�E?<@/�;���� �Ի�.�P�Z�0zm�`cc��9�0O׻ B�9��<S�<ľ
=�D=�~=���=��=2R�≠�=���=���=�P�=��=Q�=ܹJ=�=�<��޼/��ܸ��]��T������J뾭��Oy�f���"��E�����������ſ�p:��K-^�y��   �   ���-��z��-"��˓;@c9<؈O<�x-<@��;@)=; <���q���� T�� �9;�2�;X�[<�a�<8��<�=V�J=lz=E�=�'�=�w�=^��=j|�=��=$��=�&�=>i�=d��=?ʘ=�e==@.<�, �Fɽ�/-��i���w���o޾���c�N�+�h]6�<�9�G6�9j+����/��h޾ǯ�~׃��':��   �   a��ȯ�t3@�������� �S;@��;0�;@�; \S9 �B� �(9��H;�3�;�e<��<��<ԅ=
�F=�5p=�t�=b!�=T��=���=w2�=K��=e�=�3 >P��=�,�=�5�=:�=�V�=1=�5;bhH�y��B��Ŏ�����b;�����*���<��;H�~&L�~H��<�E�*��>�9�����þ�5�� 4T��   �   ���Ľ��a��ἐ1.�������:��<:��F��<�v�� ��:�<�;�G<8�<x��<�� =�XJ=��t=�=��='M�=:�=6l�=���=���=*�>��>��>(M�=<T�=P�=���=V(=@T��(�b�X5���gP����^�̾�����4�]�G�-�S��W��S�}�G���4��C�����о�����d��   �    
 �7�˽:Sm�DA��@�O���z��A*� [4��#�� f+�@�뺀��:�l�;�:^<l6�<��=D-=�EX=���=@'�=@1�=��=.��=���=���=P� >��>i>��>���=�K�=TQ�=�j�=�0%= $/�::l����8U��N���Ѿ4��*���8�~HK�w�W���[�"�W��ZK��P8�O_ �پ�8^վlU��B�j��   �   Ń�
�Ľ��a�� �((.�`����: _=:�%F� ��4��@׀:�J�;��G<��<���<�� =jYJ=J�t=/��=M��=LM�=T�=Ol�=Ѐ�=Ԑ�=7�>��>��>cM�=�T�=��=w��=�W(= ��(�b�P3���fP���G�̾X������4�j�G�/�S��W��S���G���4�,C�7�y�о������d��   �   �^�dů��-@���{�� ?T;���;�'�;��; ^W9 �A� 2,9 	I;�K�;xf<,�<���<@�=8�F=n6p=5u�=�!�=���=	��=�2�=t��=��=�3 >���=-�=6�=�=�W�=1= [5;�bH�1u�N�B��Î������8���v�*�¹<��9H��$L��H�>�<���*�=�����p�þ64��31T��   �   f��(���q�("����;p{9<8�O< �-< ��; �=; ��� !�`7� D����9; K�;X�[<�e�<h��<.=F�J=0z=UE�=(�=�w�=���=�|�=i��=���='�= j�=x��=�˘=4j==�E<�$ ��@ɽ,-�Vg���t��Tl޾��va���+��Z6���9��6��g+���� -�Te޾�į�Ճ��#:��   �   B>���J�4菼�y;|��<X�<���<8�<(a?<�d�;�ؐ��cԻ�.���Z�im� Uc�@	9�0<׻ 1�9��<<U�<��
=�D=|�~=͎�=�={R�=*��=��=���=�Q�=��=�R�= �J=�K�<\�޼������J]�TQ������t����Uv�B����"��B�������辆����6���'^��
��   �   ǻ��8ؼ m�:<��<$��<�=LW�<�`�<8�<�A�;�4���?p�8Ƽ�o�V>!�b4��k;�(I5��L ��H��4����;���i<(8=6�L=�#�=�=�h�=��=�U�=U�=:��=?˗=��U=�&�< Fo�"x�K�뽠�5�^k{�/꡾�žOU�#���>�ޯ�g���K���������I��x�r�`N/�1$��   �   �l
��D�� ��<�=�.=�71=�@=���<�5�< �~;��=�8K��4���s�I���Ƭ�͏��(���`��X���EK���M�d���:���f�<�*=r�l=�\�=zE�=�Ŷ=� �=�O�=D(�=L�[=X��<�\8��
*��O����ȞG�؀���4��g���;�˾��׾Ɣ۾��վצǾ��R9��g,s�X#7����Y����   �   �ej�(��<��%=]R=�b=H�Y=�;= M	=���<�׺�����?��V��}�½Lv𽬛������ ��1 ��M�?��$%߽k����xV�T���ϳ;`�<�`O=���=��=�'�=��=)��=fHZ=�>=@S�;pʼx�{�l�ҽ���֧E��wr����5���|��§�����A������`^���-������h��n��   �   ��<��8=6�p=�=ꐈ=ȷ{=2gO=,�=�ac<P
7���#�z���Hؽ!�zM0��M�G�b���o�iq�Fh�6T�H|7�i���۽�����`ƺ�	�<<�8=��p=W �=���=��{=4fO=,�=�fc<��6�&�#�
��NDؽ���I0�JM�R�b�l�o��cq��h��0T�Xw7��d���۽荽���@Fź�   �   �fO=��=��=?)�=�=ϣ�=�HZ=d>=�C�;�ʼ$�{���ҽd��\�E�"|r�i����8�����>ŧ����B�������[ ^���-������n���`�j��y�<��%=FYR=$�b=�Y=,;=ZL	=���< �ֺ`����?��R����½+p���r��<� �M- �:I�����߽ܠ��hkV����� �;��<�   �   �_�=�G�=DǶ=��=�P�=�(�=8�[= ��<��8��*��R����ϡG�Â��E7�� ���D�˾8�׾%�۾!�վ�Ǿ���;��1s�4'7����dĘ��t
�` ��< �=��.=851=�>=���<05�<��~;��=��C�f4�x}s��������L������X��޴���C��D�M����`㼻�y�<�2=�l=�   �   k�=Σ�=FW�=V�=̄�=x˗=�U=�#�<HQo��	x������5�tn{�$졾žX�2����?������O����ྐ���(L��V�r��Q/�7)������ؼ�Ο:D��<���<T�=S�<�]�<d�<�A�;�,���6p���ż�j�^7!��4��a;�d>5�`A ��1�������V:��j<�@=��L=�&�=��=�   �   ̺�=b��=���=;R�=V�=�R�=b�J=�H�<�޼���1��{]��R��������9���w�ȵ�E�"�iD���s��o�農ÿ��8��z*^�.��A���K�8��ny;���<L�<���<���<P\?<�`�;�ѐ�ZԻx�-���Z� Vm�0=c��8�`�ֻ a�9��<,f�<��
='D=�~=���=�=|T�=�   �   ���=t��=�'�=tj�=���=�˘=�i==P@<"' ��Bɽ`--�Ch���u���m޾����b���+�\6���9��6��h+����.�-g޾Ư�Vփ��%:����+���u�"���;Hs9<�O<��-< ��; v=; �����@$� 9��@:;0j�;��[<$p�<��<=&K=�z=�G�=d*�=�y�=U��=~�=�   �   4 >)��=x-�=^6�=#�=�W�=�1= L5;4dH�rv�9�B��Ď������9����3�*���<��:H��%L��H�-�<�v�*�H>� �����þ&5���2T��_�"ǯ�20@����@���@)T;���;p�;@�; �V9��A� $,9�I;0S�;xf<h�<ĵ�<P�=��F=�9p=�v�=`#�="��=��=�3�=���=z�=�   �   �>ƒ>�M�=�T�=��=}��=�W(=�����b��3�� gP�Q����̾���l����4�ՍG���S���W���S��G�+�4��C����о/���^�d�f���Ľ<�a����*.�`���Ԁ:�?=:�JF���C��@̀:�I�;��G<��<���<~� =|ZJ=��t=ꂏ=
��=N�=�=�l�=\��=Q��=j�>�   �   F&>3�	>��>��=���=��=��=��= z����j�����;�������0qѾ�����A��D�B�]��Sm��U#Ӿ>���4����P� /��>ӽV����P��(�n"���2�0!P���n� -��\���l���ri�`L;�X����Gi�@�v;���<4�!=re=��=�>�=t��=���=���=?0 >�>b�	>�   �   ��	>I�>B!>�?�=���=u�=I3�=�I=phٻ�b�;�罱�7�������R;\����.w�i�|o�i���w�+�ξ�Ǫ��݆�zK������˽�f�� �E�&!����~�(���E�F�d��|�O����~�J�c�<8�P��Rp�@4;�
�<��=0+\=ߌ=x�=,|�=���=�\�=fH�=6>A4>�   �   n�>R[>�l>��=8��=��=��=Ď=`s]��aL�f�ֽ��+��Ar�>Ý�m���Pᾼ����a� ��?��,��������ɴ��g{��<������@sr��%� ��Ĕ����	(�~hG�h�`��m��j��T�f�/��1���������~<<� =�w?=��z=�#�=v˲=��=z��=���=6��=(�>�   �   P/�=�E�=V�=X�=�/�=خ�=(��=�=��:
�*�aA������3Z�A������2̾D	�.��<{��z�6���ʾ��(s���]��#��?��p��,S9�d$�,�� ȗ�P�P����ֶ6��[H�z�K���?�l�%��O������ ��pK�;D�<��=��D=�.{={˗=�|�=��=d��=[�=��=�   �   "��=���=nD�=z��=�A�=Fܬ=7��= �=�u�;.��������Q�<��\w�@+�������xž�Ҿ��վ2�оE(þe��G���G3q��9��.�Si��h�U��6��sB�@���৆��D�����kǼ������)�X�*�̚��
� Bؼd#���&� `|;xg�<(��<8�)=
�`=�V�=�=脼=��=�B�=�   �   ���=X�=@F�=���=i[�=���=ĵ}=��=0B0<@����}��\ؽ�}�VN��}�i��Z����خ�'���#٬�ӽ��ۡ���p�D�?��Y�:�Ľzo����m��Z�;��J<P�G<p��; ���"�Xٝ����v��(��$��Q#�Bl���	�@�� Ϣ�x�&���:�|l<�x�<~�2=ԅo=�L�=8��=,�=�   �    1�=�g�=�(�=�=��=�ݕ=t�k= �=�Y<��y���C������8��T%�J<K�Ʃl��.��ߊ�Z�������z���[�c�5����3�ǽ��w��N�@
Z� �q<��<x��<k�<���<ur<���;Pc�4������:z�do9�j�Q��a��h�
�d�n�T�f'7��8�����*���0M<l#�<�CC=���=<�=�   �   �w�=���=b�=C��=Yǖ=tQ�=��O=i	=�`V<�*���,���½������8�4�@	G��9Q�K�Q���H�gh6��^�� ��Q��F�d��cϼ x:�ӱ<�=�P8=��C=�l:=$i=hZ�<��<�?0;�E���ܼ��*�0�d�oԌ�K������c��t��g����㡽����~>��mҼ��u�d��<ܐ=f^=�   �   K:=�Pi=�`�=���=Z�w=�W=�Q(=l��<�<��D��r�O�!������-潁P�	����;��Ju��𽱵ĽS���P3��)���N�;���<VQ:=Vi=Pc�=ܒ�=d�w=��W=�T(=��< <������O�� ������2潔S�������(��8y����ƼĽ���D\3��=�� �;��<�   �   �Ʊ<=.K8=��C=\h:=�d=�R�<h�< 0;(E���ܼ��*��d�Xь�.���⧴�^��������ݡ�<}���q>�<WҼ �t�Ĵ�<P�=� ^=�z�=3��=��=,��=ɖ=�R�=4�O=|j	=(bV< �*���N/���½������ʯ4�BG�5>Q���Q�N�H��l6��b���������d�vϼ v:�   �   �xZ���q<���<��<8a�<���< dr<@k�;{�$���(��Ry��l9���Q���a�2�h���d�:�T��7��-�x��Pٟ�`VM<,4�<KC=(��=�>�=n3�=�i�=c*�=��=,��=�ޕ=��k=��=ؼY< �y�f�C������<��%��?K���l�1��`ኾ����u⇾k�z���[�6�����ǽ �w��^��   �    ���� /�;��J<H�G<�p�; ��("�4���������(�R$��N#��g���	���0���x�&� �:0�l<��<�2=��o=�O�=ۆ�=w	�=���=�Y�=�G�=C��=x\�=���=��}=�=`=0<����h�}��_ؽ	��3N���}�i������Wۮ������۬����𣎾0�p�}@�~\���ĽNo��   �   ��U��A��B��З��͆� W�����sǼ��~����)� �*�@���
��;ؼ���`�� �|;�t�<���<�*=f�`=�Y�=6�=P��=(��=uD�=���=��=�E�=n��=@B�=�ܬ=e��=��=�h�;(	�ސ��C����<��_w��,��j���{žҾ6־m�оc*þg�� ���B6q�9�
1��l���   �   es���W9�-�|��pЗ�|����X������6��^H�F�K�~�?�J�%�M��l���@��@j�;�L�<��=��D=�3{=�͗=�~�=��=2��=��=M �=v0�=�F�=�V�=�X�=*0�="��=)��=V�= �:��*��C�����5Z�{���+���̾���)}��\���ᾱ�ʾ7���ft��$�]���#��B��   �   麶��vr��%�l���(�����"(�RkG���`��m��j���T�>�/�0����� -���~<V� ={?=R�z=n%�=Ͳ=X�=֒�=���=L��=��>��>�[>7m>x��=���=�=�=
�=��]�@dL��ֽ��+��Cr�+ĝ�*n���Q�����b�� ��@��-�������������{��<����   �   ��˽�g��"�E�(#�����(���E��d�Z�|��O��b�~�b�c��8�`N��Mp��#4;4�<��=6-\=��=x�="}�=� �=i]�=I�=b6>�4>4�	>v�>i!>�?�=��=u�=,3�=,I=ppٻ��b�T��k�7����������R;	�<���w�ti��o����Uxﾱ�ξaȪ�`ކ��zK�q���   �   �>ӽ������P���(�@"�`�2��!P�&�n�-��W���@��&ri��K;������Ci���v;���<(�!=�re=�=G?�=Ơ�=���=&��=V0 >>s�	>T&>@�	>��>.��=���=��=q�=\�=p}��H�j���I�;�#������PqѾ*�����A��D�
B�[��Jm��L#Ӿ5���+����P�/��   �   ��˽�e��2�E�V �:����(���E���d�<�|��M��L�~���c�<8��I���Dp��?4;�<�=.\=i��=��=T}�=� �=�]�=4I�=n6>�4>D�	>��>~!>@�=[��=�u�=�3�=�J=�^ٻ��b�e��/�7����������Q;�ﾏ���v��h�"o���wﾑ�ξgǪ��݆�UyK�N���   �   O���xpr�H%��z��t���B�x(�xeG�޽`��m�"j�:�T�@�/�'����� Z�`�~<�� =�|?=��z=�%�=~Ͳ=��=��=6��=}��=��>��>�[>am>���= ��=��=��=0�=�F]��^L�h�ֽ��+��@r�e�l��nO����2a�a�*?�:+��D�����ҳ���{�8<����   �   Wn��O9�4�p��l���,繼�H��h����6�LVH�4�K���?�P�%��@���������0��; S�<.�=\�D=85{=hΗ=Z�=R�={��=.�=� �=�0�=�F�=QW�=SY�= 1�=O��=Ċ�=��= ��:�*�j>��ٯ��1Z����J���̾��R��Ty����d��c�ʾC��q����]�8�#��<��   �   h�U�p,��aB�����`��� 2����`Ǽ�������)��*�ޑ��
��.ؼ������|;0z�<��<�*=��`=HZ�=��=���=v��=�D�=��=\��=F�=(��=@C�=/ެ=U��=̆=���;�������[����<��Yw�})�������vž�Ҿ��վ��о&þc��}���*0q��9��,��e���   �   h��@?� ��;P�J<H�G<��; 3�h�!��ʝ�@��d��D$��F#��`���	�\��X���0�&�@O�:h�l<؋�<0�2=��o=�O�=4��=�	�=��=<Z�=UH�=��=�]�=G��=�}=��=�\0<����}��Wؽ�z��N�8�}�B������֮������֬�~���������p���?��V�q�Ľ�	o��   �   ��Y�	r<��< ��<�u�<|��<Ȏr<p;�"�<������Lo��c9�քQ���a�0�h���d�H�T�z7�J+������͟��ZM<�5�<�KC=���=?�=�3�=Fj�= +�=��=N��=���=\�k=��=��Y<(ay�ޤC����-2���%�B8K�\�l��,���܊�ۃ���݇�8�z�8�[�~�5�l��j�ǽ֡w��>��   �   ��<�#=�U8=2�C=rr:=o=�g�<��<��0;�D�X�ܼ�*�P�d�t͌�Ӄ������[��@��O����ۡ�`|��zp>�,UҼ`�t�D��<�=�!^={�=���="	�=���=)ʖ=tT�=p�O=<p	=؀V<Ȇ*����#'���½�������4��G�*5Q���Q�3�H��c6��Z�H������&�d��Pϼ�z:�   �   �W:=�[i=�e�=x��=�x=n�W=@[(=ܕ�<�2<`�������O�'��# ���*�?O���A������t�3��Ľ���.P3��(��`S�;ܹ�<R:=�Vi=�c�=���=px=h�W=�X(=���<-<0�����2�O��������=&潄L�ԣ�������
q��w�@�Ľ���(E3�|��P��;h��<�   �   �}�=���=�=���=�˖=�U�=|�O=�q	=P�V< �*����)���	½������&�4�aG�49Q���Q�y�H�h6��^�D �������d��bϼ 1x:<ձ<�=tQ8="�C=�n:=�k=$a�<��<��0;��D���ܼ�*�j�d�ˌ�s���à���V�����(����ա�6v���d>��?Ҽ @t��Ƒ<�=�'^=�   �   �5�= l�=�,�=��=|��=x�=��k=l�=@�Y<xfy�ƧC�w����5��%�:;K��l��.���ފ�&����߇���z�Z�[�:�5������ǽ�w��M꼀Z���q<T	�<���<�m�<��<��r<Ч�;�9컠������Zo�<b9�ȁQ� �a��h�"�d�f�T��7�N!��驼0����}M<�E�<�RC=���=�A�=�   �   ���=�[�=�I�=!��=y^�=�=ƻ}=��=�Y0<̙��x�}�,Zؽ�|�^N�H�}�������خ����	٬�����ʡ��a�p�*�?��Y��Ľo�����h� `�;��J<�G<���; �p"��Н�̟�v�, �$$�fE#��]�n�	�H��\���@~&�@A�: �l<���<�2=֓o=�R�=���=��=�   �   f��=���=G�=���=�C�=�ެ=���=��=��;��{������{�<�+\w��*��E����xž�Ҿ��վ"�о:(þ	e��>���83q�m9��.�+i���U��5��qB�����Р���?�P	���fǼ� ����p�)���*����P
��+ؼ�
����A};\��<���< *=(�`=�\�=��=���=J��=RF�=�   �   �1�=�G�=�W�=�Y�=p1�=���=���=l�= ��:��*��?�����	3Z�������
̾'	���-{��p�.���ʾ��!s����]��#��?佩p���R9��#�,���Ɨ��칼�N��F����6�YH���K���?���%��A������ ��0��;XX�<b�=��D=�8{==З=!��=��=���=x�=�!�=�   �   6�>\>�m><��=\��=�= ��=�=�Q]��_L�y�ֽZ�+��Ar�Ý��l��uPᾪ����a� ��?��,��}�����ƴ��a{��<�������sr�f%�X~��������J(�xgG���`��m�&j���T���/��(�������J���~<�� =p~?=��z='�=�β=��=��=��=D��=�>�   �   a�	>��>�!>5@�=w��=�u�=�3�=�J= `ٻ�b���罀�7��������Q;R����+w�i�|o�h���w�)�ξ�Ǫ��݆�
zK������˽�f���E�� ����@�(�v�E�ȿd�D�|��N����~���c�d8��K�� Hp��74;��<.�=z.\=���=�=�}�=�=�]�=�I�=�6>�4>�   �   }�>`z>Fu>N>�-�=B��=Kۨ=t�o=<��<�λ�zB��y��}���eI��H}��ѕ��0������������kn���Ж��:��T��A'������>½&�����񱆽Rv��>]�����s���Y�!���%���!����t� ���νH��6W1�0�i��V< `=b�u=�ޡ=W�=\��=\��=��>T�>�|>�   �   F�>5f>�o>�T >�_�=|�=Ү�=�on=t��<�/���=�(#��X���BE�|x���W����D��-2��?,��JŤ��l���[|�*�N��"������6������~�����
"��⓲�Qٽ�� �J��m~���!�z�����aS��u�ʽ�j����.��_j���L<�J=:9p=.Ǟ=m¿=�A�=S{�=6S>�v>5>�   �   �>7>�I>(��=6��=�5�=��=�Mj=���<ځ��(.�}ׯ����ld9��Ci���i˚�򆥾��A��Z)������êj��4?��*�O��æ�y(��~�[� �]�����Kٞ��Ľ9�����g�<#�`����"��jO��GK��j)�p�p�Р,<�1
=�n_=�7�=է�=��=���=�p�=h7>PR>�   �   �>�M>x��=rQ�=�!�=���=m��=,�a=��<@����&��ŝ�%���a'���R��x�~��h�������� ���*�t��O�!�&�W  ��"��������E��>$��u&��G���UƢ���ƽ(��կ���0�,y�؆�}�սXۮ�����`#��Ä��;��<LA=i�=��=a��=���=���=x��=x� >�   �   ���=r��=w��=R�=$��=	J�=���=�qQ=Hg�< �L���J����սԠ�0�6�X�W�$�p��H���V����|���i�:�M�t3,��*��ʽ�����=;��]��x���X��� l��lA1�zPq��5��g���Z�ϽC<ܽ��ܽ�Pѽ,A��G؜��gq�h�"�pʣ���	�4��<��=0@V=��=��=d��= �=��=�(�=�   �   ?G�="��=UJ�=S�=^��=���=#�=�7=�ؾ<�����:�B�l��ε�m������]3��UG�^�R���T�\�L�)w;�Ě"�`����ʽ�덽�1�|�������z4��^���%� ��n����P�����j:��/����7��g%���R���Y��n*h���.�@W�@C���};���<�=�L=hy�=�=��=Dl�=��=�   �   �ܾ=���=k^�=���=d�=���=FT=�o=���<�1��h�޼h�P�mJ��t˽����J����� %��$�6����� �뽹k���>��ng�y����:��V<(�<��<`[=<�͢:�GB��Pּ>6$���U��{�؉�Hv���O��J��r�n�`�L��q$�l켸������^H<�]�<�.=��h=�Ԏ=��=;	�=�   �   ��=��=Q�=��=��=h�P=|=�^�<�;��J��\��0>E����٨�XǽmA߽��#���l�r�ڽއ�������tR���켰����7<�S�<="h"=Je=�3= ��<P9<��������؄(���N�`�k�8R��ф�W~��`���~�q���U�2G/�P����m�� �V�Ц�<�
=J�A=�tv=�B�=�   �   6h=FAu=$p=��Y=5=�=��<0��;r(���ȼ�o�F�M��!{�ߐ����婽�8���ب� ������*`S�vU��h�� va;L;�<�=�CH=h=�Fu=�p=D�Y=�5=P=�)�<`��;�_(�`�ȼDm���M�#{�ᐽ�
��-驽�<��Jݨ�;
��߷��~jS�X_��z����`;$,�<,=�=H=�   �   ��=b"=>_=Z-=8��<��8<�2�x���d�򼪉(�Z�N�d�k�zR�ф��|��ʐ��؝q�&�U��>/������[����T�ض�<�= �A=�zv=�E�=:�=/��=��=�=0�=<�P= =8g�<p��;�xJ��Z���>E�D���Nۨ��ǽ�E߽y��)���r�[�ڽ����	����~R�л������}7<@F�<�   �   �V<���<d��<PA=< ��: dB��^ּ=$�\�U���{�Aډ��w��yP���I��d�n���L��l$�(��������(|H<0l�<�.=�h=�׎=���=��=G߾=���=�`�=���=n�=���=�IT=�r=P��< (����޼:�P�FL���v˽������F��%%��$�c��������q���C���o�4��� @�:�   �   ����4� h^���%��(������P�"����=��7���:��E'���S��9Z��t)h�N�.��O���B��/~;0��<�=��L=0|�=��=�=pn�=���="I�=��=	L�=�T�=���=��=V$�=7=l۾< ����<���l��е�������E`3��XG�x�R��T���L�Bz;���"����u�ʽ��1�����   �   Ti�������xx���G1�NWq�M9��ݘ����Ͻ7?ܽ~�ܽRѽuB���؜�ngq��"�@ţ��
	�\��<�=�DV="�=�=w��=��=B�=T*�= ��=���=ά�=��=Y��="K�=v��=�rQ=Hh�< &����uL��V�սr��<�6�ǎW���p�+J��WX����|���i���M��5,�$-�׳ʽ���D;��   �   �F��C$�{&�R�G����Sɢ���ƽ/�潶���2�Dz�����ս�ۮ�����V#�����.�;@��<ZOA=�j�=��=��=��=G��=���=� >��>IN>q��=`R�=}"�=X��=���=؇a=��<����r(��ǝ�S'��@c'�z�R�.�x�I������]ᗾF���\���p�t��O���&��! ��%��G����   �   c*��^�[��]������۞�#Ľl;�$���h�4$�* �����콭O��%K��|)�8�p���,<4
=,q_=$9�=��=��=���=�q�=�7>�R>|�>�>J>���=���=Z6�=��=�Mj=D��<����d*.��د�����e9�Ei�����O̚�凥���4��@*������?�j��5?� ,�l��Ŧ��   �   Ȼ���G���z#��a����Rٽd� ������!�������S��Q�ʽ�j����.�HZj��L<hL=�:p=Ȟ=>ÿ=~B�=�{�=�S>�v>T5>~�>jf>�o>�T >�_�=��=���=pn=���< 5���=��#������CE�Px�_Ò�ڽ��%E���2���,���Ť�Am��v\|��N���"������7���   �   ������������v���]�����^s�6��q�!���%�u�!����+� �-�ν����U1�p�i�@V<4a=l�u=8ߡ=��=���=���=�>n�>�|>��>uz>Wu>N>�-�=F��=Bۨ=V�o=���<0λJ{B�Ez������eI��H}��ѕ��0������������on���Ж��:��T��A'���� ?½�   �   "����������!�������PٽV� �ߴ��}���!����ؕ��Q����ʽi���.��Qj���L<�M=�;p=hȞ=�ÿ=�B�=.|�=�S>	w>`5>��>yf>�o>U >6`�=
�=d��=2qn=��< $��.=�G"�����bBE��x���켤�(D���1���+���Ĥ�bl���Z|�}�N�b�"�����)6���   �   7'��T�[���]�����!؞�eĽj7� ���f��!����|���IL��?H��� )�@�p���,<�6
=s_=�9�=���=^�=��=�q�=�7>�R>��>�>:J>��=9��=�6�=��=>Pj=p��<����,%.�vկ����"c9�<Bi��󉾉ʚ������Q��r(��ꖉ�A�j�C3?��)�z�པ����   �   ��E�z;$�xr&�j�G�:�� Ģ�0�ƽD�潎����.�@w�҂�\�ս:׮������#����PR�;4��<
RA=�k�=\�=���=���=���=��=9� >��>tN>ҧ�=�R�=$#�=<��=,��=�a=4!�< ��6!����!���_'���R���x��|������ޗ���ޫ��ڒt��O�P�&�� � ��l����   �   �S��x�x����b��d<1��Jq��2��ʑ��K�Ͻ�7ܽD�ܽ�Kѽ,<��FӜ��]q�̬"����������<F�=<GV=#�=��=��=P�=��=�*�=w��=9��=<��=,�=��=2L�=���=�vQ=�r�<�w�P���F����սk����6�v�W��p�G��4U����|���i�u�M��0,��(�=�ʽh���l8;��   �   Xv��'4� �]�P�%���������P�r����5��<���C2����� M��0T��h��y.��AἈ�B��x~;(��<��=��L=�|�=C�=��=�n�=P��=�I�=R��=�L�=RU�=θ�=D��=�%�=L	7=��< ����)�xl��ɵ�������Z3��RG���R�N�T���L��s;���"���� �ʽ`獽j1�,����   �   HW<0�<Ȑ<Xr=<@��:8,B�$Aּ~-$�>�U���{�\҉�cp���I���C���n���L�Re$�p�����`g� �H<8p�<*.=:�h=T؎=&��=�=�߾=��=a�=���=J�=�=�LT=w=�	�<@왻x�޼.�P��D��(n˽����������%�Y~$����E�����/f���9���^�Lj�����:�   �   �=�m"=�j=Z9=���<�#9<�M�l}��l��*z(�L�N�.�k�tE�:˄��w�������q���U�B:/������V�� 5T�แ<=��A=�{v=�E�=��=���=J�=��=�=��P=$#=�o�<�ߤ;\J�lH��L3E�A����Ҩ��ǽ�:߽�����e��ڽt��������iR����P{���7<t`�<�   �   � h=BLu=p=��Y=�5=!=9�<� �;`9(�x�ȼ�a�f�M�{�@ڐ����᩽�5��
֨�#������]S��S��e����a;�<�<�=�DH=�h=�Gu=�p=l�Y=@5=f=t/�<�ڐ;XK(�T�ȼ�d��M�P{�oِ����Tߩ�32���Ѩ�����b���ZTS��J��T�� b;�J�<� =�IH=�   �   ��=���=H�=��=�=��P=.'=0w�<`��;0QJ��D���2E�ⶆ�zԨ�oǽ">߽���i!��Ak�$�ڽ↼�Ӣ��^sR�ħ켐�����7<�T�<�=�h"=f=�4=���<�9< ��|���P��&(���N�<�k�G�>˄��v��׊���q�V�U�3/�lu��G�� MR�Pȁ<�=��A= �v=IH�=�   �   ��=��=�b�=*��=��=Wć=PT=�y=��<�ޙ�`�޼ �P�$F��Pp˽�������m��B%�C�$����4��c��@k��^>���f��w��@.�:�V<P�<l��<�^=<��:BB��Lּ�3$�N�U�B�{��ԉ�wr�� K���D��ƽn�"�L�(b$����$����	���H<�|�<%.=��h=�ڎ=h¤=�=�   �   K�=���=�M�=�V�= ��=���='�=d7=��< ����*缼yl�G˵�g���^��\3� UG���R�O�T���L��v;���"�2��w�ʽ?덽1�����Њ��r4���]��%�p��L��L�P������8��M���5��Z"��O���U��B h�Ny.�x>���B���~;���<>�=tM=4�=i�={�=�p�=���=�   �   ���=R��=L��=0�=��= M�=�= xQ=Xt�<�n�$��H��_�ս���9�6���W���p�qH���V��o�|�l�i��M�V3,��*�үʽr����=;��\������t����j���@1��Oq�A5������E�Ͻ�:ܽ �ܽINѽ]>���Ԝ��_q���"�|����d���<�=bJV=�$�=o�=���=��=��=�+�=�   �   &�>�N>���=�S�=�#�=���=���=�a="�< ��4"��Ý�@#���`'���R���x��}��=����ߗ�������t��O��&�B  ��"��~���d�E��>$��u&���G�����Ţ�N�ƽ������G0��x�6��z�ս�خ�誁�#�D����S�;��<�SA=�l�=c�=���=���=���=���=�� >�   �   ��>�>pJ>���=���=\7�=��=�Pj=���< ��%.�.֯�>���c9�HCi���I˚�؆�����3��R)��������j��4?��*�9���¦�b(��R�[���]�q���#ٞ��Ľ�8�����g��"����t�����M��I��h)���p���,<�6
=�s_=J:�=$��=��=���=tr�=<8>S>�   �   ��>�f>�o>"U >b`�=5�=���=�qn=���<�#��b=��"�����BE�Gx���I����D��&2��;,��FŤ��l���[|�$�N��"������6������j�梀��!��ȓ���Pٽ�� �2��T~�j�!�G��t���R����ʽj����.�PWj���L<M=�;p=\Ȟ=�ÿ=�B�=N|�=�S>w>v5>�   �   �>��>r:	>>�9�=5��=^þ=nA�=]]=3�< hf:����C#��OBɽ"T��6$��;�!�J���O���J�H�<�V'��0��N齒g��bЛ��K��*֐�ct��ؽg7�d	0�n�V��y{��̌�ѿ���@�����p���n,y�S�P�i�#�"M꽤ď��� ��;�=-:�=�=��=el�=�;>�	>?�>�   �   ��>t�>��>Z�>!c�=��=C�=З=*{Y=b�< �H:d���;ǀ��^Ž���|� ��7�?F��K���E���7���"��
���R���/k��� ��v����ͣ���н�
��F+�c}Q�	�u�����(m���떾����v����t�6�L�Bm ��o�8����@�PZ�;�!=�=���=-�=�J�=l#>�>��>�   �   �p	>0�>�>P�=$��=��==�6�=R&M=(=�< �?9���4�t��w������"��	�+��9�I=�Y�7� �)���������˽�w���ɂ��Ph�\�p�nr���K������v���A�$Sd��\��P҉��P���R������1e�@U@�J���׽���P%׼0Q <�w=�+�=���=��=J��=���=P�>�Y>�   �   �`>�>6��=���=���=��=M�=!��=�t6=�< U̺l��4�c�E̪�������.
�B�$�<�'���!��m��T��3ֽb\��9��xK���/�<�7� !d����)�Ͻ��Q�)��I��d���u�s�|��Ex�?h�I�N�Z�-��n�OFý8kn��*��h�<z=��q=ZM�=�b�=��=n�=�u�=bt>�   �   �1�=L��=�F�=(O�=h^�=ͫ=�=�[=�_=���<@����.VT��љ�SBƽR콫[�N�B������IϽl���#{�J�3�� �X�μ܇ܼ�A�]��p����ؽ��
�x�'���?���P�,�W�U�P(H���2���w��^���T�PY����;�� =(zY=é�=�T�=,��= 9�=D��=i��=�   �   ���=|��=��=�޼=kR�=���=��`=I!=�P�<���;OU����d�M���������G�ǽR�ڽ�w��7�uѽ>H���ە�\@a�|������(E)� ����л`Dt����~�P��暽|gн���7���L'�K/�|W.�cL%�6�ѳ��̽G��p?��s�� f2;d+�<p�4=�i{=T�=�!�=���=T��=%�=�   �   ���=:`�=�>�=|?�=�T�=�UM=�=��<�_�; =,�d#ϼ�X!��VW������`���~������ů�²��͌����t�&�5�����@�@h ;��A<�<(�}<0$<�A�������T4��������u�ܽ�p��F��Я�|��&��pҽͭ�}{���w7�T�ȼ 띻��c<\� =<�B=�}=t�=v��=$��=���=�   �   ��=IK�=ݠ�=(�`=��*=���<Pd4< ё�hS���F1�t�W�� v�����ތ�ӎ��\��S߁�|d��8�İ��*��@����U<|��<��
=nd=N=�$ =|��<�Ϧ;�TU��j���T�㍽ڐ���2��0�ǽɋǽq]��$ح�����^3{�6�A�b���O�� ����3o<���<��4=tHh=�=�{�=���=�   �   ��n=�CZ=��4=F =��<��������:lF�^
t�\(��ᆓ�ꎖ������k��鄀�"5a�f�9���
�������ֻ�C<���<n(=�A=
�`=8�p=��n=�IZ=��4=�M =��< ���0�������cF�nt��$��=���!���"����k�������8a�h�9�j�
��ª���ֻ�(<�v�< "=zA=0�`=`�p=�   �   �=� =��<`��;XxU�@t���T�荽ו��37��J�ǽ#�ǽ�_���٭�����2{�ΛA��~�F�� 蓺�Jo<���<F�4=Nh=��=�~�=g�=È�=N�=ߣ�=�a=��*=D��<@�4<0���8E�����@1���W���u�����ߌ��Ԏ��^��d⁽zd�(8�J��`9������x�U<l��<v�
="^=�   �   8g}<�<p����ͺ��^4�闈����� �ܽDv�������l����rҽ$έ��{��bv7� �ȼΝ�d<� =�B=��}=���=ƿ�=c��=D��= ��=�b�=xA�=6B�=�W�=�[M=�#=���<���;H*,�$ϼ~V!�*VW�S���
b��̀���ï��ȯ�����א���u��5���㼸�@����:ȻA<���<�   �   ��л�`t����2�P��뚽�lн������O'��/��Y.�kN%������d̽����o?��p����2;2�<&�4=�m{=Q�=�#�=���=9��=
�=���={��=2��=�=�T�= ��=��`=�M!=�X�<�ت;XFU������M�����p�����ǽ��ڽ�{��;ཛྷ
ѽYL���ߕ��Ga����L����^)��C���   �   d�ܼ�H�0�]��t���ؽ�
� �'�C�?���P���W�IU�>*H�:�2���ܴ�����T��V���"�;P� =}Y=P��=jV�=���=�:�=І�=���=&3�=���=H�=�P�=5`�=�Ϋ=��=b\=Fb=���<`���輄WT��ҙ�dDƽ�T�E]��O�0����f
�UMϽ�o��l*{�r�3�� �t�μ�   �   ��7�'d�k�����Ͻ"����)�c�I�Dd��u���|��Gx��@h���N�D�-�Vo��Fý$kn�)��Ѝ<|=ܬq=�N�=4d�= ��=��=�v�=�t>{a>��>q��=���=<��=P��=��=;��=`v6=T�<�I̺����c��ͪ����
������$��'���!�fo�|V��6ֽ,_������K���/��   �   ��p��t��[N�������w���A��Td��]��,Ӊ�TQ���S��7���2e��U@�����׽����@#׼W <xy=�,�=���=��=0��=ޚ�=��>/Z>Iq	>��>">.�=��=��=���=[7�=J'M=8>�< �?9��ºt��x��!�����&�+��9��=���7�\�)�"��D����˽�y���˂��Th��   �   ����^ϣ���н���G+��~Q�.�u�F����m��k얾�����6t�G�L�,m ��o彞����=�Pf�;\#=��=h��=��=�K�=�#>f�>��>:�>��>��>��>�c�=��=��=^З=�{Y=,b�<��H:�����ǀ��_Ž(��� ���7��?F�K���E�<�7�{�"�F
�6�ὁ���il���!���   �   �֐�2u��ؽ�7��	0���V�z{�
͌�俖��@������J���,y���P���#�L꽧Ï�� �0��;.!=�:�=z��=Z�=�l�=�;>�	>Y�>�>��>�:	>>:�=E��=bþ=kA�=�\]=x2�<�Qf:h����#���BɽJT��6$�/�;�=�J��O��J�\�<�V'�1��N��g���Л�CL���   �   T����ͣ���н�
��F+�&}Q���u�r����l���떾���ᓉ��t��L�
l ��m����9�pu�;�$=g	�=���=- �=�K�=�#>x�>��>F�>��>��>��>�c�=���=��=�З=�|Y= e�< [I:����Wƀ��]Ž"��� �n�7�~>F�%K�N�E���7�E�"�,
�5�ί����j��D ���   �   p�p��q���J������Yu���A�Rd�\���щ��O���Q������/e�HS@�l��o�׽۽��׼he <2|=�-�=^��=v�=���=.��=ۊ>KZ>dq	>��>A>z�=^��= �=V��=.8�=v)M=�C�< vC9��8�t��u��D��������+�m9��=��7���)�ش����E�˽/v���Ȃ��Nh��   �   �7��d�V����Ͻ���؝)�Y�I��d�~�u� �|�@Cx�v<h���N�ͥ-�\l��Aýcn�(���<N=��q=�O�=�d�=���=�=.w�=u>�a>��>���=d��=���=���=b�=^��=ny6=0�< �˺��$�c�ɪ�H����Q�b�$�^�'�-�!�l�TS�1ֽ�Y��	���K� �/��   �   Pܼd=��]��m��Q�ؽ��
�J�'��?�4�P�6�W���T�&%H���2�����������S��G���R�;�� =��Y=���=aW�=v��=8;�=:��=J��=|3�=6��=�H�=WQ�=�`�=�ϫ=��=\=�e=��< ݴ����JNT�|͙�>ƽ�M�^Y��K���l��\��EϽ�h���{���3�  ���μ�   �   ��л�/t�����P�'㚽7cнr��s���I'�/�T.��H%���,����̽^	��e?��_����2;<�<��4=�p{=`�=c$�=��=���=q�=.��=ޱ�=���=��=dU�=ݝ�=��`=�P!=�`�<��;�+U�n����M���������$�ǽ�ڽ�r㽿2཈ѽ�C���ו��8a��������/)�0硻�   �   ��}<p:<0��쮺�(M4�?���������ܽzj�����H�������iҽcƭ� u���k7�$�ȼ�����!d<�� = �B=�}=���=d��=ℹ=���=f��=c�=�A�=�B�=<X�=�]M= &=��< ��;p,��ϼ4N!�
LW�K���[�� y��&�������k�������8�t�P�5����x�@� � ;H�A<��<�   �   �=D* =��<��;05U��a�\|T�Tݍ������+��@�ǽ��ǽQV��ѭ�����*&{���A�|v�L9���J���Yo<$��<`�4=�Oh=L�=�~�=��=)��=N�=L��=�a=ʉ*=���< �4< ~���=�����:1�W�6�u�����،�N͎��V���ف��d��	8�V��H�����V<,��<�=�i=�   �   ʰn=ZOZ=j�4= T =�'�<������������WF���s�^��r}��<���:퓽#e��I���+a��9���
�����P�ֻN<���<�)=�A=��`=��p=D�n=�JZ=F�4=nN =�<�{��H�����$`F���s�"������������e��4��*a�آ9�l�
������{ֻ d<���<
/=�$A=��`=~�p=�   �   /��=�P�=���=�a=Z�*=���<H�4<pG���/��H��41��W���u�����،�$Ύ��X�� ܁�td��8�έ�&���ൺ��U<t��<��
=e=�=>% =���<0֦;�PU�^i�ڄT��፽[����0����ǽ��ǽ�Y���ӭ�Y����'{�l�A��t�t3���Ӓ��jo<��<��4=�Sh=o��=	��=��=�   �    ��=�d�=�C�=�D�=�Z�=�bM=�+=��<ך;�,�`ϼK!�4JW�)����[��xz��c���h¯�����4���l�t�N�5��� �@��u ;x�A<4�<8�}<H&<0=��L���,T4�;���l�����ܽ�o��|��ʮ�2������lҽ�ȭ��v���l7���ȼ���� +d<�� =b�B=��}=n��=$«=���=^��=�   �   ���=X��=;��=8�=@W�=៍= a=�T!=�h�<p�;� U����b�M���������ǽ��ڽ�u�=6�9ѽQG��-ە�P?a���������B)�0�� �л�Bt������P��暽gн�����KL'��/��V.�`K%���Ӱ���̽^��~g?��a����2;�>�<��4=s{=��=�%�=|��=��=��=�   �   �4�=^��=J�=�R�=6b�="ѫ=v��=0\=�h=���<�δ���缈NT�=Ι�g?ƽ�O콬Z�JM���.���� IϽ�k��J#{���3�x ���μ4�ܼvA�`�]�wp��F�ؽn�
�L�'�O�?���P���W�lU��'H���2���ְ�a���& T�TK���L�;&� =~�Y=L��=9X�=b��=2<�==��=P��=�   �   �a>�>���=M��=���=
�=x�=m��=X{6=\!�<@�˺d�似�c��ɪ�������y	���$�ϥ'���!��m��T��3ֽ+\����.K�@�/��7�� d������Ͻ���2�)��I��d���u�&�|�uEx��>h���N���-��m�2Dý�fn�� ��X�<�=�q=�O�=re�=C��=��=�w�=tu>�   �   �q	>��>�>�=���=��=��=�8�=�*M=�E�< D9ě켰�t�5v��:��������+�_9�
=�*�7���)�ٵ�����ٿ˽�w���ɂ��Ph�,�p�Zr���K������v���A�Sd��\��>҉�qP���R�����z1e��T@������׽�����׼�^ <6{=y-�=T��=��=���=s��=�>xZ>�   �   R�>ϫ>�>Ƨ>d�=��=F	�="ї=V}Y=@f�< vI:����]ƀ�^ŽT��9� �Ы7��>F��K���E��7���"��
���B���"k��z ��l����ͣ���н�
��F+�\}Q���u�����!m���떾����d����t���L��l �Ho�|����=鼠g�;�#=��=���=��=�K�=�#>y�>��>�   �   F@>��
>*E>�p>��=�>�=�}�=`ګ=2[�=R=�C=P�A<�,�����Q��&��UJ��%���v���i���«��j��0��ڗ[�:�K��uZ��c��_F��J �t$2�zk�1/��Z紾�Ѿ�j�{������a���NB龳?Ѿ�����(����\����幽Ԑ����;W-=Px�=Z��=r��=Ο�=�n>��
>�   �   E >�y	>�>j)�=���=H��=���=�b�=�!�=��J=XN�<�q0<p=%�(����N�1[��g]�����G���%��۵���w���Qt��zP��@��(O�#K���_�����"R-�X�e� ʑ�*�����;k�侯��b���k��_��
;`i���7���<X���`��f{��!�;P�.=LB�=b+�=���=��=�>��	>�   �   3>�>�� >���=d��=Z��=�B�=߮�=6/v=�33=$��<�G�;�B�����"�F����.L���L��{���+���R����~���R��#0�
� ��8.�a�K��Ni�VQ��U��[��������־�@德Z�S��Z׾�&�����������J���%q��tM�XY<<]1=;]�= ��=���=�U�=�>��>�   �   �� >�D�=$3�=���=>��=7�=���=��=�iH=��	=|��<�L�:'�������=�p��2��)��������X���Ss�ZaI�� �����4�ܼ$����1)���흿�An	���:��.q�!������{l���ξ�ӾŊϾ��¾h����E���q�I�6�����y���ڼЕB<��3=��=ؠ�=n��=���=���=�� >�   �   O��=���=d��=;�=r��=�=~�u=rS==��=�F�< (�;@������Z�Xc9�R[���p�zNw�6n�z�U�U1�d��L����s�`�7�p�_��ü��.�>��� ۽.���HJ�Z1{�i���X���|���+���峾X�� ���F����qQ������׽@\v�HC��8Uq<^Q3=�+�=Rw�=D�=A:�=���=6�=�   �   ��=�n�='s�=?��=�7�=��R= �=8i�<�!<`�y�@Y{�DeѼ����T*��f@��M��P�ΦG��2���@�Ҽ��t�����GB;�R�;p��;@{w�� ���6�
ԛ�	���p�x�H��	p��	��;ߒ�e��I-�������|��-X�R�.�y���{���G�x�c����< B,=��=Q7�=�;�=���=0j�=�*�=�   �   �u�=���=���=�.e=�%=���<���;ؚ��沼�/�f�,�z<F�D�U�B\�ڀY�H�N��;;�^������?���c��mS;O_<,o�<ȡ�<�:�<�4�<��s;�ى�и2��z��������f,6�~�Q���d�Y�m���k�bJ_�$�I�N\-�:��̑Խ�F���*�F#�lۀ<n�=zeh=%�=�L�=���=H��=7��=�   �   �W�=�Sw=j�<=p�<��<�Q(����*1?���x�Y��������!c��E����^@c�{6����t��� ĻP��;�<�> =�R"=5=��4=��=��<`�.<��<�������Ľ,������&��/�T�0���(�>��
��`ܽ	�����i� ����h$E<L)�<>BB=Cy=lA�=75�=�Ţ=���=�   �   D�M=�Y=L��<�@1��~׼�N�����h���Dݽ����P��������/ɽ}7���}���E��!���CJ��C�;8��<v6=<�A=�f=�|=-c�=.q=
�M=�a=虙<��0�@h׼��N�Q���a���=ݽ���J��������ɽV5��a|����E��#��PMJ��(�;X��< 2=��A=2�f=��|=j`�=$yq=�   �   p��<�t.<P�<���L���ؒĽ���������&���/�ԋ0��(��@���qcܽ����*�i���� ��.E<�/�<�EB=Gy=�C�={7�=FȢ=J��=�Z�=fZw= �<=��<`�<'(�o�%?��x��{����������_���B��#�t?c��{6���$����5Ļ0��;,�<r9 =�M"=p5=��4=�=�   �   �ms;p뉼�2�������Ὂ��h06���Q���d�n�m�N�k��M_���I��^-�ܹ��ԽH��\+��B#�߀<�=zhh=��=�N�={��=h��=���=\x�=���='�=�5e=�%=$��<�D�;(u�Բ�'��x,�6F�h�U� \�~Y���N��=;�j�����,I���w� S;H9_<�c�<��<�.�<'�<�   �   $0���6�6ٛ���,t�D�H��p����_ᒾg��6/��΄��d�|��/X��.���� }���G�@�c�p��<D,=���=�8�=@=�=���=�k�=�,�=,��=:q�=�u�=6��=<;�=��R=p�=�w�< >< -y�xB{�$\Ѽ����R*��f@�h�M��P�l�G�b�2�~���Ҽ8u��C����A;�$�;@��;@�w��   �   �.�����%۽���KJ� 5{�]���Z���~���-��a糾���v���U���XsQ������׽F]v�C��Yq<�R3=�,�=wx�=RE�=�;�= �=�7�=��=���=z��=a=�=���=��=�u=�X==2�=tP�<�G�;H��읹�zY�d9�4[���p�LRw��n�T�U�2Z1���������s��7�x`��%ü�   �   n������zp	���:��1q�����y��>n����ξ��ӾI�Ͼ�¾�����F���q��6���������ڼx�B<V�3=��=ơ�=n��=���=��=5� >^� >,F�=�4�=���=��=,�={��=��=6mH=֖	=���< ��:d%�������=�p�4��񸓽����[��2Xs��eI�j�������ܼ`���f7)��   �   �M��pl�(S��U�B򇾣���'���r�־�A��[�e���Z׾d'��[��޾���J�2��	q���L��]<�^1=�]�=얽=r��=�V�={�>�>z3>>>� >���=���=���=�C�=��=r1v=�53=��<�N�;B�����P�F�����\M��@N���|��e-��@T��(�~�&�R�0'0�Ξ ��<.��a��   �   �a��E���lS-�ӹe��ʑ����[�;=��o�������󾽧�F;|i���7��<X��������y��-�;.=C�=,�=G��=��=0�>=�	>� >z	>f�>*�=^��=���=���=dc�=/"�=V�J=tO�<�r0<(>%�4����N��[��(^������H���&��ܶ��y���St��|P���@��+O��L���   �   lG��� �)%2��zk��/���紾a�Ѿ�j龗������D���B�h?ѾK���](����\����乽����ȿ;�X-=y�=���=���=0��=o>��
>b@>��
>FE>�p>�=�>�=�}�=cګ=+[�=�R=�C=�A<�����t�Q��&���J��g����������9ë�%k�����Ƙ[�R�K�RwZ��d���   �   �_��/���1R-�Y�e�ʑ����=�;��'�������󾋦�-;�h���6��";X�������Dw�P=�;D�.=�C�=s,�=���=��=G�>L�	>� >z	>t�>.*�=���=#��=���=�c�=�"�=Z�J=R�< y0<X6%�|����N�SZ���\��8���F���$�����Ww���Pt��yP���@��(O�1K���   �   CJ��wh��P��U������������#�־�?�wY���復X׾P%�����K���w�J����m���G�m<pa1=_�=���= ��=W�=��>;�>�3>>X� >��=��=���=XD�=���=�2v=�73= ��<�g�;B�����"�F����/J���J��?y��*���P��ʋ~��R�h!0�&� ��6.��a��   �   ���5���4m	���:�>-q�������k��l�ξ*�Ӿ��Ͼ��¾����>D���|q�|�6����9	��t�ڼȮB<R�3=
�=ڢ�=4��=<��=}��=a� >�� >nF�=�4�=���=s��=��=��=v�=VoH=��	=���< �:��������=�	p��/��O���㡓�WV���Ns��\I����������ܼd����.)��   �   x�.�؝��/۽j���FJ��.{����W���z���)��p㳾3�����O���-nQ�J���׽ZRv�(2���rq<�W3=�.�=�y�=>F�=D<�=� �=�7�=^��=��=���=�=�=i��=J�=x�u=�Z==��=�V�<�h�;�m�����R�x[9��[�:�p�DGw�Jn���U�O1����T��� �s��7���_�8ü�   �   ���4
6��Л���In���H�jp����ݒ��b���*��ˀ��	�|�R)X�r�.�����u����F�h�c�l�<NI,=���=':�=I>�=^��=�l�=!-�=���=�q�=3v�=���=�;�=��R=�=|�<�H< �x�x0{��PѼ����J*�V]@��M��vP�n�G�}2�.���Ҽ��t�`Ꝼ��B;�x�;`ݠ; 1w��   �    @t;h͉�x�2�?v��ʱ὿���(6���Q�l�d���m���k��E_���I�X-�D����Խm@��N�X#�T�<T�=zlh=N�=�O�=F��=���=���=�x�=��=��=�6e=�%=���<@Q�;�l��β��#�&t,�d0F���U� \�$vY��}N�R2;�F�����0���F�@�S; g_<$z�<���<�D�<�>�<�   �   @��<��.<H�<�"	�ᗈ��ĽOx��;����&���/�ԃ0���(��9�d��Xܽ�񨽬�i�P����� JE<$:�<�IB=�Iy=�D�=C8�=�Ȣ=���=7[�=[w=��<=h�<0�<h"(��k�#?���x�.z�������|\���>���섽p5c��p6�j������0�û`�;<(�<�D =tX"=0 5=��4=��=�   �   l�M=�g=짙<�0��T׼~~N������Z��:6ݽ
|�zB��Y��P��	ɽ�-��pu��حE�`��x"J��u�;м�<:=�A=��f=D�|=�c�= �q=��M=Tb=8��<@�0��f׼��N�����`���<ݽ����H��N����qɽG1���w����E����@!J�p��;@��<�<=��A=X�f=ґ|=�e�=(�q=�   �   N]�=�_w=��<=�"�<�<8�'�TX�?�x�x��t���G���TX��c;��7ꄽ`2c��o6����������ûp�;<!�<�@ =�T"=D5=��4=R�=d��<��.<@�<�6�����u�Ľ�~�����O�&�a�/���0���(��<�	�]ܽ����i�ұ� ��xKE<�<�<�KB=bLy=�E�=�9�=�ʢ=���=�   �   �z�=, �=���=|<e=J#%=T��<0��;@J�ȼ�����k,��(F�V�U�8\��rY�z|N�T2;��������6���U���S;�V_<�q�<ܣ�<x<�<6�< �s;�؉�J�2�Wz����ὢ��-,6�6�Q�`�d���m���k��I_� �I�[-�ȶ���ԽBC��#��%#���<��=�mh="�=�P�=|��=d��=���=�   �   ��=Fs�=,x�=笠=V>�=��R=j�=���<�d< �x�p{�FѼ����G*��[@���M��wP���G��2�����ҼH�t���� YB;�Y�;���;�rw�����6��ӛ�Ը车p�W�H��	p��	��ߒ��d��
-��Ȃ����|��,X�-�.�,���x����F�@�c�H	�<�H,=М�=�:�=�>�=B��=�m�=a.�=�   �   t��=R��=T��=�?�=n �=��=\�u=�_==��=�`�<���;�^�����BP��Z9�[�ʋp��Iw�zn���U� S1���� �����s��7���_�0üZ�.�����۽���HJ�E1{�[���X���|���+��f峾��ְ��뙁��pQ����a�׽~Wv�<9�� jq<�V3=�.�=�y�=�F�=�<�=X�=�8�=�   �   � >TG�=6�=��=��=<��=՘�=@�=�rH=��	=���<�_�:H�����j�=��	p��0��~���Y����W��PRs�>`I�$ �����0�ܼx���X1)����ҝ��1n	���:��.q�������pl����ξϯӾ��Ͼ��¾7����E��q���6�u�������ڼ��B<��3=�	�=���=T��=���=��=�� >�   �   �3>^>�� >���=ǟ�=���=kE�=ӱ�=<5v=�93=���<0t�;pB�����(�F�m����J���K��Oz��!+��R���~�4�R�B#0��� �L8.��a��J��:i�JQ��U��U��������־�@徬Z�A���Y׾�&�����Y���C�J����p��*K��b<�_1=w^�=]��=���=W�=��>`�>�   �   � >+z	>��>x*�=���=���=[ �=>d�=&#�=z�J= T�<�|0<p3%������N�`Z���\�����ZG��[%�������w���Qt��zP��@��(O�K���_������R-�V�e�ʑ�(���}�;h�侬��^���c��U���;Qi���7��v<X�������Dz�0+�;��.=�B�=�+�=C��=��=:�>L�	>�   �   �8>��>�>b�=J%�=1:�=�)�=�c�=?�=��}="{K=(�=���<�{G< ��:8U	���|���������L��+��0lq�p��G���y �j�Z�d��N��iK�d���ι���{���!��2���=���A���=���2�%�!�y������﴾\�����2���ν�
"�p�&<��I=�=���=�`�=F@>^�>�   �   ��> �>4� >;v�=���=��=(��=<��=���=��p=�?=�R=4�<�H/< �&9����x��[���V��`��0�{�8tR� 6O�\���s�xJO�)���i��\,F�հ���˵�����	����Lx/��L:�O>�%U:�x/�B��\&	�&o�wL���)����.��ɽ8K��9<�2L=\J�=���=QM�=ek >�>�   �   [\>o��=p?�=���=���=���=ȹ�=U�=��w=�&I=�=�t�<���<��;� 3�����[n�\d���^��(�d� 7+��z� :໰�2�����v|.�mkh���6��6��[+��X�־���x����%���/��3��0�3�%�h��Xn�kpվͦ�gt���"�`M���:���m<�ZR=⺢=&��=h��=��=�>�   �   ���=)��=&w�=�+�=��=v��=���=��^=� 0=.�=\��<P�Q<`�; �-�g	��%K�0�k���g�0�@�@!�� �H� �W:�>;���� �6������t��TϽ�7���b����A�����y�=�����:#�- �#�������TU��3���G[�i������KƼ��<f�Z=̭�=Tw�=<��=8��=@,�=�   �   �'�=:��=�8�=���=K�=��b=�,+=�V�<�+�<���;�fʺ ��"X����\���~��X���x�F��aỀ���μ;�P3<�[<�^8<`r4;��c��$�������t^=����ѥ�2/ʾ������c�%�����'��ދ��̾:'���i��c'<�F���X��o�X��<�\b=�/�=��=@��=��=���=�   �   ��=�ү=�ޕ=|n=�~+=dp�<��<pg��ĵ���伨�����,���_��|�� ߼d���X�E� I����;�Ws<���<��<<H�<�,�<`��;�~����N�'�����eyN���T]��V�¾�پH��7�l���ܾ?Ǿ�`��]G�� `X�pX� �½P�=��w���8�<��f=3�=Jd�=^��=r��=چ�=�   �   ꜟ=�_�=R�C=�8�<Щ�; �`���	��rP����.����v��ֶ���m�����D_�@�,�����x� mɺ�;<,��< l=�w=h�!=��=���<�L�;����lOk�4�ͽ9��8�M�P���A��K���󉹾�ž��ӻ����ë��nV��**`�L�+�[���J������/�;n�=-e=��=oT�=ҭ�=]&�=9�=�   �   9i=fs =��<hA����{�rx��9;۽����|�\n�����6�ѽO׫��_����/��n��@�U���i<$4�<2*=�K=�/Z=�,R= �0=��< ��;�ʺ�HNm��fȽ|��t�:�2b��
�������ː�{(��U���kt��<R�o/+�oI��/��|�Q��`�� 8+<�=�"[=T%�=R�=��=b��=��=�   �   VL=V <�㕼��M�M���B���{�y�2�UE�tFN���M�&�C��a1�������>����F��j��8B��Oe<��=hrG=$8t=�r�=�̇=.�z=f�L=jT=�| <�̕��M��y�����w�x�2�@E�xAN�֞M��C��]1����9��ꤼ�lD��:��@��Le<�=�oG=�4t=�p�=4ʇ=��z=��L=�   �   X�;�ߺ�[m�nȽڳ�\�:��b��������zΐ�%+��lW��pt�@@R�2+�fK�d2����Q�$c��x8+<=�$[=�&�=�=��=㏞=��=4@i=�{ =��<������{�fp���2۽�����w�qj��{���O�ѽ�ӫ� ]����/��l��@�U���i<d/�<*=D�K=R+Z=f'R=�0=X��<�   �   `
���Zk�
�ͽF����M��R���D��S�������Ⱦ��ֻ�!������HX��-`�v�+�R��L��D��� ,�;,�=�.e=,��=�U�=���=�(�=�;�=���=-c�=��C=LL�<��;�R`�~�	�eP���m���6p��=����h������
_���,�0�� �x� �ɺ��;<x�<�h=�s=��!=�=���<0�;�   �   l�N��d ��}N���`��G�¾*�پi��F��bo�|�ܾ{
Ǿ�b���H��GbX��Y��½D�=�p|���9�<�f=4�=�e�=���=@��=��=l��=�կ=?�=�n=և+=��<h<@������������*��Z�y�,߼�����E�@,I�0��;PKs<��<���<�>�<�!�< [�;�����   �   -ƞ�T��a=����gӥ��1ʾ�"�W��Me����5��W����;�̾�(���j���(<���rZ�X o���<�]b=�0�=��=x��=:�=L��=�)�=���=�;�=��=�N�=Z�b=�4+=�f�< <�<��;��ɺ���`X��x�����T|��������F� q� ��@��;B3<@�Z<�K8<�4;��c��%��   �   �XϽ:���b�����C��=�-{�a>����<#�H �������UV��뛖�8[��i�L����KƼ�<|�Z=���=+x�=8��=\��=�-�=:��=��=,y�=�-�=0�=,��=i��=^�^=X0=��=��<��Q<P9�; �-��a	��$K�P�k���g�(�@�p5�� �H���V:�;�f���6�<����t��   �   �k��<�6��7���,���־{��l����%���/��3�`0���%����n��pվgͦ��t��"�KM��>:���m<�[R=���=���=4��=��=%>�\>� �=�@�=���=4��=ɂ�=���=4�=,�w=,*I=�=�y�<t��<���;��2�P���^n��f�� b��`�d��@+�Џ�Q�H�2�Ī��,�.�M��   �   ����-F������̵�	�侭�	�>���x/�=M:��>��U:�^x/�q��t&	�0o�hL���)��9�.��ɽ�I� �9<4L=K�=���=�M�=�k >n�>�>��>�� >w�=z��=��=��=)��=���=r�p=d�?=�S=���<J/< �&9p��xx��]��<Y��4��p�{�X{R�>O� ����x��MO�M����   �   ��jK������ι�{��U{���!�)�2���=���A���=���2��!�9��	��g﴾������2��νH"� �&<��I=��=��=:a�=z@>��>�8>̮>-�>Rb�=z%�=Z:�=�)�=�c�=�?�=z�}=�zK=ܮ=<��<(zG<@{�:�W	���|���������M��|,��poq� p�PJ���{ �n�Z�Ye���   �   ����,F�鰉��˵������	�r��x/�VL:��>��T:��w/�����%	�n�nK���(���.�ɽ�F��9<x5L=�K�=���=*N�=�k >}�>,�>��>�� >.w�=���=��=F��=a��=ꁐ=$�p=J�?=�T=,��<HP/< j(9h���x�8Y���T��d����{��qR�`4O����ls��JO������   �   �g����6�96���*����־#����ߛ%�+�/�2�3��0�<�%�v��om��nվ�˦��t���"��I��5�8�m<�^R=���=���=���=I��=I>]>� �=�@�=���=i��=��=���=��=2�w=z+I=��=�}�<p��<p��;`�2� �� Nn�,^���X��؋d��-+��j�p,�(�2�����l{.��혽�   �   SϽ�6���b�>���@����y�<�����9#�� �ߴ�x�y��<S��Z���[�Zf�o���L=Ƽ���<b�Z=鯢=.y�=���=ܖ�=�-�=���=+��=gy�=3.�=w�=���=ֈ�=x�^=�0=b�=���<P�Q< U�;��-��N	�@K��k�H�g��s@���� kH� �X:@k;����p�6�4���Vt��   �   J�����\=�����ϥ�b-ʾ�뾧��zb����e���������̾�$���g���#<�=���N�P�n�	�<�bb=G2�=&��=U��=��=���=F*�=؂�=�;�=T��=�N�=.�b=�5+=di�<t?�<�'�; ,ɺ�����W��n��X����o��������F��3� ����;(a3<�[<pl8<��4;��c�:�$��   �   N�N��{������vN�����J[����¾a�پT����Si���ܾ9Ǿ�]���D���[X��T���½�w=��/���G�<H�f=�5�=�f�=���=��=v��=΅�= ֯=��=��n=��+=���<�<P��x���@����T������T��r�X߼Р��P�E�@�H� �;�ms<4ò<� �<hP�<�4�< ��;�u���   �   X봼�Gk���ͽT����M��M��G?������􆹾s¾��л�e�������S��%`�ֽ+����ND��Xk���z�;x�=4e= Õ=NW�=���=8)�=$<�=X��=�c�=f�C=�M�< �;�O`�n�	��cP�# ��H����n��a����f��%���_���,����h�x� ~Ⱥ�<<� �<Bq=�|=��!=�=���<�u�;�   �   ���;x����Dm��`Ƚ��^�:�}b�.��󋾨Ȑ�p%��R��2ft�{7R��*+�$E�>(����Q�DJ��8^+<$=�)[=�(�=l�=��=���=`�=�@i=�| = �<P���{��o��"2۽-���Jw��i�{�i�ıѽ�Ы��Y��@�/��\�� (U�`	j<H@�<�*=��K=d4Z=,1R=�0=���<�   �   nZ=�� <@���^�M�"s�����r���2�
E�<N�S�M�z�C��X1����M��蜼�U=���z����re<@�=6wG=�;t=0t�=u͇=j�z=X�L=.U=@ <�˕�v�M�8y��3���v�4�2��E�AN�;�M�&�C��\1�������䡼�A�����!��ke<̇=�wG=�<t=/u�=�·=ʩz=��L=�   �   �Ei=n� =�(�<�� �n���t{��h��n*۽���s��e�>w�d
񽬫ѽ�˫��U����/�PU���U�Hj<�?�<h*=$�K=�1Z=*.R=<�0=̒�<p��;�ɺ��Mm�LfȽZ��M�:�b��
������wː�<(���T��"kt��;R�I.+� H��,��8�Q�XS��(S+<�=�)[=�(�=+�=�=��=:�=�   �   `��=f�=��C=�\�<�O�;@&`��y	�WP��������%h��8���a��h����^�Կ,�ȹ���x�@_Ⱥ�<<���<�o=Nz=8�!=��=���< R�;�����Nk���ͽ���M�	P���A��7���ى��sž��ӻ�N��r���
V��<)`�9�+����FH���v�� ]�;Z�=,3e=)Õ=�W�=l��=h*�=�=�=�   �   k��=,د=�=��n=��+=0��<`@<��������P��֢����8���M�`m�<߼ț��`�E� �H����;xgs<@��<4��<K�</�<`��;�}��t�N��~�����OyN�z�J]��K�¾�پ7����el꾹�ܾǾg`��G��J_X�~W��½�}=��R��LB�<��f=�5�=g�=]��=ҭ�=���=�   �   �+�=i��=�=�=���=�Q�=z�b=�<+=px�<O�<�f�;�:Ⱥ0����W��d���Lj��������F��7� ����;pY3<�[<c8< 4;@�c���$�i���t�b^=����ѥ�+/ʾ������c�����������Z�̾�&��_i���&<����hU��o���<�`b=�1�=��=���=l�=���=�   �   ]��=?��=�z�=�/�=r�=���=T��=��^=F0=�=Dô<��Q<w�;`L-��D	��K� �k�(�g�Hv@�P
����H��X:�O;�Ǖ���6�(����t�rTϽ�7���b����A�����y�=�����:#�' ��������*U�������[�xh������FƼ\�<>�Z=H��=�x�=���=$��=�.�=�   �   8]>t�=�A�=���=���=r��=���=I�=��w=/I="�=���<쿂<0��;�2����Ln�(^���Y�� �d��1+��r�04໸�2�,���2|.�URh���6��6��W+��U�־���v����%���/��3��0�-�%�a��Nn�Qpվ�̦�t���"��L��D9���m<Z\R=ڻ�=,��=���=R��=g>�   �   6�>��>ˍ >�w�=��=��=���=,��=���=��p=�?=JV=4��<@U/< ^)9h��x��X��xT�������{�XrR�p4O������r�RJO����c��Y,F�Ӱ���˵�����	����Lx/��L:�O>�"U:�x/�@��W&	�o�jL���)��l�.�HɽdJ�X�9<v3L=�J�=y��=�M�=�k >y�>�   �   n>�G >�Q�=�=�,�=)��=\)�=eѣ=S�=�k�=p�c=$G=^y-=(F=�'=\q�<t��< �<d��<@L�<�v�<��<�V:<�����L��d��hm�v�R�%ę�nӾ6
���+��M�m�j������z������z���Pj�qL�y�*�,<�"�;t{��j�:�<ʽ�4�$ģ<z2q=�W�=<�=L?�=�> >�   �   �` >�$�=���=f��=���=V\�=�G�=�t�=k��=��o=֡Q=�}6=��=�
=h��<lu�<���<���<���<l�<�o�<hU�<�bS< m�t$��2%��zY��9M�uI����ξ�F�,�(�!6I��Jf�O}�,��������N}��f�m�H�B�'�9��g�ɾY_���o6�U�ý8���i�<0xs=ns�=OQ�=:��=P��=�   �   88�=:��=���=j�=Z��=�w�=,5�=�{=$�V=�5=�=U=�Z�<8$�<��<(��<���<�
�<���<D��<���<��<x��<@q�:Ђ��b�{�u 뽚�=��1��"¾(������>���Y���o���}��v�� ~��p���Y��=����*��Sڽ��b��n)�K屽_ż���<��y=7��=H��=RX�=��=�   �   �Q�=`�=���=�z�=H��=��y=t@G=0=F�<�&�<�e<0:(<0^
<��<�V <@�L<�<�}�<���<T8�<�� =T&�<�O�<�`*< �O���B���ŽMs%���x�`��9�� +���,��pF���Z���g��l��/h�x9[�K�F�"-�;-�����h��D�n�x]�M���N|����<�,�= �=���=
2�=j��=�   �   V��=�v�=q��=�= ?=؉�<�{<��:P�����%���⵼䋧��愼@�$�`!&��&�;@�m<���<�,�<Z=	=��=h�<���:p���ˬ��&��,Q�F����Mƾ1�����]�-�~@�L�K�#P��BL���@�&�.�2���"���%Ǿ�>��X(L�����>4h�`?��T=���=v��=`��=���=�)�=�   �   �;�=2<�=�Q=�;=�K-<X)�|~���=���p��L���֍�8d��D&x�B<O��%��Ƽ���_�;��<���<~�=��+=�y'=`=1�<h���B�*�ǽ�$��@p��ᢾ��Ͼ�!��K��I�!�},���/���,�y�"�/v�f���L�Ӿ�(��<�t���%�4������ S�;�J)=N��=��=��=��=���=�   �   &z=�+=��<���Dx�����N���߽I����*�����T�v��#lŽ�Z�� \��� �`&�@�<p�<XD=&�?=d�I=t58=�=��:<���+}�j3���4��T|�$У�(�Ⱦ��1a�l�l�������^���Fξu��p���@�iQ��>R���ܧ�hX�<H�==��=��=�ҭ=nj�=�ř=�   �   ��= <�]��&�d�］_-���$���?���R�R�[�� Z�6<N�	�9��������Ǽ��w�t��� �i���<b	=�L=�g=&f=��E=J�=�E�; ۼ�B�������4�xr����]��'�Ǿ^U־�ܾs�ؾ�0̾�P���۞�^���H�.�$��h.� ?�����<��K=��=��=$�=Ņ�=r"c=�   �   0��;<������U�Rj#�E�R���}��A������~����֞�P敾�#��h���<��.���Žz9g� 0��HH<�=BQ=\�}=t �=|�=N�R=V�=p%�;8#�^���yL�e#�A�R��}�$>��Q�������1Ӟ�9㕾!��vh��<�,���Ž�3g�x)��0N<�=�Q=��}=���=��=�R=X�=�   �   8ۼ�I��#���7�4�sr������ǾhY־�ܾ?�ؾh4̾T��ޞ�t��=�H���\��d.�`O�����<~�K=��=��=&&�=���=n)c=N�=(I <�C����d��弽J(��$���?���R�V�[�:�Y�7N�u�9�Ĥ�����K¼�2 w������ri�t�<�=R�L=*g=�!f=~�E=`�= ��;�   �   �6}��:�l�4�\Z|�aӣ���Ⱦ��Oc��!�9n���������Iξ�奄�r����@��T��hT��h᧼�V�<��==��=��=�ԭ=�l�=�ș=�#z=�+=��< ���ji��؀��D��+߽|���&����P����eŽ�U���\��� ��&�(�<(p�<.C=�?=�I=�08=2 =�:<����   �   C�ǽh$��Ep�j䢾+�Ͼ]%��T��l�!��,���/���,�L�"��w����r�Ӿ+*���u�>�%�O����� L�;.K)=팈=��=J�=ظ�=/��=�>�=�?�=��Q=�E= {-<��(��a��r=���p�E���ύ��]���x��2O�~�� Ƽhs�p�;@�<���<��=�+= v'=�=@%�<���LB��   �   ���Q������Pƾa������L�-��@�S�K�P��DL�y�@���.�e���$��1'Ǿ�?���)L�����6h��D���=��=\��=���=��=�+�=���=�y�=���=�=
?=��<h�{<�> ;p`��ꇼ����ϵ�@{��8ل� �$���%� :�;��m<���<�*�<|=Z=�=Pج<@	�:���{����   �   v%�A�x�u�����m,�;�,�frF�y�Z�y�g���l�l1h��:[�p�F�#-��-���侹i��8�n�^��M��O|���<E-�=��=���=E3�=��=cS�=��=���=�}�=���=�y=0HG=B=PV�<�6�<x�e<�T(<u
<p	<e <��L<��<�~�<$��<6�<�� =D!�<I�<�O*< �O�jC���Ž�   �   �=�X3���#¾/������>��Y���o���}��w��,!~��p�R�Y���=�o��`+���ڽ�&c��,n)� 屽�]ż��<�y=숲=��=CY�=��=�9�=���=B��=�k�=���=5z�=�7�=8�{=V�V=�5=R=$Y=�a�<�)�<���<���<���<p
�<X��<���<\��<�<䓍< ��:ȋ���{���   �   9;M��J����ξ�G���(��6I��Kf��O}����]���6��sN}��f���H�J�'�1��>�ɾ"_��.o6�i�ý����l�<�ys=#t�=�Q�=��=��=?a >�%�=���=���= ��=�]�="I�=v�=���=4�o=�Q=�6=d�=. =���<�u�<���<���<<��<H�<�l�<R�<hZS<`:m�@+��]'���Z��   �   ��R��ę��nӾ�
�!�+�SM���j������z������z����Oj��pL��*��;�q�;�z��\�:��ʽ2��ȣ<B4q=LX�=��=�?�=? >�> H > R�=X�=�,�=Z��=�)�=�ѣ=`�=�k�=J�c=�#G=�x-=�E=B'=$p�<@��<��<��<�J�<�t�<�}�<pQ:<�����N�9f��Jn��   �   �9M��I����ξ�F�"�(��5I��Jf��N}�����������KM}��f���H�{�'����*�ɾL^���m6���ýd���p�<{s=�t�=TR�=$��=2��=Oa >�%�=���=���=2��=�]�=8I�=<v�=⋈=��o=��Q=8�6=D�=8=0��<�x�<��<���<���<��<Lp�<�U�<�bS<@m��%���%���Y��   �   F�=��1���!¾����a�>� �Y���o���}�_v���~�rp�K�Y���=��~��(���ؽ��a���k)��ᱽ`Sż`��<��y=׉�=ų�=�Y�=�=�9�=���=i��= l�=���=az�=�7�=��{=�V=��5=t=�Z=e�<�-�<���<���<L��<x�<���<`��<(��<8�<���<���:x�����{�	 ��   �   br%���x�����;*���,��oF�b�Z�;�g�C�l�2.h��7[���F�� -��+����f����n��Z��H���2|�D��</�=�=���=�3�=Y��=�S�=��=���=
~�=ɚ�=f�y=�HG=�=,X�<�8�<��e<`\(<H~
<X	<�q < �L<|�<І�<��<?�<�� =8+�<�S�<Ph*<X�O���B�4�Ž�   �   Ţ�WQ����,Lƾ*��������-��@�t�K�/P��@L���@�<�.�j������"Ǿy<���$L�ħ��V*h������#=G��=俯=���=ք�=6,�=��=�y�=��=��=�
?=��<��{<�K ;0\��燼 ��,˵��u���҄���$���%�P_�;�n<��<�5�<0=d=��=0�<@ �:���������   �   Єǽd�#�>p��ߢ���Ͼ������p�!�y,���/�w�,�U�"�%t������Ӿ�%��W�t���%���������;�Q)=]��=t�=~�=���=���=?�=7@�=n�Q=�F=8}-<X�(��`�r=�^�p�GD���΍��\��x�J/O�h���ż�^�P��;�*�<��<(�=��+=@}'=�=�8�<P���B��   �   �#}��.���4��P|��ͣ�F�Ⱦ5�P_�a��i�W�����Q��-Cξ#ꩾ�m��5�@�bI���K��@ǧ�j�<��==�=��=�խ=�m�= ə=n$z=��+=��<����h�E؀��D���
߽�����%�����O����4dŽ�S��	\�t� ���%���<p|�<�I=Ĺ?=��I=v98=&
=�;<H����   �   �ڼ>������O�4�� r�� ��'����ǾzQ־�
ܾV�ؾ�,̾&M��؞�=����H����p���.��ꉻ8��<H�K=`�=<�=X'�=Z��=�*c="�=�K <|B��"�d��弽&(���$���?�U�R��[���Y�u6N�Ƽ9����������B�v�(����i�X��<�=��L=v�g=:*f=B�E=8�=�t�;�   �   �^�;L⼻���uE��`#�4�R�D�}��:����J�Ϟ��ߕ����&h�i�<�.'��Ž�%g�t���v<��=�Q=��}=�=��=��R=f�=�+�; "����?L��d#�%�R���}�>��7�������Ӟ��╾� ���h�0�<�!+�P�Ž/g�8���c< =$Q=��}=��=��=$�R=�=�   �   ��=hi <x/��F{d��޼��#��$�'�?���R��[���Y��0N���9�N����������v�������h�T��<�=��L=�g=�(f=��E=��= M�;�ۼ�B��i��� �4�^r����Q���ǾIU־�ܾN�ؾ�0̾�P��5۞� ��-�H�<����.����Ĥ�<.�K=	�=|�=-(�=Ɋ�=�.c=�   �   :)z=�+=�*�<@H���\�;р��<���߽����� ����^K�G���\ŽxM����[�|� ��%���<\��<�J=ҹ?=��I=�78=�=��:<8��x*}�23꽺�4��T|�У��Ⱦ��,a�f�l�x�����0�Fξ-�~p��E�@��O��VP���ԧ�$a�< �==~�=��=u֭=�n�=�ʙ=�   �   �@�=�B�=��Q=�N=��-<��(�XG�Ld=���p��<��|Ǎ��U��"x��#O�����żXG����;T0�<��<��=r�+=B|'=4=�3�<���B���ǽ~$��@p��ᢾ��Ͼ�!��I��F�!�x,���/���,�m�"�v�:����ӾB(����t��%�����X��o�;�N)=|��=2�=��=x��=��=�   �   ���=�{�=���=��=�?=��<(|<�� ;80�hч�����L����b�� �إ$��F%�0��;�n<Ď�<�7�<Z=�=��=0�<�ߎ:,���������Q�=����Mƾ,�����\�-�}@�K�K� P��BL���@��.�#���"���%Ǿ�>���'L�Ҭ���1h�`)��R =?��=n��=���=Y��=--�=�   �   �T�="�=~��=2��=e��=t�y=�OG=R=�g�<�H�<��e<�y(<0�
<�-	<@� <��L<T��<���<H��<0@�<�� =�*�<�R�<�d*<H�O�B�B�b�Ž:s%���x�Z��4���*���,��pF���Z���g��l��/h�t9[�E�F�"-�/-�k���h����n�]�:L���F|�L��<�-�=k�=f��=4�=��=�   �   B:�=���=v��=wm�=O��=F|�=:�=`�{=��V= �5=j=>_=�m�<X5�<���<��<<¹<0�<H��<D��<X��<,�<\��< ��:����{�U 뽏�=��1��"¾%������>���Y���o���}��v�� ~��p���Y��=����*��<ڽ��b���m)��䱽�\ż���<P�y="��=l��=�Y�=>�=�   �   Xa >>&�=:��= ��=���=�^�=0J�=Rw�=��=�o=�Q=��6=��=@=��<�{�<��<� �<���<��<Hq�<�V�<�dS<`	m��#��%��sY�|9M�rI����ξ�F�+�(�!6I��Jf�O}�-��������N}��f�j�H�>�'�6��[�ɾL_���o6��ý���k�<�xs=�s�=�Q�=���=$��=�   �   �[�=��=,�=���=m*�=�x�=v%�=�K�=|�="h=�V=��J=��D=�C=ҋF=��L=��T=X*\=4`=Z�[=ިH=�:=�K�<p�����N���㽭F�:Ù�}�ݾ�z�aB�@�o�ݍ��I��2����f���ʽ��f�����~��~�����n�ع@��0�LL׾�u���=0����P��HU
=��=]r�=v��=��=�   �   �,�=ل�=`U�=���=Dκ=X�=���=x��=T�e=zoN=�==r3=�}/=j1=��6=�5@=�*K=�U=�=\= 7Z=�vI=p4"=D��<�Q���>D�Y5ܽ�@��I����ؾ���s�>���k��Y���{��5���g:��Γ��q@������^��
����j��8=�,d�ӾwO���+�ؔ���l�ZQ=C�=�Ϳ=~��=���=�   �   �u�=r�=S��=>R�=qS�=���=�o`=�v8=��=���<��<���<���<X<�<�7=��=�".=|fA=FP=OU=�CK=g*= #�< ���%��ƽ�2��5��'�˾	�
�� 4�(�^����
T�����!���;��h��ۤ�X`���򃿮>^�
3��B	�2�ƾi.��D���n���T���=P��=P��=�+�=X��=�   �   ���=��=6�==q�=v�Z=��=���<��W<�r�;`��������� �5����;5O<(��<<��<>7=��9=�K=P*L=��5=��<@L�;�8鼂٤���� y��Ŷ�E?����#��K��:q�K���b������V����6��]ԉ�	�q�xK��#�&��F-��y�m��2�s�@ǡ�vS*=�T�=:p�=J�=��=�   �   ��=Zl�=">i=Fh=�>�<�(^��%����
��?8�nZR��X�>TJ��J+��*��P�� EY��7<���<ι=N�8=VJI=�ZA=��=���<�Q]���s�h���d3Q��s��oپϔ���1�TT�ĕr�aW�� ���䏿�^��&ą�D�s�U�z�2����0پԱ��/J���
-1���<��==�%�=&M�=�p�=�R�=�   �   ���="�>=�J�< 첺 �漌�_�r
gɽ-��U����5彬�ɽq(��vPt�n��P�v����;$�<
�=�t?=��I=tB4=̟�<�(T;� �uc���Y$��}�^��"��ko�F%3�1�M�Ѳb��Sp��?u�~�p���c�`O��4�4���0�������~�A"�TW��(�ϼ���<�+P=��=�_�=(�=���=�   �   ��=�GX< i��TV��t��hX���) �1�:�#RM��U�ZCS���F�.�1���+l��D��@�L��I����;pk�<`�+=�XL=H�K=zN%=8I�<�1:��<f� t�`<@��싾���6��Q��C '�]�8��vD�e�H��6E�0L:��)����OS������ߏ��rF���Sg� _����<��^=���=�=�=o=�   �   p��;O��[�����l�'��(X�3��O���ʖ��j���������@���j��s=��j��Z���pZ�H.��8�C<��=�F=�E]=��N=z�=x�M<�O��vS���j�~<K�����X��Q�޾ڍ���w��5*�Ox�|��n��p�侧ϼ��Ɠ���X����p����}����<��=d�f=(!�=�T�=4G]=�q=�   �   ����;��{���B������|��s��վsI侣:��c�5پ�ľ먾	N��gHU���i^���@>�������<ڰ5=��f=�p=:`S=�=�Q�;����3������B�����x����Vվ�D��5�)_��0پ�ľ�稾bK��8DU����Y���:>�������<��5=��f=��p=�ZS=��=��;�   �   �Z���n�BK��
���\����޾[����0���,��z��������供Ҽ�ɓ�/�X������������<P�=��f=�"�=�V�=�M]=z=p��;�3�kS����r�'��!X�t��R�������S~��*�������<����j�Go=��f�qU��<iZ�|$��0 D<��=�F=�C]=v�N=��=�hM<4e���   �   �{�?A@��ʹ���������"'�2�8��yD�>�H�c9E��N:��)����cV��] ���᏾@uF����Xg��p����<��^=���= �=��=o=��=uX<M��^CV� k��_M���# ���:�{KM�e�U�=S���F���1�����d�=?����L��=�� �;o�<��+=8WL=h�K=�I%=P<�<�T:�vHf��   �   �]$�!�}�?a�����q��'3��M���b��Vp��Bu�+�p� �c��O���4����53�����~��B"�VY��d�ϼ���<�,P=��=/a�=V�=���=S��=T�>=0a�< C��`��<v_��堽�\ɽ����J��5��"彤�ɽ�!��,Et����H�v� ɹ;d�<�=ft?=�I=6?4=(��<�S;�)�yi���   �   <7Q�sv�� rپ����1�� T�R�r��X��u ��揿�_��?Ņ�0�s��	U�Ȏ2�����پ߲��x0J�佬.1�@�<n�==�&�=nN�=�r�=EU�=΂�=�o�=�Fi=|r= V�< �Z������
�p08�.KR��X��FJ��>+�,���񐼠�X�س7<ȴ�<z�=��8=pII=�XA=@�=��<Pl]���s�R����   �   �y��Ƕ�B��U�#��K��<q�g������������V����7�� Չ�I�q�t	K��#�-'���-��W�m����s�����hT*=bU�=Jq�=K�=� �=���=4�=h�=�t�=��Z=�=���<P�W<�ɂ; ��l���X�� �3�P�;�KO<���<l��<(9=ȅ9=�K=()L=��5=��<�'�;�D鼟ݤ�����   �   7���˾1�
�B"4���^�U���T���������f<�����ۤ��`����=?^�f
3�2C	�u�ƾ�.��@��En��Q�ʝ=��=6��=�,�=���=�w�=R�=x��=�T�=AV�=½�=�v`=�}8=��=\��<���<���< ��<E�<B;=0�=>$.=^gA=vP=|NU=�BK=e*=4�<���%%��ƽ�2��   �   �J���ؾl��h�>���k�/Z��|�������:��6����@������;^��!����j��8=�d��Ӿ-O����+�ѓ��P�l�S=�=zο=N��={��=�-�=��=�V�=��=�Ϻ=��=`��=6��=��e=�rN=�==�t3=�/=@1=� 7=�6@=�*K=�U=D=\=^6Z=vuI=�2"=���< k��
CD�8ܽ��@��   �   �Ù�U�ݾs{��aB���o�Vݍ��I��V����f���ʽ��f��∰�M��D�����n�Z�@�|0�wK׾�t���<0��}������W
=ノ=s�=��=���=h\�=|��=��=��=�*�=>y�=�%�=L�=��=&h=�V=F�J=8�D=x�C=<�F=ڧL=>�T=�)\=X`=f�[=��H=�9=(H�<������N�w���F��   �   J����ؾ���z�>���k��Y��]{������:��h����?�� ����]������j�8=�Zc�� ӾVN��R�+������l��T=��=�ο=���=���=�-�=
��=�V�=��=�Ϻ=�=r��=K��=�e=sN=t�==,u3=��/=�1=�7=`7@=�+K=�U=j>\=�7Z=�vI=P4"=@��<�X��@D�"6ܽ��@��   �   b5��ӏ˾��
�~ 4���^����S������o ���:�����Dڤ��_����0=^��3��A	�S�ƾ�,������j��X>��=5��=���=<-�=��=�w�={�=���=�T�=aV�=ݽ�=�v`=�}8=:�=h��<,��<x��<L��<�G�<�<=��=(&.=jiA=�	P=�PU=*EK=h*=h$�<���b%�D�ƽr2��   �   ��x��Ķ�>���#��
K��9q�������򍟿w���:����5��GӉ���q��K�>#�^#��+����m�V���s���X*=�V�=ar�=:L�=:!�=$��=q�=��=u�=D�Z=r�=���<�W<�΂;���Pd���N���U3����;XTO<���<���< <=�9="K=�,L=��5=��<�Y�;5�hؤ����   �   �1Q��r��umپ�����1��T�דr�HV������㏿8]������s��U�_�2���"پ\���0+J�\�~#1���<��==�(�=�O�=fs�=�U�=:��=9p�=>Gi=�r=�V�< �Z�$��:�
��/8�PJR��X�\EJ��<+�����쐼 �X�@�7<���<(�=��8=�MI=�]A=P�=< F]��s������   �   �W$�E�}�8\������m�k#3��M�b�b�FQp�=u���p���c��O�m�4����-�����x�~��<"��P���ϼ�<�2P=�=�b�=O�=E��=���=��>=,b�<@5������u_��堽�\ɽ���`J�����`影�ɽh ��|Bt������v���;��<|�=Ry?=��I=�E4=���<�eT;��d`���   �   �o�X9@��ꋾ������f��	'���8��sD���H��3E�]I:�� )�S���N��5���܏��mF�����Fg�0��h$�<��^=�=��=��=r	o=��=�wX<L���BV��j��,M���# ���:�RKM�/�U��<S���F���1����c뽱=��4�L�p6��P.�;(x�<��+=]L=L�K=tR%=�Q�<�:��5f��   �   �N��zg��8K����U����޾���~����'��u�������Ԑ侔˼�3Ó�߃X�Ь��� e���<�=��f=�$�=LX�=xO]=T{=���;L2�)S��L��[�'��!X�i��D�������<~��
��Ө���<���j��n=�@f��S���eZ�����D<��=tF=DJ]=��N=�=x�M<�A���   �   L��.����S�B�=����u��%��վ�?��0�AZ�,پU ľ�㨾�G���=U�~�EQ���,>�P[���<ظ5=D�f=�p=�bS=��=0[�;��z3��h��ՏB�����x�����Mվ�D便5�_澰0پ�ľ�稾K���CU��NX��7>���� ��<µ5=��f=F�p=�dS=x�=���;�   �   p#�;p��L��|�뽐�'�2X�!�����������/z�����ꤘ��8����j�i=��a�EL���YZ���0*D<��=� F=�J]=��N=��=��M<tM��S��^j�d<K�z���X��J�޾׍���t��/*�Ex�n��\��C��nϼ�nƓ��X�ް������v����<(= �f=�$�=�X�=�R]=.�=�   �   z�=��X<\7���5V�c���C��S ���:��DM���U�26S�M�F���1�إ��Z�06��"�L��#��pe�;ԁ�<��+=�^L=��K=`Q%=$M�<�,:��;f��s�D<@��싾���/��O��A '�[�8��vD�a�H��6E�(L:��)����$S������ߏ�rF�����Pg�@D��|�<v�^=���=��= �=�o=�   �   !Ą=j�>=�r�< ꯺���g_�^ݠ�vSɽ���/@��{��彬�ɽV���4t���X�v�p �;(�<�=�{?=��I=�E4=h��< AT;��c���Y$��}�^����io�D%3�0�M�Ҳb��Sp��?u�|�p���c�XO�۫4�$���0�����(�~�}@"�$V����ϼ��<�/P=j�=�b�=(�=ԧ�=�   �   ���=�r�=�Mi=�z=�i�< �W��R�
�!8�&;R���W��6J�r/+������א��%X��7<8��<�=V�8=�OI=L^A=2�=D��<@M]���s�*���M3Q��s��
oپ̔���1�ST�ƕr�bW��!���䏿�^��$ą�A�s�U�o�2����پ�����.J����*1���<̡==�'�=�O�=�s�=�V�=�   �   P��=!�=��=�w�=[=R�=l��<(�W<p!�; A����`��� �0��A�;�qO<���<��<�?=��9=K=.L=��5=��<pV�;�6�?٤���� y��Ŷ�A?����#��K��:q�K���b���������W����6��]ԉ��q�rK��#�&��(-��6�m�����s� ����U*=V�=r�=bL�=�!�=�   �   nx�=z�=���=�V�=yX�=U��=l|`=�8=��=� =���<x��<���<�R�<�A=�=�).=
lA=�P=PRU=*FK=�h*=T%�<���6%�S�ƽ�2��5��#�˾�
�� 4�'�^����T�����!���;��i��ۤ�X`��~򃿪>^� 
3��B	� �ƾT.����n��8P���=9��=|��=-�=I��=�   �   �-�=V��=&W�=���=�к=�=���=���=$f=XvN=ȧ==|x3=��/=�1=R7=�9@=�-K=��U=�?\=�8Z=�wI=N5"=d��<@N���>D�D5ܽ�@��I����ؾ���s�>���k��Y���{��6���i:��Г��r@������^��
����j��8=�)d�ӾkO����+�������l�R=��=Aο=>��=���=�   �   /��=*F�=�h�=d��=�a�=���=�=�N`=�F=�4=�s,=dA-=6=R�E=plY=ro=�b�=�ʊ=`}�=�q�=�u=!6=�Δ<�n���զ�
�'�Ќ��־���!�K��`��6v��O����ӿ�X����[3������B翔�ӿͺ�����hg���I�6$��pϾ�݄�S��,[q��:�;��H=E=�=�f�=��=�   �   ��=��=p!�=㭳=7��=iW�=��d=��@=�j%=��=|/=|�==��,=��C=��]=�v=,��=�=__�=�t=��7=0I�<���� ����_#� �����Ѿ?�� +H��	�����`���Zп�{�t�￢�����Nw㿖-п���$	���Q~�2�E�T��D˾Q遾P��8-g�pK�;�K=��=�]�=n��=�   �   �;�=T��=,��==L�=Mt=,�==�L=P��<��<��9<�t$<�B<lv�<�ѿ<�9=jU'=�K=ʽj=Bw=:܁=�5p=4<=|�<H}o�tg�����'��T�ľQS�=��{r������خ��ƿFؿv�*�F,�toؿZƿx����<��>q��l;�2&
��%��c�r�,(�z�I�p3<P�P=�؟=4�=���=�   �   ��=B7�=��=NFB=�}�<�XG< n}�p^��4*ڼz�����+������@T;�ɑ<`� =�Z2=42X=�l=N&g=fA=� �<`����yd��s���b�Ui��������+�t8]������S��!ӵ�<�ƿ��ѿտ��ѿ�&ǿv/��ˈ��C���>�\���*����;:����W�5)��+�P؀<LBX=t��=P��=�x�=�   �   m8�=b�Z=�=(
(<�h��\�hyu����pQ��cĽ�½����h#��ƍk�����������;H�<f=�HG=0�V=�C=�a=�a�;޿���ν��=�-ۖ���۾y���(B��o�ˍ�h.���w���U���ܽ������
���ѡ�zX��2zp�WnB���
9ھ5B��6�����`�Ƽ<��<��^=��=�7�=���=�   �   ��4=hժ<p���|�#�;H���>۽N�d#%���5��J=���:�,l.����;���Ao���h���C��t�<�=�;=	A=��=d9�<�J��O���,��Dt�6Y�������#�#*K�lq�ӭ��>�������⢿�(�� ˗�����s��L��$���������&�r���م�(#�4��<��a=��=�ь=�x=�   �   �GL<d ����w�^�ֽ^�ƽI���s��܊��)���Ú��I�����K��IY� T-�+`���尿0�,�D����<�=b�5=,�,=��< �\9��.�0�ѽ��8������iǾ<��h�$��>E���a��x�ʃ�~���:���`z��d��lG��'�����aʾdԏ�0,;��ҽ�]$��u�;��=�V^=�s=��[=K=�   �   p�׼�N��� ��'>�Lp~����H����ѾX�ྺ����+�վ����}������S�N��������G-��!��l��<^�=��5=�K=2�<�h��"|��#���kN�����8kɾ�e������1��@D�uP�j�T��]Q�z�E���3�����a�՛ξ党��V�`��)`��d_���ʞ<2�*=R=��G=�M=0�<�   �   �������qP�1����캾NI�}��G���K��� �,;�p[��5��A��w��+_����]��W�����<���H�;���<�\5=r�;=��=@.D<��¼�����\kP�M���'躾D侚��3���H��� �%8��X�@3�==�^t��S\��V�]��T��~������_�;���<4[5=��;=��=�D<��¼�   �   �,��KqN�1ĕ��oɾ�j�����1�DD��xP���T��`Q���E���3���xc���ξG���m�V����8c��f���Ȟ<0�*=R=�G=<U=��<��׼�E���� �!>��h~�����f
����Ѿ���]�����b�վ>���́������w�N�8�N���F@-�@������<H�=��5=�G=h$�<�+h�^0|��   �   `�8�ⱍ�smǾ���6�$��AE�6b���x��˃����S<��dz�f
d�oG��'�A��dʾ-֏��.;��ҽ�a$��j�; �=,Y^=,�s=��[=�S=�tL<���4�w���ֽ���I���s��؊�`%��e����E���
�����CY�,O-�=X��y馽h�,�P,�dȒ<4=��5=r�,=��<  U9@/�yҽ�   �   �It�w\�����f�#��,K�Aoq�������s��䢿�*���̗�i���# s���L���$�H���I���t�r���څ��(����<��a=a�=Ԍ=�x=��4= �<�a����#�m>���3۽�G��%���5�D=���:�'f.�m���~���g��Ă�����`��`#�<@=��;=�A=V�=�.�<lZ������0��   �   �ݖ�Ԯ۾t��+B���o��̍�0���y��jW��]޽�6���V��&ӡ��Y���{p��oB���q:ھ%C��C6�ᙸ�<�Ƽ��<��^=��=�9�=t��=�;�=2�Z=Ɩ==(<H�g�L�gu���jG��)YĽm�½	���g���k�<�|ㅼP7�;�<�=LJG=
�V=L�C=v^=�6�;���0�νF�=��   �   �k��������+��:]������T���Ե���ƿb�ѿ#�տ��ѿ	(ǿm0����������6�\�8�*�޷���:����W��)�,��ـ<�CX=���=���=�z�=_�=�:�=��=�OB=,��<��G<`�|�C��$ڼ�����������0t� �;4֑<$� =^2="4X=Vl=�%g=nA=���<�辻��d�(v�c��   �   F�ľ�T�� =��}r�򟔿�ٮ��ƿ3Gؿ��+�)-�6pؿ�ƿ����;=���>q��l;�`&
��%��o�r�(���I��8<��P=�ٟ=q�=0��=�=�=���=���=LO�=
Tt=��==>U=ص�<���<�:<H�$<H�B<L��<�ݿ<�>=4Y'=̢K=��j= x=3܁=�4p=2<=4�<��o��j���M)���   �   �Ѿ*��5,H�~
��������P[п8|���'��C�￞w��-п3���,	���Q~��E��S�*D˾�聾����*g��[�;� K=��=�^�=p��=5��=h��=�"�=���=��=mY�=:�d=`�@=fo%=�=|3=�=:=4�,=��C= �]= �v=g��=��=_�=�~t=��7=�C�<���������a#�I����   �   �־e����K��`���v��dO��!�ӿ�X���]3�����B�W�ӿ�̺�����g��r�I��#��oϾ"݄�-���Wq�Q�; �H=>�=<g�=!�=���=�F�=,i�=ɨ�=Xb�=F��=V�=�N`=8F=&�4=�s,=A-=�6=ĄE=�kY=Jqo=ub�=�ʊ=�|�=q�=~�u=j6=Dʔ<pt���צ�:�'��Ќ��   �   �Ѿi��?+H��	�� ���C��jZп>{�
����@�￩v��,пj������P~�&�E�'S�C˾0聾����'g��l�;&"K=���=�^�=���=]��=���=#�=���=#��=yY�=X�d=��@=�o%=4�=�3=d�=�=��,=^�C=��]=��v=ƈ�=o�=�_�=�t=.�7=�G�<���� ���b`#�r����   �   �ľS��=�\{r�����خ�ƿZEؿ�
�)�;+�cnؿKƿt����;��l<q�!k;��$
��#��o�r��%���I�I<��P=�ڟ=�=���= >�=Ē�=���=fO�=6Tt=�==vU=4��<t��< :<�$<��B<���<<߿<�?=^Z'=�K=�j=�y=#݁= 7p=
<=��<�|o�bg�����'���   �   �h������!�+�r7]������R��(ҵ��ƿ��ѿj�տ8�ѿ~%ǿ.��������*�\���*�����7��b�W��#��#�D�<�GX=���=���=8{�=��=�:�=��=�OB=���<؈G< �|�|B��xڼ�� ������ho� �;hّ< � =`2=j6X=�!l=�(g=fA=��< ����wd��r���b��   �   ږ�!�۾o��V'B�)�o�ʍ�--���v��2T��۽� ���H	��VС��V���wp��kB����5ھ�?��H�5�ʒ��X�Ƽ䴻<0�^=��=;�=$��=f<�=��Z=4�=x>(<0�g��K��fu����?G���XĽ�½��������~k��}��߅��H�; �<L=xMG=ڟV=
�C=�d=�w�;�����ν�=��   �   TBt�fW������]�#�+(K��iq�r������񾟿ᢿ'��8ɗ�S����s�4�L���$�����V����r���	Ӆ���� ��<�a=!�=DՌ=Nx=��4=x�<�]��X�#�I>���3۽�G��%���5��C=�T�:��e.���.~���f���������P���t)�<�=Ԉ;=�A=�=�@�<DB�������*��   �   ��8�Ь���fǾ���Y�$�><E���a���x�Rȃ�<|���8��;]z�d�yiG�$	'�=���]ʾ4я�,';��ҽ�Q$��þ;�=�^^=��s=0�[=(U=�xL<�����w���ֽ
���I���s��؊�U%��W����E���
������BY��N-�5W��H覽��,� ��ϒ<~=
�5=Z�,=p��< Za9n�.��ѽ�   �   8���gN�����gɾ�a������1��=D��qP���T�ZQ�
�E���3�����^�[�ξ2����V�����X���G��$ޞ<��*=DR=��G=�W=�<��׼�E���� �� >�}h~�����a
����Ѿ���Q�����H�վ�������r�����N������X=-��᣻԰�<~�=~�5=�P=`<�<��g��|��   �   ����_���fP�X����亾�?���h���E��� ��4��U�V0��7꾴o��YX����]�JO�v��$�� ��;|��<�c5=8�;=�=�6D<4�¼����̵�BkP�E���!躾D侘��1���H��� �8��X�23�=�3t��\��ս]�T�T}������}�;D��<za5=�;=�=PGD<��¼�   �   0�׼�?���� ��>�Bb~������Ѿ������w���վI���L}��������N������:1-�����켶<,�=�5=&P=�7�<0�g��!|��#��hkN�����0kɾ�e������1��@D�uP�f�T��]Q�r�E���3����na���ξ����z�V�����^���X��0Ӟ<��*=�R=��G=[=x<�   �   ��L<���w�1�ֽ��|�I���s��Ԋ�*!�����eA���������;Y��H-�M��ঽʁ,���
��ݒ<J=��5=d�,=��< �^9&�.���ѽb�8�����yiǾ9��g�$��>E���a��x�ʃ�~���:���`z��d��lG��'����waʾ3ԏ��+;��ҽ*[$�0��;N�=]^=r�s=��[=�Y=�   �   ��4=l��<�	��2�#�@6��0*۽lB��%�K�5�L==���:�{_.� ��es��D]���y���u� ����8�<J=��;=A=��=?�<G��� ���,��Dt�,Y������#�"*K�lq�ԭ��?�������⢿�(�� ˗�����s���L��$�����v���ɪr���ׅ������<4�a=#�=0֌=�x=�   �   �>�=��Z="�=@f(<ȧg��=��Vu�����=��OĽ7�½�������nk��o��ǅ����;\!�<$!=�QG=��V=��C=*e= s�;z��H�νh�=�#ۖ���۾w���(B��o�ˍ�i.���w���U���ܽ������
���ѡ�xX��+zp�NnB����8ھB��� 6�������ƼD��<��^=C�=�;�=o��=�   �   2!�=�<�=��=�VB=���<��G<��{�x)����ټB��T~�����٤� B��D�;T�<�� =�e2=�:X=*%l=+g=�A=L�< ����xd�ts���b�Ni��������+�r8]������S��"ӵ�<�ƿ��ѿĎտ��ѿ�&ǿv/��Ɉ��A���8�\�}�*�ֶ�� :����W��(�R*��܀<<EX=m��=���=|�=�   �   �>�=���=���=�Q�=~Yt=^�==�\=���<4��< 1:<�$<� C<���<��<FF=�_'=ΨK=��j=�|=Mށ=�8p=j<=p��<Xyo�%g�����'��P�ľOS�=��{r������خ��ƿFؿx�*�G,�uoؿZƿx����<��>q��l;�+&
��%��:�r��'�l�I� 9<8�P=�ٟ=��=���=�   �   ~��=��=�#�=��=B��=�Z�=��d=$�@=�s%=d�=8=��=�	=p�,=� D=��]=P�v=���=h�=h`�=D�t=��7=�J�<���������_#������Ѿ>��!+H��	��
���`���Zп�{�u�￣�����Nw㿕-п���#	���Q~�1�E�T�~D˾F遾6���,g��P�;�K=���=n^�=���=�   �   ���=��=�c�=Ԯ�=�M�=�\g=�;=�=���<b�<x��<�2�<<�=�)=X�K=,o=Z��=�c�=���=��=q}=��(= ��;ʴ<�����ij��T��W�3�F�����P��a)˿�����R�%S����Q�Z@����l�쿵ʿ���J���6�C�\�
�ͷ�)4\�q۽0e꼰'�<R��=歮=:9�=�   �   L��=}��=�l�=��=�8z= �F=Z�=�>�<Dת<hq�<TR�<x��<���<��	=�*0=(X=bg}=�B�=j��=%��=d�z=�g)=p��;�a3�C���d�>E��v7��;C�v����k���ǿ������7��i���w�b�������������ƿ�C��m��Er@��H�w���W�uԽ�,ۼ�3�<:F�=�a�=� �=�   �   ���=�=
�=�nc=a#=�T�<�&< w��Ș�h>]���X�H���9Z��"<��<�=<�D=�n=4ф=���=hmq=�+=P�4<����ݽ�pT������h8���u�����ƽ�J޿D�������5�9���N���������ݿ�=���3���s�V%6�W� ����2H�SM��ȯ���<+}=�A�=X��=�   �   �{�=<gz=��5=�k�<�JQ;(���xi��aU��2��c��T���0r�HqA�
� ���X�C�;0��<�H#=p S=�j=9`=ښ+=���< i�	���;��,��Ϸ�P�'�A.`�BՎ��/���#̿`�������������2��%&翡l̿$(������*	_���%���$Η�d�0�����0�\��,=D�u=A��=���=�   �   �;P=`�=�e�;�j��j�P��[��B`ڽ�����|��h!���	������ں�����@:�8O<�=��4=0=D=T�'=HK�<�{��!����n��є̾
���D�m|��I��N���'Ϳ��߿�6���d�쿸�࿍ο���I����\|��D�e�[^ʾ?���P���}��z��X=�g=bl�=�+�=�   �   ��<x����1�ϼ��Z ��q*� _P�L�n�L������NL����u��4Z�^�6�u��ǉʽ:�t� $ɼఖ;��<�:=�w=���< - � �G�_�)V�#}��g��q�%���U������O��k9������7j˿�NϿ0�˿����^��
e����H	W��m&�$���̧�NS����`L,�Ћ�;B�=�=P=��T=�)=�   �   p㎼��q���޽D(���c��=����������̾�
Ҿ�fξ^¾5i���,���_q��6������}������@��:l��<�=���<�*"<$�Ӽa;��0� �r6������ޡ�,�-�ָW�����Ǒ�!۟�T����V��:����⠿��
A���Z���/������þH���� ������е�X5~< =V�,=��=��f<�   �   䄽�R��d�B����e����Lؾ�����:���}����k �0j �|޾�۶�f���O�����K���#���;���<t5�< h�<�����v=���ٽ�N>����H�̾;�^)��
J�Jfg�Z�~��膿嵉��u��vW����i�;�L���+�xg	�	�оF���L�B�����B� ?}�p�<$6=���<�kE<�^���   �   �����J��S��~ƾ������ Y/�&�A�
N��R�gO���C�b�1�Z���� �O̾�i���S�]��ṡ�������@<`��<�H�<`�n<�ou��v��x����J��O���yƾ����k�`U/�K�A�N��R��O�&�C�8�1������ ��
̾�f���~S�v���ȇ�@����@<�}�<�@�<xdn<@�u�|�v��   �   sT>�����ر̾��)��J�Tjg���~��ꆿ����w��dY��A�i�:�L�;�+�xi	��о����s�B��ས�B�`\}���<\9=<
�<ЎE<�E���ۄ��G����B��
������GؾU����7�����P�`��vg ��޾�׶��b��'	O�5���F������;���<41�<L^�<`܎���=��ڽ�   �   z9������Y��-.�V�W�����ɑ�_ݟ������X��`����䠿����B��iZ���/�^���þ�	��� �r���<յ�`6~<�=�,=��=�'g<8Ȏ�(oq���޽v=(��c�R9�����j���y�̾YҾ�aξi¾�d��)��JYq��6����x��`���@Q�:��<�=P��<"<��Ӽ�A���� ��   �   K���~����%���U�\����Q���;��̻��ul˿QϿG�˿����`��~f��C���7W�o&�A&��VΧ�>S�)��^N,�p��;@�=�AP=��T=P�)=�ë<(��^�1�g����S ��j*�HWP�	�n��������.H��K�u��-Z�_�6�u����ʽ̽t��ɼ��;�<<<=�v=Ը�<@� �z�G�!��;.V��   �   �̾
�#�D�^|�dK���O���)Ϳ��9���L��q��ο���U����^|�C�D��e��_ʾ���Q��}�@�z�:Z=�g=�n�=�.�=`DP=	=p��;PK���P�lQ���Tڽ������/��R��	������k������p�9�`0O<=(�4=�=D=��'=�C�<�*{��&�����	���   �   ���&�'�0`��֎�:1��\%̿��֥�������n��4��V'翜m̿�(��F���
_�I�%�_龚Η�׿0�,���h�\�|.=�u=��=2��=�~�=oz=2�5=0��<�R;�j��jY��PU��)�������}��xor� cA��� �x�X�p��;��<TM#=XS=�j=�8`=�+= ��<@u�v���;��.���   �   ��>j8�g�u�����ǽ��޿����z���6����NO����������ݿ>��+4��|�s��%6�s� � ���H��L�� ů����<`-}=C�=��=ҝ�=n��=7�=,vc=�i#=�g�< �&<@��`l�X]�x�X� ���X�x#<�!�<�=��D=��n=�ф=.��=�lq=�+=��4<��p�ݽ�sT������   �   f8��<C�"����l���ǿ���D�����η�Rx�������ʱ�����ƿ�C��	m��r@��H���W��sԽ�'ۼ8�<NG�=�b�=."�=���=��=hn�=��=.=z=�F=��=xI�<<�<|�<`\�<���<���<Z�	=@-0=, X=�h}=�B�=}��=״�= �z=�e)=�k�;|f3�LF��d��F���   �   ����F���Q���)˿�����R�5S���}Q�>@�|����Tʿ���쭂���C���
�5̷��2\�<۽x^꼸,�<M��=���=�9�=R��=C��=:d�=J��=1N�=f]g=��;=��=@��<0b�<0��<L2�<��=p�)=��K=Do=���=[c�=��=�=To}=��(=��;<�<�a���>kj��U���   �   �7� <C������k���ǿ��鿴����&���w���Q��>�����1�ƿ�B��wl��)q@�H����	W��qԽ�"ۼ�;�<�G�=8c�=l"�=п�="��=zn�=��=8=z=�F=��=�I�<\�<L|�<�\�<���<��<��	=�-0=� X=Di}=GC�=ڄ�=J��=<�z=2g)=`|�;�c3�=D��d��E���   �   ��qh8� �u����(ƽ��޿|���O��]5����N�f��������ݿr<���2��J�s��#6�$� �;���lH�$I��4���\��<�/}=�C�=���=$��=���=Y�=Vvc=�i#=�g�<h�&<@���k��]�H�X������W��#<�"�<��=��D=��n=�҄=���=�nq=�+=��4<�����ݽ�pT����   �   �쾪�'�U-`��Ԏ��.���"̿,�濤���P��������0��r$�	k̿�&��d���_���%����˗�(�0�����|\�43=�u=��=���=M�=�oz=��5=���<�R;�j��JY�bPU��)�������}�� or�zbA��� ���X����;���<�N#=&S=j=�;`=ڜ+=���<�e����;�,���   �   |�̾�]�D��|��H���L��^&Ϳ��߿5����T�쿭�࿖
ο�
�������Y|���D�c�B[ʾ���rM���}� 4z��_=вg=�o�=�/�=TEP=�	=���;�J����P�XQ���Tڽ������ ��9���	�p��>���޲��L��@�9�x7O<B=��4=$AD=��'=Q�<�{� ��C�����   �   �{��!����%���U�^���?N���7������#h˿�LϿ��˿ϱ���\��c��N}��@W�k&� ���ɧ�uS����A,���;|�=�EP=��T=�)=ƫ<����1�G����S ��j*�@WP� �n��������� H��&�u��-Z�"�6�*���ʽ$�t��ɼ`��;�<(@=&|=D��< ��H�G���>'V��   �   �4��E���?���-�D�W���� Ƒ�*ٟ�4���KT������Z࠿�	��?��_�Y���/�P����þ/��D� ����� ���\~<=Z�,=��=�.g< Ǝ��nq�y�޽f=(��c�N9�����f���u�̾RҾ�aξV¾�d���(���Xq�l6����w��|������:��<=��<`="<��Ӽ�7���� ��   �   dK>������̾3
��)��J��bg���~��憿�����s��VU����i���L�t�+��d	�k�о������B�����B� �|���<�?=��<��E<|B��Iۄ��G����B��
�����GؾU����7�����L�X��kg ��޾�׶��b���O�����E���p=�;��<�?�<Lr�< m��Vo=���ٽ�   �   Wr��%|J��L���uƾ(�����=R/���A�NN�,�R��O�J�C���1�H���� ��̾�b��mxS�N������h��� �@<,��<TT�<`�n<(fu�z�v�yx��n�J��O���yƾ����l�aU/�K�A�N��R��O�!�C�0�1������ ��
̾�f���~S����cǇ�X�����@<؊�<LS�<ؗn<XRu�B�v��   �   �Մ�*@����B�s������dBؾ�����4�p�����{���Zd �޾�Ҷ��^��,O�����=��L�� }�;���<PD�<r�< ����t=���ٽ�N>�򒑾>�̾9�])��
J�Lfg�\�~��膿䵉��u��tW����i�2�L���+�ig	��о�����B�u
���B� �|�$�<H>=<�<�E<D4���   �   X���"bq�H�޽*8(���c�w5������z���-�̾��Ѿ\ξ¾�_���$��8Qq��x6�y����n����� ��:Ф�<"=x��<X;"<��Ӽ�:��� �`6������ڡ�*�-�ָW�����Ǒ�#۟�U����V��;����⠿��A���Z���/����|�þ���� ������ɵ�I~<=��,=��=�Eg<�   �   �ӫ<X`� �1�����N ��d*�_PP�^�n�刁�z����C����u� &Z�>�6�(���vʽ��t���ȼPF�;�-�<2E=4=���<@���G����V)V�}��^��m�%���U������O��l9������7j˿�NϿ1�˿����^��e����@	W��m&��#���̧��S���佌I,� ��;��=�EP=��T=~�)=�   �   �JP=�=��;2����P�mH���Jڽ�������������	�!�����쩇�&��(�9��_O<�=��4=&ED=�'= S�< {�� ��H�\��Ȕ̾���D�l|��I��N���'Ϳ��߿�6���e�쿹�࿍ο���H����\|���D�	e�?^ʾ���P���}���z��\=
�g=�p�=71�=�   �   ��=�tz=\�5=��<��R;�Q��K��@U��!������u��,^r��RA��� �XtX��;�	�<,V#=�
S=`!j=�>`=�+=H��<xe�o��p;��,��ɷ�N�'�@.`�BՎ��/���#̿`�������������2��&&翠l̿#(������%	_���%���
Η��0�/���0�\�0=��u=E��=���=�   �   
��=��=j�=�{c=(p#=@w�<�'<�ൺ B�(�\��`X� \� fU��C#<D3�<��= �D=��n=�Ԅ=���="qq=�+=��4<p��&�ݽ�pT������h8���u�����ƽ�K޿D�������5�:���N���������ݿ�=���3���s�R%6�P� ����H��L��0ů�4��<�-}=�C�=���=�   �   ���=���=?o�=3��= @z=��F=��=�R�<4�<���<Lg�<|��<H��<^ 
=�10=�$X=�l}=�D�=��=f��=D�z="i)=���;\a3��B���d�<E��v7��;C�v����k���ǿ������7��j���w�c�������������ƿ�C��m��Br@��H�n���W��tԽL+ۼ�5�<�F�=�b�=K"�=�   �   ���=�˯=�O�=�j�=�&W=�`!=���<�9�<H�4<��<��<�/Q<��< O�<<�(=��W=�a�=�]�=)�=kː=L�l=zd=`-�Z⚽*%.�r��������4��vy�8��)Sο�n����y�$�Mt4���>���B�Y�>�KW4��r$��C���F�̿=P���v���0�)������i"��l�� �;�;=Ǔ=�g�=�   �   o�=셦=��=�4p=x]5=�V�<�Ɋ<�(�;�]� 5���T[��n�:8�<U�<Z,=t�;=��k=L{�=郑=x��=�hh=ƛ=��������)��%���𾟮0�\�t��<����ʿGF���5��!��C1�};��?�&�;�z;1���!�������eOɿ����o�q�s�-��A�����G�LX{���K;D:=m/�=���=�   �   ���=�;�=�^]=��=��< Hs:�|���zw�j)��#��'	���� ���<t��<��%=|�Z=I{=&�~=C[=
�=�-��!������;��Y��ڽ&���g�}󘿙����:�'����s)(�ݲ1��5�2�1��T(�^��9���}�����¹��FEe��1$��ܾn9��%Y��)`�@<�;�7=��=%2�=�   �   ��l=��2=���< �W9Ġ̼�K��t��,&��A�н��ڽ��սyM½B.���q�Fr�x�A��O3<�?�<�a6=�1Q=B=C=J� = �z���]�S���{��H˾^>�WS�����밿�vֿ�z��8[��W�S�"�'&�5.#����>�������jֿ+~��hK���Q�e�dǾ~s�"����7� �<8�/=<|u=�=�   �   Z�=��<�{��:�_�Y���k ��� �Ϊ:���K���R�&�N��?��=(���	�ާν�X��^�@�]�Hg�<��=j=��<��;��$���߽~U��
��ٝ�(L9�k�v�H���@�����޿Ʀ���F	���R��$���	�
�����߿.2���휿͞v�މ8�����n��~�N�h�ѽ�;���X<� =�I= <=�   �   �ho������������9�vl����n�������A�� ���B������U�u�"�C��@�X����J��i� 8<�e�<���<ȵ<��ѼN�����)��k��۾���ohQ��ǅ��t���ʿ���ؿ�����?T��\��e�� \ڿ63��Z���Pu���R�&��Hrھ���Q.&�LU���񡼤*�<�?=�;=$ �<�   �   �bJ���̽�R$���i��d�����2ݾ�������~�-�������p4¾1ܞ���t��.�݇�*?o�$����_�;@u�<�VB<h�>� �c�����U�]����������@*�,][��䆿o���`���9ſn-п�:Կ��п�ƿT ��:����>���e]�B�+��S��i6����]�����F Y��I��j�<��<�^< <6��   �   ��ٽ��4�턾�d��2�{F�k� �M2�v�=���A�X�>��&4�nr#���/��,ƹ�)Ӊ�VW=����vl�����g�;h�B< x�94����R��53�g���r������,�pU��N}�-R���J���_��)������^����ޑ�PA��	[X�-}.�����C¾�`���a!�J�������&�: 3p<H/<�aN���R��   �   c�2�nn��.¾�b �>!���@��]��rs��������󞁿��u��_�<�C�O�#�����kƾ_��I{8�]ս^�B��@'�Hg<_<�x	�:T6�=\̽��2��j��I���` ��!���@�[]�ns�k��J���������u�4�_���C���#�A��[hƾ����w8��ս��B�`9'�b<�L<�	�|`6��d̽�   �   Ə��ܓ����,��sU�pS}��T��.M���b������|����������!C��^X��.�~���F¾�b��rd!�T������@8�:pAp<0J<P8N��R���ٽ8�4��脾�_��;�C��� �I2�S�=���A�^�>��"4�o#�	�S��C¹�&Љ��R=����bl���� p�;��B< ��9����Y��,8��   �   p���d����C*��`[��憿���{c��i<ſ)0п�=Կw�п}�ƿt�����u@���g]�0�+��V��l8��b�]�����&#Y��I�Tp�<h�<'^<�6�XRJ�0x̽ZL$���i�`������,ݾ>���h������
����ᾬ/¾6؞�G�t��.�����4o�P����x�;du�<�JB<��>�j�c�U�����]��   �   �۾&���kQ��Ʌ��v���̿�|�ؿ��쿢����V���^�����
^ڿ�4��ψ��{v��wR�z��&tھ8���/&��V�����.�<D=^B=h3�<`�n���?���B��Y�8��	l�9����h������l<������=�������u���C��;�������J� �h�((8<�i�<���<�<��Ѽ������)��n���   �   ����N9�j�v����C��� �޿0���*H	�P�����G%���	�����`�߿m3���P�v���8�[���o����N�j�ѽ�;�X�X<�� =h�I=|<=,�=�<X\��bu_�G ��Qe ��� �W�:���K��R���N��?��7(�U�	���νOQ�����B]��r�<��=�j=��<P��;<�$�s�߽�U�����   �    @�UYS�2����찿Zxֿ�|��I\��X�u�"�?&�6/#�t�����#����kֿ�~���K��ħQ��e��dǾ�~s�y���H7�8�<*�/=h�u=��=��l=�3=4�< (e9��̼X�K�k�������н �ڽ��ս�C½�%���q��e�XgA��o3<XK�<�e6=�3Q=<=C=D� = �{�Т]�����{�0K˾�   �   X�&���g��������O<��'����T*(���1�[5���1��U(��������~�\��� ����Ee��1$�)�ܾc9���X� (`��L�;n7=��=*4�=c�=�>�=,f]=��=P��< v:��{����
j��\)�F�#��	�d������ $<���<��%=УZ= K{=��~=FB[=ƅ=�N��E$��Z��V=������   �   ��0���t�O=����ʿDG��&6���!�LD1��};�.?���;��;1���!�������\Oɿm���/�q�0�-�}A꾤����F��U{� �K;�F:=�0�=P��=��=���= ��=�9p=�b5=`b�<l֊<�\�; m[�p��@�Z�� �:؞<\]�<�/=�;=��k=�{�=��=8��=Lgh=n�=`��������)�A'���	��   �   W4��wy�����Sοo��S����$�st4���>� �B�E�>�&W4�sr$�������Л̿�O��v�H�0�
��6���2h"��j����;0";=ȓ=�h�=6��=d̯=#P�=3k�=�'W=na!=��<�:�<��4<�<0�<H.Q<��<�M�<\�(=��W=a�=]�=��=�ʐ=n�l= b=�-�m䚽�&.�Y���$����   �   �0���t��<����ʿ7F���5���!�~C1��|;�M?���;��:1��!� �����Nɿ�����q�Z�-�F@�˅���E��R{��L;�G:=1�=���=(�=ԇ�=6��=�9p=�b5=pb�<p֊< ]�; j[�0����Z� $�:��<�]�<0=Z�;=0�k=|�=g��=���=lhh=��=8������ç)�\&��<��   �   ��&���g�<�5���Q:鿣&�p���((�$�1��5�U�1�T(����u���|�¬������wCe�_0$�أܾ�7���V�"`�0l�;7=y�=�4�=��=�>�=`f]=�=x��<�v:@�{�����i��\)��#��	�����(���%< ��<^�%=��Z=FL{=R�~=jD[=Ĉ=�+��!�����;��:���   �   �=�QVS�K���_갿�uֿ�y��zZ��V�T�"�&�-#�|��4�����iֿ�|��J��ؤQ�cc�|aǾ7zs�R����6�P�<О/=Ђu=��=��l=`	3=��< be9l�̼<�K� k�������н��ڽ��ս�C½[%��Bq��d��cA��s3<�M�<:g6=�5Q=4@C=x� =�#z���]�Ŀ�@�{��G˾�   �   ��K9���v�D�������:�޿����E	�������"�`�	�������߿30��윿ݛv�x�8�����k��>�N�
�ѽ�1��X< � =B�I=8<=V�=��<�[��8u_�@ ��Ne ��� �X�:���K�ߧR���N�
�?��7(�0�	�I�ν�P�����+]��v�<~�=�n= �<�4�;��$���߽U��	���   �   "۾E���fQ��ƅ�	s���ȿ���ؿâ�i����Q��ZY�����zYڿ�0��B���|s���	R����lnھ���)&��N�� ܡ�|=�<�H=~E=H7�<��n�b�����5��Q�8��	l�7����h������i<������=��������u���C��;������J���h�P38<�q�<��<��<�}Ѽ������)�cj���   �   ���������>*��Z[�Pㆿ�
���^��b7ſ�*п88Կ.�пr�ƿ����ᡠ��<���a]�>�+�O���2���]������Y�(�8�<T(�<�3^<@6�*QJ��w̽BL$���i�`������,ݾ?���h������
��s�ᾗ/¾؞��t���.����2o�����p��;���<@kB<s>���c�G���L�]��   �   E���������*,� mU�cK}�P��UH��w]������d��Ѕ��0ܑ�?��WX��y.����w?¾V]���\!����������:H^p<8]<@,N��R�8�ٽ�4��脾�_��7�C��� �I2�T�=���A�[�>��"4�o#���;��$¹��ω��R=���转l�H���P��; �B< \�9����8N��#0��   �   ��2��g�������] ��	!���@���\��is�'����F����u���_���C���#�9��acƾ����wq8�սޟB��'�Ў<xy<�g	�~Q6�f[̽A�2�j��?����_ ��!���@�\]�ns�m��J���������u�/�_���C�v�#�3��9hƾ���7w8�lս��B�x%'��~<`v<�]	��K6�qV̽�   �   ��ٽ��4��儾�[��d�2@�[� �jE2�a�=�j�A�<�>��4�Lk#���F��"����ˉ�!L=���轞l��萼�̸; �B< a�9�����Q���2�N���d������,�pU��N}�/R���J���_��*������]����ޑ�MA���ZX� }.�����C¾�`��Wa!������� ��:�Wp<xc<�N���R��   �   �FJ�ap̽DG$�F�i�)\�����"'ݾ7���+���������V��*¾NӞ���t�=�.�qu�(#o��k��@��;���<@tB<�t>�ڙc������]����������@*�+][��䆿p���`���9ſo-п�:Կ��п�ƿS ��7����>��xe]�6�+��S��D6��P�]�F����Y�`4�dz�<�)�<@B^<��5��   �   �n����0���4��'�8��l����Od������07��� ���8����@�u�R�C�h5�×����J�0�h��W8<L~�<ػ�<��<�~Ѽ���]�)��k��۾���ohQ��ǅ��t���ʿ���ؿ�����AT��\��e���[ڿ43��X���Lu���R���*rھ����-&��S�� 顼<7�<�H=�G=�A�<�   �   |=�< D��<f_�����_ �f� �q�:���K�4�R��~N���?��0(��	�N�ν�G��N��g\����<��=�s=H&�<@@�;��$���߽>U��
��՝�&L9�l�v�H���@�����޿Ȧ���F	���R��$���	�	�����߿+2���휿ƞv�Չ8����qn���N�O�ѽJ8���X<�� =��I=�<=�   �   ��l=f3=P�< �o9 h̼0�K�gb��M��[�нd�ڽ��սs9½�����p�pU�0/A���3<�_�<4n6=(;Q=DC= � =��y���]� ���{�}H˾\>�WS�����밿�vֿ�z��8[��W�S�"�)&�5.#����>�������jֿ)~��fK����Q�e�dǾ�}s�W���� 7��<8�/=$�u=��=�   �   ��=�@�=Hk]=B�=��<�qx:��{�L��^]�xO)�ܙ#��	�d฼�W��M<t��<�&=��Z="Q{=8�~=rG[=0�=���] ��ʳ��;��S��ڽ&���g�}󘿘����:�'����t)(�޲1��5�2�1��T(�_��8���}���������AEe��1$��ܾ[9���X�(`�N�;7=?�=05�=�   �   `�=l��=)��=H<p=>f5=�j�<��< ��;��Y��·���Z���:�< i�<25=��;=<�k=�}�=慑=�=�jh=N�=���������)��%���𾞮0�\�t��<����ʿFF���5��!��C1�};��?�'�;�z;1���!�������dOɿ����l�q�p�-��A�����G��W{� �K;�E:=�0�=p��=�   �   ��=Dw�=���=��T=�=���<h�<@������XSH� e2�`�����;� �<��<��3=f�g=��=$Ԏ=!<�=ʣM=xx�<x�����ܽ�a��������Z��1���'Ŀ����PY���-���E�nZ�!\h��Um�IVh�vCZ�ЍE��"-��]�eb��¿�<��[vW����M���TX�m˽�[����<�Tr=��=�   �   ��=�Ў=�p=�3=@u�<��8<@�]�x�x�\뼼pؼ V˼8��ȟ�@�;��<$�=ʢL=�x=��=R�=�iH=t;�<�����ֽ�v\��p��D���V�����^���
u������*�K[B��9V���c�n�h���c�T,V�3B�?*�� �9���޾�������S�P��et���\S��cŽ�ݪ�$��<�l=a��=�   �   Dy�=��\=H=��<@����0����(���e�&U��ҙ����Bvt��r=���� $�O4<D�<��8=��^=�b=��7=X۟<��м�Ž*CM�^����0��$K��ߋ��&��^���
�V'"��8�hYJ�@�V��H[�B�V���J��8���!��(
�C�F���2m���uH�����K��4E�c���Q���b�<TuZ=��=�   �   $/=���<`�V;�tżPzZ�����&�ܽX��W���
�t���o����Wq���y�b��@��d�<J�=��+=�3=4��<�y��91���5����]���a�8������Mӿ��z����(�0�8��C���G�]�C��;9��(��)�����̋ҿy3��C�}���6��&���d�.�}9���~U��<&:=d�L=�   �   ?O<�g��G��д��_��z/�ZXU�v�s�σ�����+���Cx�8c[�!�6��i���Žzi�80����;��< ��<�]}<( i�����U��,���jcھo�!�{a����������}�����y#���,��(0��6-��@$�(g��!�u������Ԉ��aI`� � ��׾-��:[�
`|�������<BT=Ȼ�<�   �   ̋�E��{��M?5���r�p��������kȾѧ־�	ܾ�ؾ}�ʾ8�������{� >��0�,����$����#<�<2�DVN�����f^��派��dx>��}�@à�Uÿ>]� � �d���W��9�����y����%濬�Ŀ�����5~�ҍ>��0�?����C[�� ;=��ᔻ��v<��<�DC:�   �   �s������XZ�9m��v���8
쾥 	�T%�D"���%���"�����|�𾳓ƾ�����b�LU�2����,���I� ��8`k׻�>�E���x*�_���پDg�~O�$���\���0��h׿��w����^��U����f�wٿ���X���������P��0���پK���K)��B���@� �P�@��; ������   �   �*�-`m�W��x�ᾆ]� +��D���X��8f��)k��Mg�v�Z��1G���-���~��R����jt�����Z��f�(��fg� �X����j������R�yפ�t��@p"�g�Q�|&��7t��D
���M����ǿ/�˿h�ȿ�ʾ��ܮ��I��Ă�HDT�P$�7;�!q���~T�p>��i�����|��0r:��4�v���   �   n�j�#|�����!'���D��j�I���6���r2���^��4᛿C铿�"���Tm���G�z� �����n���Eo���������9��<���5���������u�j��w��-��#�[�D��
j�����~����/���[���ޛ��擿� ���Pm�Q�G�ʺ �����U����@o����g���V7�H�<��5���
�����   �   vۤ���s"�c�Q��(���v����zP����ǿ5�˿O�ȿU;�:߮��K���ł�/GT�HR$��>�s����T�(B�(�i����\���S:��(��	���$��Xm�&R������Y�+���D���X��3f�	%k��Hg��Z��-G��-���ҵ澵����et���V���(��`g��"黠d����j�	��R��   �   �پj���O�D������n3��_
׿'�꿬����a��\����i��ٿ���'���'�����P��2��پ�L���M)�iD�� A���P�`��; �����9j������PZ�kh����������s!�A"���%���"�@���������ƾ�����b��P����B�,���I� 0�8��׻$F�K��~}*�9b���   �   <��W{>�=�}�eŠ�|Wÿ�_俠� ����qY�l;���{� ��0 �_�ĿV����7~�h�>�2������E[���d;=�0ϔ��v<���<�F:n輣���n���75��r�`�������eȾ��־Mܾ� ؾ��ʾ3��������{�%�=��+�O락\�� �����#<<�B�T^N�0��k^��鴾�   �   ��!�X a�ȵ������c����K{#�+�,��*0�58-�FB$�?h��"���!»������J`�� �K�׾����[�.`|����؝�<fZ=���<�lO<��f��	G��Ŵ�$Y�Bs/�PU���s�tʃ�🇾������w��[[���6�jd��Ž�i�����Q�;���<���<X}<�i�ޟ����������fھ�   �   t�8�~�����$ӿ0
������(���8�Y�C���G���C��<9���(�W*�������ҿ4��$�}�}�6�~'��𛾤�.�59��wU���<�:=��L=l,/= �<�_W;�UżhZ�������ܽ?������Y��,j�X��Yh���
y� ���ȧ�r�<��=$�+=�3=�}�<H���Q5��4�5�Ɓ��}����   �   �&K������'�������
�L("��8��ZJ�e�V��I[�6�V�K�J�$8�!�!�)
��C俎���]m���uH�����K���E����`M��Dh�<�xZ=C�=*|�=��\=�&=3�< <�����J�(���e�=M���������&ht� f=��������l4<�O�<��8=2�^=Үb=��7=X֟<��мŽ�EM�X���2��   �   \�V�a���P���v���+�*��[B�z:V�N�c��h�a�c��,V�eB�?*�� �.�￫޾�����9�S����s���[S�bŽت�x��<�l=쓓=ݶ�=�Ҏ=bp=x�3=���<�8<�G]�yx��ۼ�X�׼�G˼�*������;��<D�= �L=Z�x=��=�=hH=06�<���ֽ$y\�Nr��Q���   �   ��Z�l2��`(Ŀ;����Y� �-��E�KnZ�<\h��Um�.Vh�FCZ���E�D"-�V]��a�n¿�<���uW�^���L��SX�˽�T���#�<�Vr=��=ң�=�w�=���=��T=�=���<��<����H���RH��e2������;d�<��<n�3=6�g=��=gӎ=C;�=��M= s�<������ܽ��a�%���P���   �   W�V�����y���u����g�*�[B�l9V�&�c�ؚh�>�c��+V��B�b>*�f �4���ݾ�𺑿?�S�L���r���ZS�8`Ž8Ӫ����<�l=;��=��=�Ҏ=�p=��3=���<��8<@G]� yx��ۼ�P�׼�G˼�*��0��@�;,�<x�=P�L=��x=4�=��=>iH=�9�<���/�ֽ�w\�@q������   �   �$K�gߋ�;&����ƣ
��&"�8��XJ�K�V��G[�"�V�h�J��8���!��'
��A����$l���sH�g���I��PE���(D��<n�<�zZ=��=�|�=&�\="'=T3�<�8�����D�(���e�<M����������gt��e=���x���n4<�P�<h�8=L�^=Z�b=
�7=�ܟ<0�м�Ž8CM�X����0��   �   ��8����T��mӿ�������(��8���C�-�G���C�*:9���(�z(������ҿ�1����}���6��#��p훾�.�\4���]U��'�<�:=��L=x-/=4�< eW;pUż�gZ�������ܽ@������T��!j�3��*h��N
y�z��`§�(t�<j�=J�+=�6=��<�u��A0��q�5��������   �   z�!�"a� ���P�������|�s��ux#�!�,�d'0�-5-�u?$��e�W �&����������F`�� ���׾����W��T|� ��ܧ�<�]=���<PqO<��f�*	G��Ŵ� Y�Ds/�PU���s�xʃ�򟇾������w��[[�~�6�Gd���Ž�i�@���_�;� �<��<�m}<@�h�͙��#��M���bھ�   �   Ȅ��v>�s}}�����OSÿ2[��� ���OV�88����'x�O��j�<�Ŀ؊��12~��>��.�Я���>[�U
꽸.=�P���(�v<�<��F:|k�A���n���75�
�r�a�������eȾ��־Mܾ� ؾ��ʾ�2��}���Y�{���=��+��Ᵹd�� ྻ��#<�"<�6QN���d^��䴾�   �   �پ�e��{O���������.���׿D��{����[��&����c쿀ٿ��矣������P�.�8�پ�G���F)��:��4��P�`�;��������i��S���PZ�eh����������u!�C"���%���"�<�������܎ƾ�����b��P����z�,���I� d�8�=׻�8�]A��pv*�6]���   �   �Ԥ� ���m"���Q��$��r������J����ǿ0�˿^�ȿ�Ǿ��ٮ�DG������H@T��L$��5�m��hxT��4���i�D袼�� >:��%�����$�ZXm�R��|���Y�+���D���X��3f�%k��Hg��Z��-G�
�-�����澔���+et�����T��(�(��Ig�0��K����j����&�R��   �   ɐj�at������ ��D�j�~������-�� Y���ۛ�	䓿���Km��G�6� ���������e9o�R���}��)���<�p�5����;��{��4�j�w��$��#�]�D��
j����������/���[���ޛ��擿� ���Pm�I�G��� �����1���A@o�J�������1�X�<�0�5� ����������   �   � ��Rm��N��ٽ�"W�� +���D���X�
/f�8 k� Dg�W�Z��)G� �-�[���澺����]t����`L����(�X,g�����J��r�j����_�R�_פ�f��>p"�f�Q�}&��8t��F
���M����ǿ0�˿h�ȿ�ʾ��ܮ��I��
Ă�=DT��O$�;��p��~T��<�F�i��󢼐*���6:�������   �   Uc������JZ��d������������l"���%���"�\����-��"�ƾ����b�kJ�ĝ����,�ГI� �8 (׻H9�MC��nx*��^��vپ@g�~O�%���]���0��i׿��z����^��U����f�uٿ���U���������P��0���پ�J��K)��@���:�`FP���;�~������   �   X�[���ve���15���r��������_Ⱦ��־�۾��׾��ʾ]-��k����~{���=��%�᝽Ė�������#<�5<���QN�[��ff^�v派��cx>��}�@à�Uÿ?]�!� �e���W��9�����y����"濪�Ŀ�����5~�ɍ>��0����uC[���J6=�������v<PȂ<�H:�   �   ��O<��f�f�F������S��l/��HU�l�s�ƃ�c���'섾�w�gS[��6��]���Ž��h�X���P��;d�<���<�|}<`�h�����������Zcھk�!�|a�	�������	��}�����y#���,��(0��6-��@$�&g��!�s������ш��[I`�� ��׾����Z�v\|���`��<_=t��<�   �   <2/=D�<��W;=żYZ��맽��ܽ����|�A����d�ӥ��]���x����Z����<��=��+=j;=T��<r��	0����5�l��O���^�8������Nӿ��{����(�1�8��C���G�^�C��;9��(��)�����ʋҿv3��>�}���6��&�����.�98���oU�0$�<�:=�L=�   �   �}�=D�\=�,=0B�<@��� ��ʻ(���e��E��5�������Xt��W=������8�4<�a�<v�8=��^=�b=��7=��<��мŽ�BM�O����0��$K��ߋ��&��^���
�V'"��8�hYJ�@�V��H[�C�V���J��8���!��(
�C�D���0m���uH�����K���E�����L���i�<dzZ=m�=�   �   W��=pӎ=�p=��3=���<@�8<��\��_x�μ���׼�8˼����k�`A�;H*�<�=�L=��x=��=�=lH=?�<X�５�ֽ�v\��p��C���V�����]���
u������*�K[B��9V���c�p�h���c�T,V�2B�?*�� �:���޾�������S�M��[t���\S�:cŽ8۪����<��l=��=�   �   H�=�Є= H]=(� =���<`�; �� ���<4��� ��z�ܐ����D�`�;X��<�g=�F=V�r=�I�=h�p=D_)=�?�;:�P������澢�1�ت��.���a�Ӄ�%�+�V�J��i�����Ŋ��������B����|h��I��a*�Q@�t�߿$���)|�a�.�"P⾔��w'���7���M<@�@=�"�=�   �   }
�= �q=J�>=t��<(�A<�_λ�����5�&C��Y:���Lռ��,��o�;��<L5(=��Z=��r=�/e=~G#=@��;�J��~�w膾bV��..�d{��/����޿M$�E�(��F��hd���}�Kć����fʇ���}��d�,'F�_�'��
�iܿk=����w�3v+���ݾt�����>)2���J<j:=2P|=�   �   ��S=�h(=�.�< �;X���d�7������Ĩ�-?��
�ǽ�½K1��R*���J��aڼ _�@��<Vj=��<=�A=�(= ��;�s9�Tt��h|���Ծ�l$�_�m�/y��!�ӿ
K� �z8<�eSW�l�n��~��?���~���n��fW�p�;��t������ѿ>��j��"�R�о|�u�ө����"�H�><Zr&=��W=�   �   ��<��%<�D����@��A��J�潺`�L)���8�"�>���:�:e,�������t��FX�,����;�X�<��=:�<`?�;�� �Tp� �a�j𿾠8�=�X�1Ք��i¿6`����7,��C�`%X���e�Yk�Vjf���X�V�D��,�O�����Ņ���ד���V�u�MǼ���[���ٽ�L��<��=<j=�   �   બ��V�����q���U,�_z\�I����+��k�������؀�����i���bb�f�2�N������\�)�HZ-���<�`<�W�:|S�S����Q@�����P �yR>�%p������P�ؿ��7���-���=�04I��tM�)�I�f�>�g�-�����9�H�ؿ�V�����<=�z� ��k��i�;�߶�غ鼠J�;P2�<��_<�   �   �	T�Jʽ�H ��wc�P!��1ɷ���־��ﾑ���v��� �� �hھ�[��uΘ�ގj���&���ս@i�L似�����l��������y��T�ؾc ��c_�A���	6��"p�(��C���Q"��+���.��#,��[#���������<������by_�z �I�׾K ��9��8#��p�ļ@h�� ��<b���   �   �{潾j9�>������)m�P���G"�,�3�z�>��C�۵?��"5��K$�:�����������?e?�����˄�h���t���D?ɼ�g��S�eU�S���w^��&6�:�r��K���\�ۿ�����7���6l��5��1�%����ݿi��
���at���6�������deT��'��_�4S���
d��[༎�x��   �   A�A��ޑ��J̾����(�-ZI���f�(�}�!\��%��`솿���&i�<L�&'+����Rо�ٔ�t&F�m��O���_���м�*��b��z�������ƾ����r?��|u��d��Ұ��"ȿ��ڿ濈��翌:ܿ�"ʿ˲����x��KA�#�I-Ⱦ�؂��B��ߩ�ʍ&�@ż�F ���{�����   �   V���Ҿ+��͛:�~�f�Ɵ��h���<��p߳�ns��c���:������XP��V�i�d"=����}�Ծl��;�9�W�׽Pc��/��|���0_�AԽ/37�V���	Ҿ�����:���f����0e���9��Fܳ�Gp��Y���b���]
��N����i�L=�A����Ծ�����9���׽dc�p2�������:_�YԽ 97��   �   K�ƾ����v?�|�u��g��հ�&ȿ�ڿ9����:�翟=ܿb%ʿ|Ͳ���>x�*NA��$�
0Ⱦpڂ��D��᩽z�&��ż&> �
�{�H�齗�A�,ڑ�&E̾r����(��UI�|�f�ɩ}�]Y��Z"���醿����!i�FL��#+�!��#
оj֔�"F����L��^���м�*�i��$������   �   �`��)6�F�r�
N������x�ۿ ����9����n�C7�&3��'��2�ݿk������Qdt���6���������gT�*�L�_��L��h�c�F���x��p潬c9����v����f辌��^C"���3���>�&C�i�?��5��G$�����쾬�������(`?�zy�HǄ� ~��X���|FɼL�g�uZ�3jU�����   �   �e ��f_�P���y8���rῼ�����S"��+���.�}%,�>]#����������������2{_�� ���׾R!��7��#����ļ@���@���I��,�S�R�ɽ�A �foc�>��^÷�[�־���a���� �9� ���	ھ�V��,ʘ��j�H�&���ս<i��ּ�P騻�򷻈�༁���9���{��5�ؾ�   �   
U>��q��������ؿu�����O-���=�+6I��vM���I���>�� .����:���ؿ�W������==�(� �il��-�;�>߶���� m�;�?�<(�_<�D��6F�*���gd��gN,��q\��ۃ��&��${��{����{������d��b[b��2�0���𥽌�)��9-���<�`<@$�:�X�����U@�c���>��   �   ��X��֔��k¿Pb���9,���C�''X���e�&k��kf�J�X�o�D��,�������z���pؓ�P�V�u��Ǽ���[�p�ٽ�J��!<@�=Pq=4&�<��%<�'��ȟ@�X7��s��.Z�E)���8���>���:��^,����>
�<l��&�W�(��@S�;�c�<��=�:�<�,�;� ��t佐�a��m:��   �   `�m�kz����ӿ�K�	 ��9<��TW��n�l�~�G@��N�~���n��gW���;��t�ˈ��ѿn��j��"�J�о0�u����L�"���><fv&=��W=�S=�p(=0B�< �;�۰�`�7�Y���仨�&6���ǽ9½5)��#��.J��Lڼ��^�h��<
o=��<=�A=�'= ��;y9�rv��k|���Ծ�n$��   �   �{�m0��Ș޿�$���(���F�vid�v�}��ć�	���ʇ���}��d�L'F�h�'��
��hܿA=����w��u+�?�ݾ�����$&2�x�J<,m:=�S|=n�=��q=��>=���<دA<0"λP���l��N5���B��Q:�����>ռ��,����;P��<�7(=.�Z=T�r=�/e=�E#= ��;ƧJ�����醾.X�0.��   �   ̫�M/���b�%��z�+���J��i����� Ŋ��������"���i|h���I�-a*�@���߿����(|���.��N⾰ ��*&���7� �M<z�@=�#�=�=:ф=pI]=d� =輹<p�;�������d3輾� �{򼸑��h�D��u;T��<�f=��F=��r=I�=��p=�\)=�'�;@�P�� ��� �k�1��   �   �{��/��ӗ޿Q$�8�(���F�Mhd��}��Ç�C���ɇ���}��d�e&F���'��
�
hܿ�<��t�w�
u+��ݾ(�����n#2���J<>n:=HT|=��=ȵq=��>=Е�<�A<P"λP���l��T5���B�~Q:�|���>ռ`�,���;���<(8(=��Z=��r=d0e=,G#=���;��J�l��膾�V�1/.��   �   (�m��x��ȗӿ�J�� ��7<��RW�h�n���~��>����~���n��eW�N�;��s����F�ѿ��j�P"��о.�u����&~"�@�><�x&=�W=��S=
q(=�B�<��;�۰�\�7�Y���컨�,6���ǽ8½*)���"��J�,Lڼ �^�`��<�o=��<=dA=0*=���;�s9�bt��h|���Ծ�l$��   �   ��X��Ԕ�#i¿6_�����6,���C��#X�V�e��k��hf�'�X���D���,������
����֓�V�V�Os��ļ���[���ٽdC�h4<6�=0s=t(�<�%<�&����@�L7��s��3Z�E)���8���>���:��^,����
�l����W���� [�;�f�<��=8A�<�T�;�� �Do�I�a��￾-8��   �   bQ>�`o��������ؿ@��&��@-�]�=�e2I��rM�4�I���>���-�z��g8���ؿU��u ��f:=��� ��h��9�;��ض�t��Й�;G�<�`<@:��|E�����Td��iN,��q\��ۃ��&��({������{������d��S[b���2���8�b�)� 3-��<�+`<@�:�O�?����P@���������   �   �a ��a_����x4��3n����݉�P"�Q�+���.��!,��Y#�b��-�����������v_�� �Z�׾_�����Y����ļ���������D����S���ɽ�A �^oc�;��a÷�`�־���f���� �8� ���	ھ�V��ʘ�ʇj��&�4�սPi�Ѽ�PǨ������t�%�������w��v�ؾ�   �   ]��$6���r��I��䱻��ۿ����@6�%��dj��3��/��!����ݿAf���|���]t���6����Ո���_T�?��}_��9��h�c�(>�j�x�p�|c9����r����f辎��`C"���3���>�)C�i�?��5��G$����쾖���z����_?��x��ń�xu��,����2ɼl�g�qO�&bU�G����   �   ѻƾ���_p?��yu��b���ϰ�! ȿ��ڿ}���v��*7ܿgʿȲ�m��^x��GA����(ȾՂ�J=��ש��&�$�ļ.8 �L�{�$��D�A�ڑ�E̾p����(��UI��f�˩}�_Y��["���醿~���!i�@L��#+���
оC֔��!F�b��J���W�h�м\*��^�����w���   �   ����Ҿm����:��f�䚈��b��7��Gٳ�(m��2���M���o��gK����i�6=�����Ծ�	����9��~׽��b�L�������*_��Խ�27�5���	Ҿ�����:���f����2e���9��Hܳ�Ip��Y���b���\
��N����i�D=�5����Ծ���N�9���׽�c� !��ܥ��t'_��ԽR/7��   �   �{A��֑��@̾ƣ�Z�(��QI�
�f�ݤ}��V������憿��|i��L��+����mо�є�F�����C��jO�L{мD*��`�����R����ƾ����r?��|u��d��Ұ��"ȿ��ڿĕ濊��翌:ܿ�"ʿ˲����x��KA��"�-Ⱦ^؂��A�mݩ�.�&���ļ06 �޴{�l���   �   �h�k^9�J�����,a�U��?"���3�}�>��C�Ԭ?�5��C$�(��t��	��������X?��m���� `��उ��,ɼ��g��Q�sdU�,���n^��&6�:�r��K���^�ۿ�����7���8l��5��1�%����ݿi�����at���6���r����dT��%뽒�_�0@��`�c��4�8�x��   �   ��S��ɽ�< ��hc���W�����־��ﾀ���L���� �
�ھ�P��Ř�:j��&�7�ս��h�x���Ђ������Dp༈�������x��7�ؾc ��c_�A���	6��$p�(��D���Q"��+���.��#,��[#���������9������Zy_�n �#�׾ ��h��� ��0�ļ@���&���6���   �   @����9����7Z��.H,�ij\�J׃�,"��v��<���vv������_���Rb�}�2�����好�t)� -���<`F`<�i�:�M�x���mQ@�{���H �vR>�%p������Q�ؿ��:���-���=�14I��tM�)�I�g�>�f�-�����9�F�ؿ�V�����<=�l� �jk����;�,ݶ�0�鼐��;pJ�<p`<�   �   83�<&< ����@��.��I��\T��>)���8���>�J�:��W,���J��a����W�H���p��;$y�<��=�K�<�p�;�� �o佛�a�Q𿾚8�<�X�1Ք��i¿6`����7,��C�a%X���e�\k�Vjf���X�V�D��,�N�����ą���ד���V�u�.Ǽ�0�[�\�ٽzH�,<��= v=�   �   ��S=�u(=�O�<�;�ư��7�8��������-��,�ǽH	½| ������I��1ڼ��]�Ȯ�<�w=��<=�A=>.=@�;2q9��s��h|���Ծ�l$�_�m�/y��"�ӿ
K� �{8<�eSW�l�n��~��?���~���n��fW�p�;��t������ѿ<��j��"�A�о<�u� ����"�(�><�w&=J�W=�   �   ��=d�q=D�>=���< �A< �ͻ��&��b5� �B��H:����x.ռH�,����;̔�<t=(=�Z=��r=�3e=VJ#= ��;��J��~�j膾[V��..�d{��/����޿L$�E�(��F��hd���}�Kć����gʇ���}��d�,'F�`�'��
�iܿj=����w�0v+���ݾd������'2�h�J<�l:=T|=�   �   ��y="f=Ԧ5=t�<�&<����X�ü܈���8��F�r�<��s�"׼�_.�P*�;�t�<_'=�W=fak=8�U=��=@e��"č�z�+�������I��ӏ���¿(���:�5A�r;f���������o��������ؕ��i��f7e�r�?����(e��*����2��y�F�; �朾��&�Vۄ��C��|�=tod=�   �   �}f=��K=l=p��< B� ���>!�~"[�~��F����e���Qb��,+�Pɼ����p<d�=.A==6�W=��H=� =����zg��� (�n����i��^E�K�� ���������c�=�n�a��߂�����ej��6F���p��d���A���v�`�hp<��b��f��ҽ��Ë���B����������"�İ����̺�=aW=�   �   ��*=���<84<��R�X��㸃�>�����׽�h�͒�����2ܽ&��L��H-��?�����;���<�U=� =��<ptû����u��������C�:��텿����a�r����3���T��u��-��m�������1���U��,�u��T�E�2������Q��������z8�mu�{J���A� �q�@����<D9/=�   �   ��<Pd��l���v����Խj ��40�L�J���[��8b��]�M��}3���%�ܽ4��� �� ����bS<|۵<���<����g�T	��'����ܾ.�)�\�t�w���fٿ���z�$�o�A�C;^��v��փ�b���K��|w���^��)B��~$�v��F�ؿ$���s�%(���پ`݁�6��nX��x��X��<��<�   �   &��J�_��0ɽ@���N�� ��O,��\���߹��{��H����鮾p=��@|��
�S�����ҽ�p���ȼ@?U���;�?��J��8�2Ic��Q��+S��tW�铿tD��o��)+��:+���B�y�V���d��i�(e��W�T�C��,�T���<���偓�kxV��R�n���_�!����=��� f�; h�8�   �   ����$���NgA��+��ߩ���KԾ_���C	��=�̈�����K
����PL׾⬰������nF�������Ƒ� J��<❼p2�d0Ľ��:�S̞�B����B6�18|��ӥ�%oп���%��\&�(F6�A�E�C�A�A\7��'�r�Y���Eѿ�/��<M|���5�����W����Z8�Al��P((��ڈ��-������   �   ���
L]�T��Ӿ�X�?k ���8�%�K�90X�.�\���X�:&M��a:��]"�;��o־mΠ�k�a�Z��^譽��A��7�r�%�Q���$�bN{��^Ǿ�����N� ����@���!ҿ�r���|
��*�^����"��& �\)�t��������ӿ%f��3���ECO����MǾ�~z�L������V����󼤉7��Ч��   �   =f�D奄?�C����?�cd��+��쎿L/���6��L��������^��W�f��A�e��>q�b����i�J.�����`�M��i*�2�s���ؽ�W<���� ��;�!�4�X��p������#ƿj�߿
B���� ��@��A�*���e�῎
ȿ����]���X�Z���"���径�����<���ؽ�4q�>O&���G������}��   �   ,ȧ�a��$�p�S�	T���˙�����Ѿ�efɿcLͿ�ʿt��O��Ia��+���~�U���%�����i���T\�m[��{��vfC�4�B����3Z��ç����b$��S�jQ���ș��|��7ξ��bɿ�HͿ�ʿS��|���^������U�J�%�����f��=Q\�BY��y���gC�J�B�������9Z��   �   �侒�!�b�X�As�������&ƿ��߿�E��� ��B�tC�����t��6ȿ֚��4���<�Z���"���徐���j�<��ؽt4q��J&�b�G�B���bx��f�]ꩾ�8�r��s�?�Hd��(���鎿=,���3��Y����ݏ�0\����f�_�A�e���l^��ڴi�+�(���B�M��l*���s���ؽ#]<������   �   |��&�N�<����C���$ҿ0v���~
�	-�|��׷"��( �.+���[�����ӿ�g������uEO��	�PǾr�z����������,��}7�ȧ����,D]�P�
Ӿ4U�g ��8�6�K�+X��\���X��!M�i]:�Z"�8��j־�ʠ���a�^��H㭽^}A�.7�N�%��ě���$T{��bǾ�   �   �E6��;|��ե��qп2������^&�XH6�RA�LE�h�A�'^7���'���>[���Gѿ+1��@O|�I�5����������[8��l���%(�<ψ����Rs�g������_A��&��5����DԾ'���B?	��9�Ʉ����G
������F׾��������hF����h}��$��<C��`㝼d2�\5Ľǲ:�`Ϟ������   �   �wW��꓿�F���,��<+���B���V�a�d�R�i�F*e���W���C��,�F��k>��������yV�ES�o����_�Z��Ο=�X��0��; T�8�	���_�!%ɽ>�g�N��� '��lV���ٹ�v������4䮾�8��x����S�����ҽl
p���ȼ �T��;p$?�^J� >�TMc��T��OU��   �   ��t����hٿ�����$��A�8=^�8�v��׃�~���L���}w���^��*B�a$�����ؿ�$��U	s��(�p�پ�݁���lX��Y��ؓ�<��< -�<����4���l��3�Խ���-0�{�J�r�[�k0b��]���L�Ww3�T��q�ܽX���ƪ�p����zS<��<���<@����g����)��ݐܾ-�)��   �   �X��_c�k��܍3���T���u��.��X��v���H2���V���u���T���2���$�꿉��������z8�fu�TJ��@A�X�q����l��<�>/=��*=x��<�:4<�nR�������� �����׽�^�Ĉ����1�۽���E��@<-�p,��@��;<��<6Y=d� =���<��û� �����Y��0����:��   �   �K��"����������6�=�f�a�i���I����j���F��Fq������i�����`�sp<��b��f���ѽ��Ë�_�B�����z�����"������̺D=�dW=ԁf=��K=6=̠�< O����5!��[�y��~���/a��<Ib�P%+��ɼ���p<>�=
C==�W=>�H=
 =����j���(�ܹ���j��_E��   �   Bԏ�r�¿����t:��A��;f����������������ו��i���6e��?�6���d������{2����F���� 圾!�&�:ل��߷���=vqd=��y=�f=B�5=!�<�&< �����ü*��$�8��F���<�lt��#׼�c.��!�;@r�<�]'=h�W=�_k=*�U=`�=�~��Lƍ���+����0�{I��   �   QK��M����������V�=�B�a��߂�q���j���E��^p��Ց��������`��o<��a��e��ѽ���u�B���������y�"����� O̺x	=~eW=T�f= �K=X=���<�L�4���5!��[� y������.a��DIb�H%+��ɼ��h�p<��=dC==��W=�H=Z =�����h���(�󸜾(j��^E��   �   �텿���\a�&��=�3���T��u�-����������0��U����u���T�%�2���5�����q���y8��r�H��?���q�`����<P@/=��*=���<�;4<`nR��������$����׽�^�ӈ����/�۽����D��<-��+�����;���<6Z=�� =���< mû�������������+�:��   �   ��t�����eٿ@����$�i�A��9^�V�v��Ճ�H���+���yw���^��'B�J}$�R��]�ؿl"��s�.(��پ>ہ���dX��0��@��<�"�<�/�<���ҁ��l��.�Խ���-0���J�|�[�r0b��]���L�Rw3�M��M�ܽ"���$������P�S<X�<`�<�����g���%'��Z�ܾ��)��   �   �sW�E蓿OC�����2*��9+��B���V�΁d���i��%e���W�N�C�� ,�֗�l:�r��"����uV�\P��j��u�_���N�=��~�0��; �8(��@�_��$ɽ3�j�N���'��tV���ٹ�v������6䮾�8��x���S�����ҽT	p�T�ȼ �T��];?��J��6ｷGc��P��WR��   �   =A6�$6|�Lҥ�kmп������8[&�GD6��A��	E���A�Z7��'���V��ACѿ�-���I|���5�d�������U8��d��l(��������p��񓽈���x_A��&��5���EԾ-���F?	��9�̄����G
������F׾�������XhF�B��v|��6��<:���՝�� 2�N-Ľ��:��ʞ�0����   �   ��R�N���?��fҿp��{
�4)�e����"��$ �R'����0�����ӿc�������?O�"��IǾ�xz��������n�����ly7��Ƨ�~���C]�C�
Ӿ5U�g ��8�:�K�#+X��\���X��!M�h]:�Z"�8��j־|ʠ�l�a����᭽�xA� 0���%�������7K{�~\Ǿ�   �   Ǹ��!�P�X��n������� ƿh�߿�>���� �	?��?�j������Jȿ����ڥ��'�Z�J�"�\�徕����<���ؽ*%q��@&���G�>����w�~f�Gꩾ�8�p��t�?�Kd��(���鎿?,���3��Z����ݏ�/\����f�Y�A�[��yl�h^��l�i�h*������M�Hb*�H�s��ؽ�T<������   �   ����q��$���S�WO��Nƙ��y��"˾��_ɿyEͿ&ʿ���@
���[��m�����U���%����`b��@J\��S�-q���XC�{B�&��(��2Z��ç�r��^$��S�kQ���ș��|��:ξ��bɿ�HͿ�ʿR��y���^������U�?�%�p���f���P\�LX��v��r^C�8|B�\���	��.Z��   �   �f��橾*4�w��̗?��d�k&���掿T)���0��N���ۏ�`Y��υf���A����:fY��
�i�%�����Z�M��]*�8�s�_�ؽ2W<�������4�!�3�X��p������#ƿl�߿B���� ��@��A�*���b�Ή
ȿ����Z���P�Z���"�i��A���$�<��ؽ�,q�C&���G������t��   �   ���P>]�uꝾ�Ӿ.R�vc �ŋ8���K�A&X��\���X��M��X:��U"�V4�nd־tŠ���a����.٭��lA��(�8�%�������M{��^Ǿ�����N� ����@���!ҿ�r���|
�+�`����"��& �[)�s��������ӿ#f��.���;CO����MǾD~z�8��O�����أ�t7������   �   �듽�����YA��"��~���`?Ծ�����;	�6�Ѐ���D
�S���@׾^����󈾕`F�,��1s���y�l'���ɝ�@�1��-Ľ�:�̞�%����B6�08|��ӥ�'oп���&��\&�)F6�A�E�C�A�A\7��'�p�Y���Eѿ�/��7M|���5���������Y8��i�� (�����i��   �    ���F�_�%ɽ��u�N����B"��*Q��Թ�9p�������ޮ�K3��>s����S����ҽ�o�0�ȼ�T���;��>��J��6ｚHc��Q��!S��tW�铿tD��p��*+��:+���B�|�V���d���i�(e��W�T�C��,�T���<���こ�fxV�sR��m��|�_��转�=���pϮ; ��8�   �   |;�<0����u��d���yԽ+�'0�J�J���[�j(b��]��L�p3����ūܽR���ޙ�2��@�S<���<��<�c���g���U'����ܾ)�)�[�t�w���fٿ���z�$�q�A�D;^��v��փ�b���K��|w���^��)B��~$�t��E�ؿ $���s�(���پ)݁���HjX�pC��T��<�(�<�   �   ��*=���<�X4<�HR��������6���3�׽U��~��{��۽����<��b--���� M�;�<Da=�� =���<`QûN�����v�����?�:��텿����a�r����3���T��u��-��n�������1���U��+�u��T�F�2������Q��������z8�^u�ZJ��NA��q� ��ػ�<�A/=�   �   �f=��K=.=̨�<@������.!��[��t��ۢ��l\���?b�R+���ȼб��H�p<J�=TH==��W=��H=� =`~���f��� (�^����i��^E�K�� ���������c�=�n�a��߂�����ej��5F���p��e���A���v�`�hp<��b��f��ҽ��Ë���B���������a�"������̺�= eW=�   �   �q_=ZNJ= �=|��< ��9�������t�J�Ʀn�~�{��q��O�D��l���׺М�<�=d�A=�V=ަ?=�_�<X�r�����kB�LX������T[��'��9ӿ;����+�Z�R�#�}�v��x6��nҳ��<��.ͳ����}-����|�K�Q��y*�~���fѿYߚ�~[Y�RW�}����>�"���GJ����<�oH=�   �   T�J=
:.=hy�<8�<�}M�F�	��W��;��.)���x���n������.�]��`� �n��>�;���<�~%=B=0�1=(��<h�t��n��xB>�ͺ��m�dUW��r��}Ͽ�d�G�(�J�N��Zx��(��b`��������Ƕ���U��������w�&�M�!�'������Ϳ�>��	vU�|��2����:�\�����L�`"�<b�:=�   �   R=�0�<�1�: �ȼ&V�����5ս���^z�03��7�s�����ؽ�d��"x_���ۼ@������<�8=J�=\L�<��~��]���R2��N�����Q�K�(����?ſ3���� �m�C���i�Jއ�/����������������/Ti�*C��u�6Z���Ŀ����!J�5���R��./�����X���<��=�   �   �X�;�w��<�Iϩ�d�����$�߄H���d��6w���}�%x��f���J��'�� �vF���G��������;�Rp<�<\�����R2 ��B����򾲙9�J=��3���E�!�4�2���S�d�t�ŀ��AS��'��Ì���Ԉ�Ku��"T��2����O���s�����h8������\r��*���z���1<�y�<�   �   ���S��0���.���i�3ܑ��˫��q��s�;p�Ҿixξϕ���K��0����Xm��12�����|����J��WO��߻���
�~��=
���~��^Ӿ��"�ek������gѿ}���u�*T:��U���k�4�{�Ԁ�g^|�e�l��U�Y�:����R��Cѿ&b���@j�[�!���ѾK&|���X�v�E��Ђ��(-��   �   ���B-���[�JX��E����������� �$��!����i!	��Iþ�\���_��&�������N��.��T���[e��A�p�R�bJ������[G��Y�������k���C�4���F���R�XqW��S�'�G���5�` ��	�>��P��|b��:#G��s�.{���:Q�m�<�^�0��<lἄ�F��   �   ��$�ثy�+��8�����; 0�6%J�Ӹ^��l���p���l�W�_�F�K�2�1��P�y�'����|��y'��ν<v��2�FpX��ẽ�$'�Ն���`ܾh;"���a� ��<����������$�xC-� �0���-���$�6������X��K����:b��l"�EUܾB<���J&�[ٸ���S���,�to���ɽ�   �   �x��?�������#)�?�Q�y��܍�0����P��2}������sD���͎��{���S�ɧ*�9��¾��Ă��(�zͽWЁ�,�]�����&i���"U��4���[���1��	m���������`�ֿ5��_F��q��� ������,��Xmؿ�۸�㶗��Xn��e2�cG�������fU��"���˕�DH[����YʽO<&��   �   �}��r4�4��mg�����E���w��v�ο 9ڿ�P޿��ڿ�Ͽ��������o-���2i��[5�v������Lw��`�{���&�y���x��·��x�?�u�y��H1�	4��hg���qB��gt����ο@5ڿCM޿��ڿ��Ͽ�����,+��/i��X5�J�j����Hw��^�����x�y�2�x��ȷ��}�6�u��   �   .a����1�1m�zÖ�ו����ֿ��gH�t���"������/��2pؿ2޸�ܸ���[n�2h2��J��6���qiU�%���˕�dC[�&���Qʽ�6&��t���󼾍���)�c�Q��y��ٍ� ���8M���y��Y����A��.ˎ���z���S���*�������B�.(���̽$ρ���]�����[p��*(U��8���   �   l>"�d�a������g�㿯�� �#$��E-�Y�0��-���$���S��)�S��ڥ���<b��n"��Wܾ�=���K&��ٸ���S���,��ro���ɽn�$�V�y�����������0�: J���^�H�k�@�p�^�l�^�_�ƃK�C�1�=M���"����|�yu'�"ν��u�2�\tX�v溽�('�����oeܾ�   �   �^G��[��v��r���l�����4���F���R��sW���S�N�G���5��a �	��⿅Q���c���$G��t�v|���;Q��㽜�^����X��wF������&�:�[�%S��$�������V���� ��$�n� �ź��	����Cþ_X��r_��!�G�����N�l'��U��"ae��F���R��M��J���   �   rk�v���jѿ���/w�(V:�U�|l���{�eՀ��`|���l�C�U���:�����Eѿ
c���Aj�3�!���ѾC'|�	��v�P;���C����,����DI��Ց�m�.���i�ב��ū��k���;	�Ҿ:rξ����F������Qm�z+2�����g����@��@O���߻|����~�h@
�k�~�@bӾG�"��   �   �>��=5���G�T"�¿2���S���t�����T��q��퍒��Ո��u��#T�׵2�n��(��xt��k����h8����G���@r�[)��P z��2<4��<���;��v�x�<��ĩ�������$��|H�$�d��-w���}��x�*�f�a�J��'�� �>���G�D쎼`��;�`p<H�<��������5 ��D�����՛9��   �   V���dAſ����� ���C�>�i�=߇�:��������������������Ti��C� v��Z��Ŀ+���"J�2���R���/������zX�L�<��=�=�C�<���:��ȼNV�����+սX���t��-��2�������ؽS]��fk_�(�ۼ�����	�<h<=��=K�<Р~��`��U2��P�� ��(�K��   �   �s����Ͽ;e��(�:�N��[x�1)��
a������r	��4���$V�������w�3�M��'����{�Ϳ^>���uU�!�������:������L�\)�<V�:=ֵJ=V?.=���<�<�\M�2�	� W��6���#���s���i�����8�]��Y���n�Pa�;���<Ā%=�B=ؿ1=���<��t�aq���D>�Y������VW��   �   o(���ӿ����+�϶R���}�Kv���6���ҳ��<��ͳ�l��D-����|�٠Q�&y*�#���eѿ�ޚ��ZY��V�n
��Z�>����8:J����<�qH=~s_=PJ=��=`��< .�9h��������J�F�n�T�{��q�pO���n��@)׺,��< =ЯA=>�V=��?=<Z�<�r��	��(mB�dY������U[��   �   	s���Ͽ�d�M�(�;�N��Zx�](��`������b��,���1U��������w�>�M�a�'�����Ϳ�=���tU�m������̿:�󨡽��L��+�<�:=Z�J=�?.=��<@	<�\M�4�	�W��6���#���s�� j�����<�]��Y�`�n� b�;L��<�%=rB=��1=t��<0�t��o��JC>�_������UW��   �   ����?ſ˩��O ��C�ړi��݇�w������	������ ������Ri���B��t��X��rĿ䔐�& J�۶��P��H/������jX�<$�<@�=�=�D�< ��:��ȼ>V�����+սf���t��-��2������ؽL]��Dk_���ۼ@���H�<t==d�=<P�<��~��]���R2��N�����9�K��   �   �<���2���D�s �\�2�o�S�҉t����R�����s����ӈ�u�� T���2����?��)r�������e8����Ɯ���n�%��h�y��2<���<���;��v��<��ĩ������$�}H�-�d��-w��}��x�.�f�`�J�ܑ'�� ��=��G�hꎼ ��;�ip<��<H����󎽴1 �gB����'�9��   �   k������fѿ���ut��R:��U���k���{��Ҁ��[|���l�-�U�b�:�7�����Aѿ@`���=j��!� �ѾL!|�*���v�@.��#��X�,����H�����e�.���i�ב��ū��k���;�Ҿ>rξ	����F������Qm�b+2�����ᣓ�:?��5O��{߻򱼞�~�j<
�b�~��]Ӿ�"��   �   �YG��X���������i�w��x�4�b�F���R��nW�~}S���G���5�+^ �G	�b�⿬M���`�� G�Qq��w��`5Q�\�⽄�^����O�(uF�����v&��[�!S��$�������Z���� ��$�o� �ƺ��	����CþPX��A_��!�V�����N� �LG���Ue�Q>�L�R��H������   �   �9"� �a����C�����\��3��$�FA-���0���-���$�#����l忂���衕��6b��i"��Pܾ�8���E&�Ѹ�ĹS�j�,�no�C�ɽ�$� �y�����������0�= J���^�M�k�D�p�a�l�`�_�ǃK�A�1�8M���"��z�|�u'���ͽ��u��2��hX��ݺ�4"'� ����^ܾ�   �   2X����1��m�Ӿ��Y�����ֿ���D��o���
������(���iؿ�ظ�2���OTn�;b2��A������h`U����wÕ��8[�B��~Oʽ�5&��t���󼾇���)�c�Q��y��ٍ����;M���y��\����A��.ˎ���z���S���*���Ҿ��	�z(�i�̽�ˁ��]�[���
d��U�I2���   �   �u��/�14�8eg�����?��iq����ο�1ڿ�I޿6�ڿ�Ͽ5�������X(��&*i��T5��t���LAw��X�`���8qy���x������w���u��x��>1�	4��hg���tB��jt����οB5ڿFM޿��ڿ��Ͽ�����*+���.i��X5�=�;���5Hw��]�h����wy�B�x������u���u��   �   r�����J)�r�Q��y��֍�}��J���v�����N>��)Ȏ�`�z���S�a�*�G	���������(�|�̽�Ɓ�.�]�P���yf���!U��4���[�� �1��	m���������`�ֿ8��`F��q���"������,��Tmؿ�۸�඗��Xn��e2�<G�������eU����oǕ�J;[�޻��Kʽp2&��   �   ��$��y����7�龢���0��J���^��k���p��l��_��~K���1�?I�]�Q����|��n'�\�ͽ�u��2�jeX�'޺��#'������`ܾ`;"�}�a���;����������$�zC-��0���-���$�8������V��I����:b��l"�Uܾ�;���I&��ո���S���,�fho���ɽ�   �   a񴽶!���[��N�������q�x��n� �$�!� �����	���=þ(S���
_��_��N��	��:��2Se��>潓�R�$J�����z[G��Y�������k���F�4���F���R�YqW��S�(�G���5�` ��	�=��P��{b��2#G��s��z���9Q��㽖�^���缌G��lF��   �   p���A��"��O�.�E�i��ґ������e����;��Ҿ�kξ���
A��w���Hm��#2�<������(0�@	O��<߻<豼`�~��<
�X�~��^Ӿ�"�bk������gѿ~���u�*T:��U���k�5�{�Ԁ�g^|�e�l�~�U�Z�:����R��Cѿ#b���@j�P�!�[�Ѿ�%|�����v��1��p��H�,��   �   `��;��v� �<�R�������h�$��uH�\�d��%w�S�}��x��{f���J�'�x �A3����F�TΎ���;(�p<�<���m򎽔1 ��B����򾬙9�J=��3���E�!�4�2���S�f�t�ŀ��@S��&�����Ԉ�Ku��"T��2����O���s�����h8����ٞ���q�%(��p�y��2<x��<�   �   @=�O�<���:��ȼ�	V�0���U#ս�����o�x(�0-�Z���1�ؽgT���[_�x�ۼ�?����<�D=V =�Y�< �~�\��R2��N�����O�K�(����?ſ4���� �l�C���i�Jއ�0����������������/Ti�(C��u�7Z���Ŀ����!J�-���R���/�}����vX�#�<��=�   �   *�J=�A.=H��< <GM���	�X W�r2��2���n���d������v]��P�H�n����;���<b�%=�B=��1=���<`�t��m��<B>�����k�cUW��r��|Ͽ�d�F�(�J�N��Zx��(��c`��������ƶ���U��������w�%�M� �'������Ϳ�>��	vU�x��"�����:�������L��(�<Ȉ:=�   �   DN=p8=<k=0�d<P`ƻԼ�2��l�n����������Hn�p�5��+ۼ z廘�T<$��<&4=h�I=��1=���<�̩�<��?{P��!�������f�1У���ܿ��%4��g^�h����`�������� ������G����5���f���]���3�ُ�1ܿ:��2�e����麾��N��E���៼8м<�6=�   �   �i8=��=|ҹ< �/;hɟ�Ȧ)���y�����*��2q��α�_❽<}��g-�<秼�K�:�s�<��=dV4=Dk#=ݤ<TǪ�����%L�w\������b�����Wٿ���W1�"Z�σ�Y͚�\�������uI��庻����;���R���×Y��q0��>��~ؿ_V����a�V,�R0��8WJ�	���������<�'=�   �   N�<��<`F��r~��(z��l��ɞ��~
�^��V���9�k2�������~��%�P�׻0�r<���<���<(�j<X��P��v�?�,}������uV�mט��ο����(�aN�>�w���������)��:����<�����蹐�lhw�^�M�4�'�z���οK����U�����q���>��[���ʦ���{<�	�<�   �    15:϶�N`�����	�x+3��JX���u��h��ȇ�����^�v��{Y�څ4��!����=e�U�� �ǹ�~#<�{;�=��)����,�-����u ��C�(	����̒���W��<���_��߁��w��*�����]L������
���$`��<�3�^,�����7���A�B�X����᛾�h+�S���0���`��;�4<�   �   j�(��6�������=�,�{�I���;����̾��ھ��߾;۾Nc;������'s}��?����⤽J=-�䬗�PL��l式������ꇾz��+��\w��Ǩ�y�ۿ d	�ۀ&��iD�Pna�Hwz��ׅ����������z��a�u�D�m�&�(s	�ђۿ효�|�v�y?+�8H߾zE�����G�����ݼ��<�Z���   �   ��ʽ9�!���l�C頾]�;:����Q�	����)��M-��*�%; �J��Ӻ����ξ������n��F#��
ͽ��m�(A���2Ƃ�C���5'b��a��b���8R����q����;���'��>��Q��_���c��Z_��{R��B?�v=(����af�>������R�i��
���nMa����,��,��8��ʬi��   �   "3�����黾�Q����aT:�~�U��j���x��}��	y��k��FV�3$;��}�(���!���򆾢v4��+��{��,!P��]x� �νҁ4�� ��1��Vz+���m�<���ȤſK-�J��>��[�,��Q6���9�&�6�;-�qR�f$����k)ƿ�.��u:n�.�+����
ڕ��4��ͽ.v��uM��݉�
��   �   �׊��ZɾR�	�	3���]��T��hj��曣����x꯿������𕿵߃�ը^���3�!z
�pNʾ����rD5�Saέڒ���~��䨽(Q
�� e��D����S�;���y�A���y��/�� �����
�	\���z���C�H���x��׼���=��Ӳz�n%<�����%e��?
��w���<}�9瑽*
�,P4��   �   ؗƾ�A�g>�f9t����� ��w&ǿ�Sٿ��I&�ZW�y�ٿ
�ǿ�����K���3u�#?����;Ǿ�0��	&��̽��%ˍ��	̽.�%�Mȃ�ђƾ�>��b>�Y4t����������"ǿ�Oٿ���b"鿗S���ٿ��ǿʱ��6I���/u�?�E���7Ǿt.���&�݄̽<�~΍��̽2�%��˃��   �   ����;�f�y����������"�����
�@^��
�����E�����s��Y����?���z��'<�D
�H����(e�A
��w���7}�⑽��J4��ӊ�@Uɾ��	��3���]��Q��Cg����������篿K���@݃���^���3�zw
�|Jʾꂋ��@5�L]�oْ���~��訽�T
��e��H���   �   }}+���m��✿��ſ�0�A��r��,�?T6�m�9���6�^-�IT��%�6��{+ƿ�0���<n���+�e�龁ە�64�v�ͽ�v��mM��։�Q��3�Y��仾�J�����O:�E~U�s�j��x�T�}�Zy���k�!BV� ;�~z����������r4��%⽻x��B P��ax��ν�4�������   �   <R�ҁ��������<���'�l�>���Q��_���c��]_�R~R��D?�?(���Rh�@��A���?R����c����Na����*��̳������i��ʽY�!��l��㠾�;ր���M����5�)�tI-�f *�7 ����\����ξ�����~n��A#��ͽ$�m�&=�@��Ȃ�ɶ���+b�;e��Ϲ��   �   `w��ɨ��ۿ�e	���&�lD��pa�&zz�Yم�f������Y {���a���D���&� t	��ۿܛ����v�\@+�HI߾�E����������ݼ�a<��B����(�J,�� ����=���{�����5��_�̾�ھ�߾��ھ>];������'k}�p|?���9ۤ�3-�䠗���K�@p弡������쇾�	�k�+��   �   �
����� ����X�f<���_������x���+��-���M�������
���%`��<��3�D-������������B�����6⛾�h+�%��������Ğ;H84< 
8:���� `��徽x�	�$3��BX��u�d��|Ç�����v�tY�X4�����f/e��@�� iĹ��#<��{;�B��l����,�e���.w �%�C��   �   �ؘ���ο����(��N��w��������+��I����=����������?iw���M���'�����ο&K����U����oq���>�"Z�� æ���{<D�<�]�<�<`粻Dp�dz��c��s��Uy
�������i4�S-��u�Ȑ��*�~���`V׻��r<,��<���<��j<���{���?�&����wwV��   �   ����Xٿ���)1�	#Z��σ�	Κ����6���J��X���e���o���l���ӗY��q0��>��~ؿ'V����a��+��/��$VJ�.���� ����<�'=�n8=@�=h߹<`0;L���J�)�r�y�O����$���k���ȱ��ݝ��}��`-��ۧ�@��:tz�<°=NW4=�j#=�٤< Ϊ�p����'L�^����}�b��   �   �У�8 ݿg� &4�h^�����-a��G������ ���m�����{5��Nf����]�$�3�{���ܿ���?�e���躾�N�3C���ڟ��ռ<6=N=8=�l=�d<�Uƻ�Լ�2�l�,���������In�<�5��-ۼp��x�T<0��<�4=��I=`�1=���<�ө��>���|P��"��P����f��   �   ���Wٿ���^1��!Z�σ�#͚��������H��A���`�����������ƖY�q0�0>��}ؿtU���a�9+��.���TJ�y���<���࣭<ڑ'="o8=��=�߹<�0;0���T�)�~�y�T����$���k��ɱ��ݝ��}�x`-�Xۧ� ��:�z�< �=�W4=�k#=`ܤ<�ɪ������&L�]��G��o�b��   �   Lט�նο���H(��N�h�w�	����ߢ�)��-����;������Ḑ��fw���M��'����ο�I����U����o��w>��V��غ��P�{<��<�_�<H�<�䲻&p�bz��c��|��_y
�������r4�X-��u�Đ���~��� S׻P�r<D��<(��<�j<T��6����?�9}�����suV��   �   ���o�����W��<���_��ށ�xv���(��c���J��<�������"`�<��1�4*��D���ȥ���B�����ߛ�le+�����H�����;8A4<�a8:(�����_��徽t�	�$3��BX���u�%d���Ç�$����v�tY�U4������.e�0?�� �ù��#<�|;X7�����A�,�����6u �\�C��   �   �[w��ƨ�5�ۿHc	��&�{hD�ala��tz�qօ�f������z��a�T�D���&��q	�i�ۿ񘨿V�v�=+��D߾�B����������ݼ�P<�h=���(��+�� ����=���{�����5��f�̾�ھ�߾��ھD];������k}�[|?����ڤ�n1-�`���8�K�pb�C�������釾?��+��   �   7R��~������ ��9��'��>���Q�_���c�%X_�RyR�`@?�d;(���bc�<�����YR���d�Ha�0���$��T��
����i��~ʽ�!�Ƨl��㠾�;ـ���M����9�)�xI-�i *�7 ����\����ξw����~n�}A#��ͽ$�m�p8����Â�ܭ���$b�5`��8���   �   �x+��m��ޜ���ſ�*����i��=�,�`O6�k�9���6���,�>P�p"�7��u&ƿf,��h6n��+�5��|֕�o4�w{ͽ��u�4fM�uԉ���X3�;��仾�J�����O:�H~U�w�j��x�Z�}�^y���k�#BV� ;�|z���������q4�u$�\v���P�*Vx��νD4��������   �   @��ׯ;�u�y�4���� ��;�ῶ�����
��Y�]�F���A�H���Ҟ⿘��� ;��!�z��!<���}��Je��:
�Vo���,}�zޑ���߽sI4�nӊ�'Uɾ��	��3���]��Q��Dg����������篿M���@݃���^���3�qw
�\Jʾ����@5�[��Ւ�p�~�>਽~N
�X�d��A���   �   n�ƾQ<��_>��0t�K���
����ǿdLٿ�促鿲O�*�ٿG�ǿ}���FF���*u��?����2Ǿ�*���
&�M{̽�鍽ƍ�F̽1�%� ȃ���ƾ�>��b>�X4t����������"ǿ�Oٿ���f"鿚S���ٿ��ǿ˱��6I���/u�?�9���7Ǿ(.���&���̽$퍽�ƍ�E̽��%��Ń��   �   �Њ�:Qɾ!�	�Y3���]�aO��~d������j����㯿�ꬿy���ꕿaڃ���^�5�3��s
��Dʾ�~��:5��RὩВ�d�~�3਽�O
�$ e�QD����K�;���y�@���z��0��#�����
�\���{���C�H���y��ռ���=��Ͳz�e%<�o�����%e�Z>
�~s��P/}�6ݑ���߽�E4��   �   �3����߻�HE��v���K:��yU�R�j�f�x���}���x�,�k��<V�Y;�Uv�}�������놾�j4��⽱o��vP�nRx�t�ν��4�u ����Lz+���m�;���ǤſL-�K��@��\�,��Q6���9�'�6�<-�rR�f$����i)ƿ�.��n:n� �+���龳ٕ��4�d�ͽ�v�FeM�xщ���   �   �wʽ�!��l�~ߠ���;qz���I����߿)��D-���)��2 ����������ξ��un��:#�u�̽�m��-�X������\���P&b��a��Q���8R����p����;���'��>� �Q��_���c��Z_��{R��B?�v=(����`f�>������R�Y���󺾉La�����'���� ���i��   �   �v(��$���L�=�і{�*��R0��e�̾��ھD�߾�ھ�V;���������a}�ot?�2�}Ф��!-� �����K�<X�������BꇾL���+��\w��Ǩ�y�ۿ!d	�ۀ&��iD�Pna�Jwz��ׅ����������z��a�u�D�l�&�(s	�ϒۿ뚨�y�v�n?+�H߾'E���������t�ݼ(H<�p1���   �   �::@����_�ݾ��	��3�$;X�Ĵu��_����������I�v��kY��w4���ޛ���e��!�� ���X�#<�g|;�.����� �,������u ��C�'	����̒���W��<���_��߁��w��*�����]L������
���$`��<�3�`,�����6���;�B�;����᛾:h+�⯝�������;�O4<�   �   �f�<�#�<ࣲ��e�Dz��[�����\t
�W�����.��'��k�|�����~���p�ֻ(�r<��<`��<��j<����	����?�	}��{���uV�nט��ο����(�bN�>�w���������)��;����<�����蹐�mhw�^�M�4�'�y���οK����U�{��vq��
>�Z��4�����{<��<�   �   �o8=|�=�< W0;����f�)�j�y�Ĩ������f���ñ�j؝��}�6W-��ʧ����:���<��=�\4=�o#=��<�ª��~���%L�h\����� �b�����Wٿ���W1�"Z�σ�Y͚�\�������uI��亻����<���R���ėY��q0��>��~ؿ_V����a�R,�B0���VJ�K��� ��d��<��'=�   