H   F�`)�Z#@                        ���+BY@                        �{�"TQ@H      6       �        �   �p�����������׽� ��3�d�'�E�5��9?��hB��9?�9�5�P�'��3��� ���׽����
����o�� ����Ž����+Y�gL��1`���M9����*��￰���f>���i���������a��*��x���Y�� b��(���C����i�hg>�d��[�,�����O9�Ab���M���-Y�V��Žn����   �   bd��hg����ŽKK�e��L^%���9�ȠI���S��dW���S���I���9�5^%�C���J�x�Ž�f��{c���򟽾�Ƚ����JW����b����]6�����)X��!f�HA��8;��pe��.�����>9�����?������9��a��q/���qe��9;��A�Xg�6Y������N_6�j������LW�����Ƚ.����   �    ����ӽN+ �����9�k{W���q��`������`������`����q�O{W���9����+ ��ӽ#���҂����Խ����R��՝��쾭�-�~�w�}��R��N\�n!2�0&Y����k���xN��\��ZE������N��ԗ������ 'Y�*"2��\�{�� ��+�w���-�ޗ�ם��	R�R��k�Խ����   �   8��@��e3�cx[�S0���6������鹾�zþ��ƾ�zþ�鹾����6��@0��1x[��d3���j��
޽���W��I�J�L���۾�� ���d��7��.�Ͽx��^H$���F�t�k�
a���v���o���R��p���v��da��2�k���F�I$���B�Ͽq8��$�d�Ϫ ��۾dM���J�������9޽�   �   �?%���L�������>%��y�۾�g�����Q��� �N��~��}g��f�۾&%��x��������L�x?%�8���U�~�xmB������ƾc	�"�L�N����y��� �p�x�0���O�J~m�����%x��՜��Ex��ڤ���~m�\�O��0���!z��'�����L�v
�5�ƾ9���oB�5��V�Ț��   �   �Ka��l��􎵾���S>�{�$P1���@�>K��vN�9K���@�P1�{�E>����Ҏ���l���Ka�:�5����΀���;��+y�9�����EX1���s�9��;Ͽ7���l4��H2�^�I���]��j�&�o�D�j��]���I�xI2��4�4����<Ͽ�r�s�yY1���������-y���;�с������5��   �   �2���žS�����f=��\���w�a���C���E�A���\�����w��\�T=�|���R��V�ž�2��Nl��8@�IO.�ڎ8�db�o���*վ�.�٫L��������6ؿ�/���0!(��)7��A���D��A��)7��!(�T��Z0�ؿå������L��/�q,վ:p���eb��8�,P.�>9@��l��   �   LBʾ�����*���T�h��Wڔ��/��$���娾����ᨾ�����/��Mڔ�^���T���*����Bʾ���,�k��D�M?:��lO�����6��3���v&�eO]�9S������i�ӿ����j!	�H���S�����S�z���!	�7����ӿ3����S���P]��w&�����7�����nO�X@:�wD���k�Q����   �   %x�..��1`�oy��v����=¿/�ٿ��y������u�����%�ٿ�=¿h���by���1`��-.�
x�N�¾�����a�*�A�V�A�a������¾�u��*.�x-`��v��y}��O:¿��ٿ��}������������ٿ�:¿~��mw���.`��+.�fv�!�¾�����a�|�A��A�U�a�����¾�   �   |y&�5S]��U��Z�����ӿL���t#	�v��V���V�r��n#	�=�����ӿI����U��S]�^y&�;!��>9��/��nO�?:��D���k�>���>ʾ
����*���T����kה��,��ă��m���������������,���ה�C��x�T���*����G?ʾ?��� �k�D��?:��nO�z���9��v!���   �   �L����{���9ؿ�1���p#(�,,7�`A��D�\A�&,7�h#(����1�%ؿi�������L�81��-վ�p���eb�(�8�N.��5@��l��/����žCM�����.�<�\�s�w�����[���_�t��������w��\���<����{N���ž0��_l�7@�O.��8��fb�7q��,.վV1��   �   A�s�Q���Y>ϿC���:6�K2���I�v�]��j��o���j�p�]���I�K2�.6�-���C>Ͽ=����s��Z1�N��I����-y�F�;�2������5��Fa�di�����4��;�Rw��K1��@���J�rN���J�\�@�ZL1��w��;�#��a���,j���Ga��5��������;�{.y���������Z1��   �   跌��{���"���F�0��O��m�����y��b����y�����ڀm��O�8�0����"{��Է��n�L����ƾN����nB��}�xT�җ��;%���L��������t ����۾pa��<���������l���a����۾!��5���p����L��<%����2U��~�	oB�������ƾ ���L��   �   �8�� �Ͽ����I$���F���k�Nb��!x��gq��8T��bq��x��Fb����k���F��I$������Ͽ�8����d�� ��۾UM��w�J����p���޽o{󽊮��`3��r[�-���2��� ��A幾!vþ�ƾCvþ�幾� ��E3��|-���s[�la3�f���|�8޽������J��M��V�۾<� ���d��   �   � ��ض�:]��"2��'Y�����{����O�����nF��}���O��r��������'Y��"2�,]���࿣ ��D�w���-���쾾֝�	R�^����Խ󀶽�����ӽL( ������9��vW���q��]�����]��-��^��/�q�NwW�R�9�>��) ��ӽD���
�����Խ˥�t	R��֝����-�l�w��   �   Y��Cg��A��9;��qe��/������9�������?�������9������/���qe��9;��A�&g��X�������^6�������KW�*����Ƚ� b���d����Ž�G�@���[%��9��I���S�bW� �S�b�I�m�9�l\%�̦��H���Ž�e��c��󟽤�Ƚ���LW��������_6������   �   �+������g>�|�i�	�����a��E��w���A���a��珥����f�i��f>�����n+��y��@N9�a��
M���,Y�r��!ŽR����o��؍��X���=�׽�� �d3�)�'��5��9?��hB��9?�b�5���'��3�� �Q�׽h���掗��p��:����Ž���-Y�<M��Xa��cN9�����   �   aX��Uf�ZA��8;��pe��.������8��m���{>��i����8������.���pe��8;�JA�8f�HX�����-^6���������JW�����Ƚ���a��vd����Ž{G�>���[%��9��I���S�bW�%�S�g�I�p�9�j\%�̦��Hｾ�Ž�e���b������Ƚ��%KW�������P^6�*����   �   ]����\�!2��%Y�����Ζ���M��g߶�HD��c߶��M��Ŗ�������%Y�!2�\����E��>�w���-����w՝�jR�P����Խ#�������u�ӽ6( �}����9��vW���q��]�����]��4��^��6�q�RwW�N�9�4���( ���ӽ����8�����Խ����R��՝���쾪�-�f�w��   �   7����Ͽ���G$��F�(�k�)`���u���n��\Q���n���u��!`���k���F��G$����q�Ͽ�6����d�� �m�۾�K��2�J�����꽮޽�z�R��a`3��r[�-���2��� ��H幾*vþ	�ƾKvþ�幾� ��G3��{-���s[�Oa3�2��K|�޽��꽐����J��K����۾?� ��d��   �   �����x��;�T�0�:�O�N|m�f����v��J����v��a���@|m�,�O�H�0���"x�������L�����ƾ8����kB�/|�]S�'��t;%���L��������r ����۾va��A���������q���a����۾!��0���b����L�{<%���T��|�UlB�v���ɛƾ��5�L��   �   F�s��D:Ͽ>���*3�dG2�d�I�T�]�^�j�>�o�Z�j�L�]�Z�I�ZG2� 3�(���-:Ͽ��"�s��V1�8���ڂ��j)y�V�;�M~����%�5�/Fa�Bi��m���+��;�Sw��K1��@���J�rN���J�b�@�]L1��w��;���O���j���Ga�M�5�������;��)y����w���W1��   �    �L����M���ؿ�.�^��R(��'7�bA���D�^A��'7�H(�T���.�ؿ;������ߩL��-��(վ�m��Vab�/�8�2L.��4@�l�Z/��؀ž2M�����,�<�\�w�w�����_���c�w���������w��\���<����lN���žG0���l��5@�*M.���8��ab��m��)վ�-��   �   �t&��L]��Q��k����~ӿ�����	�T���Q�����Q�P���	������~ӿ[����Q���L]��t&�Y��r4������iO�=<:�D�j�k�箘��=ʾ�����*���T����mה��,��ǃ��q���������������,���ה�C��v�T���*����?ʾ诘��k�CD�1=:�wjO�:���4������   �   �s�\(.�`*`��t��{���7¿W�ٿ6쿵���+�������/�M�ٿy7¿{���t��F*`�@(.��s�$�¾y���{a�9�A���A�z}a� ����¾�u��*.�s-`��v��z}��Q:¿��ٿ�쿂��� ����������ٿ�:¿~��mw���.`��+.�Pv���¾��a���A� �A�y|a����_�¾�   �   ;ʾ���I�*�*�T�����Ԕ��)���������2�����������)���Ԕ�����T�3�*�����:ʾ׬����k��D��;:�njO����6�����~v&�\O]�7S������k�ӿ����l!	�J���S�����S�|���!	�9����ӿ3����S���P]��w&����e7������kO��<:�dD�a�k�����   �   -���}ž�H��$����<��\���w�󤆿����}�������w��\���<����H��j}ž�,���l��2@�K.��8�'bb�}n���*վ�.�̫L��������6ؿ�/���2!(��)7��A���D��A��)7��!(�T��Z0�ؿ¥������L��/�,վ�o���cb�?�8��K.�&3@�0l��   �   �Ba��f���������P8�t�@H1���@�<�J��mN�7�J���@�8H1�t�B8����܆���f��CBa�m�5���m}�G�;�:*y�Ń��� ��4X1���s�8��;Ͽ6���l4��H2�`�I���]��j�*�o�F�j��]���I�xI2��4�4����<Ͽ�k�s�iY1����)���7,y���;�q~������5��   �   �8%���L�6��A���i��,�۾�[��1�����&�����+���[���۾S��'�����~�L�|8%���R��{��kB�����J�ƾL	��L�M����y��� �p�z�0���O�J~m�����&x��ל��Ex��ڤ���~m�\�O��0���!z��%���|�L�`
��ƾ����XmB��|��R�����   �   Yw�ʫ��\3�Cn[�?*���/������Ṿ�qþd�ƾ�qþṾ����~/��-*��n[��\3�|���v�޽���|���J��K��ߩ۾�� ���d��7��0�Ͽz��^H$���F�v�k�
a���v���o���R��p���v��ea��4�k���F�I$���D�Ͽq8���d��� ���۾M��ՁJ����K���޽�   �   �����ӽ$& ����D�9��rW��q�V[��Z��[��V��N[���q��rW� �9�����% ���ӽ����~���Խƣ�R�e՝�Ε쾥�-�~�w�}��S��L\�n!2�0&Y����k���xN��\��[E������N��՗������ 'Y�*"2��\�}�࿁ ��)�w���-�����֝� 	R� ����Խ\���   �   La��lc����Ž6E�ˤ�$Z%��9���I�l�S�__W�h�S���I�ݞ9�Z%�����D�~�Ž�b��b`�����Ƚ��-JW����R����]6�����(X��"f�HA��8;��pe��.�����=9�����?������9��a��q/���qe��9;��A�Yg�5Y������L_6�Y������5LW�z����Ƚ���   �   0Q��H��q���ӽ����{t�Ns$�%�2�̏;���>�J?;�� 2�L�#�X��[{����ѽ4����*��@4��$/��ﾽj�
�T�ί��0,����5�l���|�����꿚��r�:���d�\��㢡�[���)k������n������С��)���e�0[;��d�C�뿏���U��<r6�`t��ު��ЛU��L��>��|Y���   �   d�������q��O�+d"�BJ6��E�^�O�/S�؊O��PE��t5��i!�`�
����w����Ơ������h��ʻ½S$�9R�|���4t�R�2�?�~��������~���7���`�F�����A�� ��H������s����>���O���Aa�88����ٳ�����`�3�2������S�l�kŽ����   �   �F����Ͻ����E�.�6���S�Աm�l��)���$���`\��ᰀ���l��R�^�5���� G��+�ͽ���f����ν���dM��l�����j*��s�����Ĩܿ���>�.���T�Bp~�~0���a��C������)���iL���+��(�~�5U��?/��0�[ݿL�����s�B!+����YJ���N���x�нBѲ��   �   ���VV0���W�U�������&����������$þPſ��A��E���T���4L��ldV�d�.�|��F���׽�0����h�E����(1׾Ă��p`��X���G̿�]�Po!�b>C�B=g�*���� ������Fq��\���J���_��\g� EC���!�B���̿���� a����ؾ�ڑ��G�j�^U潈�ٽ�   �   vZ"��pI�` |��/������XؾSX�U�$�m���
�@����l׾/��wN���iz��H�d"!�Z���������=��ԅ��¾A@�
�H�"0��_D���,�$���-���K��i����M����u��4U��O����h���K���-����\C�u���i��s7I�I���KþDl���?�d�����

��   �   �}]�6�������Rݾi�'��%u.�8�=���G���J�8SG��Z=���-��[�F��T7ܾ����XK���/\�%e1�%��|����7���s�����:��C.��o�7��p�˿�������v/�.qF�X�Y��uf��j�xf��Y���E�P�.��{�ŗ����˿=3��,�o��M.������{����t�Wg8�S������{2��   �   ����ET¾,S���r�:�T�X���s�,����>��_�����82����r�B�W�CE9�L��\.��n������w�f���;�\*�g4��]��r��k/Ѿ]��z I��ׅ�yޫ�q�Կ�����i�А%��94���=��
A��=���3� %����l���mEԿk���}���I����ZѾm����;^��5��+��<�l
h��   �   ��ƾ����(��iQ�Z(|�4�������ٶ��✻�����^���F��������: {�0�P�&h'��M�r/ƾi���!�f���?��K6�%2K�*����������^�#��Y�Q��(pcп�?���Z��\��pH�����"����Y�b�Ͽ�`������6Y�t_#�4��T孾����mK�U�6��l@�	�g�����   �   �B�%W+�x�\�V������a��k�ֿ��迂�󿉽���������տ�����[���ӈ���[�g�*��� ��'��Q<����\�7�=���=�5]�+w�����@��S+�H�\�|S�������]���|ֿ��迗�󿥹�����翽�տۢ��7Y���ш���[� �*��� �h%��;����\���=�-�=�58]��y�������   �   =�#�ϯY�����𭿮fп-C���~������J����$�8���[��Ͽ�b������^9Y�8a#���ﾽ歾�����mK��6�Qj@��g������ƾ���(�7eQ�E#|�S���w�������w���E����Z���C��3��J��{�ωP��e'��K��,ƾ�����f���?��L6�84K������������   �   �#I��م��૿i�Կ�����k��%�<4�x�=�<A�l�=�ʻ3��%�:������GԿ��������I�K��R\Ѿ$���<^��5��+���<��h������O¾xM��Vo��:���X���s�d���;���|������/��.�r�.�W��A9����*���j��r�����f�k�;��[*�m�4���]��t���2Ѿ����   �   #�o�(9����˿ �����y/��sF��Y�hxf���j� f�DY���E���.�$}������˿c4��Ժo��N.�����B|����t��f8����[��.x2��x]����C����Mݾ1�t��q.���=��G��J��NG��V=�/�-�|X��}��2ܾE����H��g,\��b1�&�����J�7���s��	��6>���.��   �   �1��YF��</꿘����-���K�i���т��lw���V������څh��K���-�����D��u��:j��X8I�ѥ�Lþ\l��,?� ����� 
��V"�{kI���{��+��3��bSؾNR�jR�� ��i�M�
�<�Q~�Xg׾+��CK���dz�H��!���������k�=�օ�c�¾�A�l�H��   �   �Y��|I̿_��p!�@C�L?g�b���"������r������^���`���g��EC�2�!������̿����\!a�9��ؾ�ڑ�G�W�4R�0�ٽ����Q0�2�W���殕��"��0���,��Y þ����u=���������|I��`V���.�������׽80但�� �E�Y��Y3׾^���r`��   �   ����A�ܿ���Z�.��T��q~��1��c��a���������1M��n,����~��5U�@/�"1�K[ݿp�����s�>!+����J��L�N����н!β��B����Ͻ�������6���S���m����V���T����Y��Z����l�'�R�5����C��<�ͽ�������4�ν����M�n����Fl*�rs��   �   � ����n�~�7���`���� ��������֨��[������?��P���Aa�88�����翤��������3����7����S�(k��Ž������좽�������3��a"��G6�d�E���O�k,S�M�O�uNE��r5�*h!���
�P��ۮ���Š������h����½.%��:R������u�k�2���~��   �   ±�C������:�N�d����$�������Bk������n��R��VС�b)����e��Z;�,d�����������zq6�>s�������U��K��=��bX��:P��FG�����>�ӽ���2t�s$���2���;���>�^?;�� 2���#�����{��_�ѽ����h+��-5��<0��]�I �3T�����P-��O�5�慁��   �   ������~���7���`�-���������������B������/>��]O���@a�:78�\����<��@�3������.�S��j��Ž��������뢽�������.��a"��G6�j�E���O�q,S�S�O�wNE��r5�)h!���
�H�载����Š�J���Dh����½�$��9R�荠��t򾮹2���~��   �   a�����ܿh����.��T�ro~��/��,a��T���������JK���*��j�~��3U��>/�0��Yݿ�����s��+�����H����N�����нSͲ�)B����Ͻ�������6���S���m����[���Z����Y��`����l�,�R�5�����B����ͽc��٤���ν���[M��l������j*�ws��   �    X��G̿|]��n!��=C�<g�P������Q����o�������^��Pg�ZCC�8�!�*���̿�����a�C�8ؾ�ؑ��G���\P��ٽf�����Q0��W���宕��"��4���6��_ þ����}=���������|I�� `V���.����9����׽l.�����E�����0׾k��p`��   �   x/��qC���+�P����-��K��i������mt���S��㼀�d�h�t�K�ڶ-�:���@�s���g��5I�}��ZIþIj��{ ?�e��x��o
�V"�8kI���{��+��/��dSؾSR�nR�� ��i�R�
�B�Z~�\g׾ +��?K���dz��H�z!�2�����ۺ���=��Ӆ�B�¾�?��H��   �   @�o��5����˿������du/�@oF�
�Y��rf�2�j��f�JY�H�E�B�.�"z�Ɣ���˿.1���o�K.������x����t��c8�ي�*��ow2�Ex]����.����Mݾ.�u��q.���=� �G�	�J��NG��V=�4�-�~X��}��2ܾ7����H���+\�Db1����Ȯ�l�7��s�h��79��.��   �   �I��օ��ܫ�c�Կ���Bh���%��74���=�>A��~=�F�3���$��������yBԿ�w����I����LWѾ�����7^��5��+�_�<��h�j����O¾eM��Qo��:���X���s�g��<���|������/��5�r�0�W��A9�����)���j��=�����f�A�;��Y*��}4��]��q���-Ѿ��   �   ��#���Y����쭿�`п�<�>�l��D��@F��� ����gU�'�Ͽ�]������"3Y��\#�ȍ�⭾����RiK�H�6��h@�g����N�ƾ���(�2eQ�B#|�S���x�������{���I����Z���C��5��K��{�ωP�}e'��K�z,ƾE����f�5�?��I6��/K�֐��(������   �   l>��Q+�=�\��Q��m����Z���yֿG�����Ƶ�� �����*�տ����KV��sψ���[���*�b� �~!��8���\�R�=���=�h3]��v������@��S+�B�\�zS�������]���|ֿă迚�󿫹��������տݢ��9Y���ш���[��*��� �%���:��M�\��=�T�=�n2]�ou�������   �   ��ƾ���l(��aQ�|�ᓒ�����t���2���㌾�eW��O@����n��	{���P��a'��H�M(ƾ@�����f���?��H6��/K�u�������n��L�#��Y�M��&mcп�?���\��^��rH�����"����
Y�e�Ͽ�`������6Y�d_#�����䭾j���rkK� �6��g@�Ĝg�����   �   +���xL¾I���l�j
:�~�X���s��|��?9���y������,�� �r�w�W��=9���K$��Mf�����f���;��W*��|4�?�]�@r��/ѾE��m I��ׅ�wޫ�q�Կ�����i�А%��94���=��
A��=���3� %����o���oEԿm���|���I� ���ZѾݮ��:^��5��+��<��h��   �   �t]�#��Ρ��,Iݾ|�>��_m.���=�ÈG���J�_JG�[R=�!�-��T�az��-ܾ٭��JE���&\�w^1�^��*����7�U�s����:��2.���o�7��p�˿�������v/�0qF�\�Y��uf��j�zf��Y���E�T�.��{�ȗ����˿=3��(�o�xM.�d���%{��I�t�e8����.��Ju2��   �   �S"��gI���{��(��8���Nؾ�L�iO���pf���
�
��\x��a׾l&��HG��]^z��H��!�G��������.�=�
ԅ�¾*@���H�!0��_D���,�$���-���K��i����N����u��5U��Q����h���K���-����aC�u���i��l7I�3���Kþ�k��?�ۺ�����
��   �   ��P�=N0���W�X����������������þ[���9��x���f���>F���ZV�Y�.�&����콦�׽A+���.�E�����0׾����p`��X���G̿�]�Ro!�b>C�B=g�)���� ������Gq��[���I���_��\g�EC���!�B���̿���� a���oؾFڑ�x
G���P�@�ٽ�   �   X@����Ͻw������6��S�+�m�-	�����������V�������l���R��z5�d���<���ͽ}������y�ν����M�~l��ʹ��j*��s�����èܿ���@�.���T�Dp~�~0���a��C������*���iL���+��*�~�5U��?/��0�	[ݿM�����s�:!+����J��@�N����н�̲��   �   V���ꢽ����l���
�`"��E6��E�%�O��)S���O��KE�,p5��e!���
���轓���à�����9f��"�½�#��8R�^���%t�L�2�=�~��������~���7���`�F�����A�� ��G������s����>���O���Aa�
88�� ��ڳ�����[�3� �󾥀����S�xk��Ž�����   �   �倽Rh������Ƚ�%�R�
�0���h)���1��4�V:1��;(�gb����_���ýb����ᆽͷx��·�L����Z��G��̙��H,�̤u��Ȩ��߿�V�v�0���W��2���̖�/����(��$���G.��E������Ũ����X��2�VY��������w�ܓ-�
f뾇���HK���{w���l���   �   �?��q��\���:޽�����-�%�;�V5E� 3H�̋D�ٝ:��S+���(����ٽjx���۔���������G��\���4F��ȗ�~�uN)���q��+��y�ۿd,��.�&�S�~a}������ѥ����=d��I��Yݥ�Iғ�&~�N�T��/���D6ݿ�j��8�s���*��羄����7I�@ �d���W���   �   h����}ĽZ�<��-�h0I���a�d*u�ٲ������zP��ϼs���_��F��+����vr�
����\�����ž��^?�peA�) ��]۾�t!�Ҁf�����k�ѿ�����%�l?I��7o�����2=�������m���`�� ��E���P{o�<�I��&����)ӿ����'h�,�"�4nݾ٫��5D�����iŽ*����   �   k1�B���p'�jM��Xu�VT��1؟�桭�x`��9���䵾����X���
����xr��DJ�ݸ$��$��lݽu]ɽ�oսAW��:�$7����˾�A��T�듒��@¿)��B{��9�:=Z���z�Z����2������\����>���Rz���Y�H"9�N�������ÿ@L��&V��J��v;����	=������ٽ|�ͽ�   �   ��$a?��o�%�����8�;�Z�D����*��B����*Y��
�徸�˾�>��瑾�}l���<�y��n� �Ԃ����	�U23��%}�*R�����]v>�1=��cI����޿��	�<[%�2SA��\���r��
������>�����q��$[���@���$�~�	��߿���������A?���Ԝ��St��R5��
�����$���   �   KqR��&��P�T�Ҿ�<��Tg��%��m4��=��@�@2=��3���$��@�s���zsо&��	���d�O�|/'�}������C-�N�f�C����x��/%�Ìc��g���!¿��<���&��O<���M�\�Y���]�*
Y�LM��G;�D	&�N�2k�Q���r`����c�u�%��R꾂أ��sh��.��j����d)��   �   �D��7̸�W1�2���1��+N���g�,!|��n�����5��{�`�f���L�G�/�L����~��쌾�GZ�Te1�W� ��*�!�Q����dmƾ��	?�ۄ~�Ϝ��.�ʿ�������0\+�n14��7� �3�^�*�������R���ɿ��D�}�H�>�����ƾZ����R���+�22"�U3�rf\��   �   ���4�������@G�p�V����ќ��6������^���3���o��ٛ�ޗ��J,n��E�$������M�������iZ��y5�qe,��`@���s���L��}q���N��K��׮����ƿ��� �Ч�
����j�.�
� �b��s[ſٲ��J����N����N@�,���"�s���@��-�py6���[������   �   n���[�"�;�Q�����`1��
m����̿�ݿs远��Y���ܿ�8˿�!��H��&ԁ��P���!��k��<.���ǆ�9IQ���3�'�3���Q��;���񵾩���4�"�?�Q�:����.���i���̿p�ݿSo������翻�ܿ�5˿	����Pҁ��P�c�!��h��2,��\Ɔ�AHQ���3���3���Q�
>��l����   �   8t�U�N��M��������ƿ�濶� �ة� ��̷�d��
��	 �5���]ſѴ��ס��N�f���B㾃���`�s���@�r-��v6���[�����������A��o<G�:p������Μ��3��ן��][���0���l��n֛�����Y(n���E�����������̘��}Z��x5�f,��b@�h�s����G���   �   �?���~�/����ʿO��������n^+��34�L7�R�3�X�*�^��f���T���ɿ�����}���>����ƾ���R�Ļ+�>0"�(3��a\�lA���Ǹ��+�����1�F'N���g��|��k��N�����)�z��f�͟L��/������n���錾EZ��c1� � ��*�u�Q����npƾ���   �   ԏc��i��$¿�����&� R<�n�M��Y���]��Y�lM��I;��
&�z�m������a��+�c���%��S�'٣�th�z�.�i�9��m`)�NlR��#��!�/�Ҿ�6���c�.�%�vi4�1�=���@�.=��3�m�$��=�V���Yoо��������O�l-'��������D-���f�f����{�82%��   �   �>��EK���޿T�	��\%�&UA��\�J�r���쨃����q�`&[�`�@���$�L�	��߿蟮�@����B?�l��S����t�ZR5��	�����Y����<\?�Õo�\�������;2U� ����'��?����pS�����@�˾�:��䑾�xl�2�<��� � �Ł��,�	��33�R(}�VT��L���x>��   �   H���CB¿9���|� 9�?Z���z�����%4��D��������?��:Tz���Y�#9�������Lÿ�L���V��J��v;馊�q=������ٽP�ͽ�+�ĭ��l'�#M�NRu��P��Cԟ�����\���4���ൾ����У���򌾮sr�d@J���$��"�^iݽ�[ɽJoս�W���:�y8����˾8C�'�T��   �   ������ѿ�����%��@I��9o�r���6>�������n���a�����џ��|o���I�<�&����jӿ1���(h�)�"�
nݾ����d4D�����gŽ,�������(yĽXT8��{-��+I���a�)%u�*���N����M���s�2�_�[�F��+�Q���n�@����Z��$����� @��fA�`���^۾v!���f��   �   �,����ۿ-��.��S��b}�����ҥ�[���d������ݥ�|ғ�Z~�`�T��/���6ݿ�j��ӵs���*�z�������6I�d����V���=��jn��D���6޽������ -���;��2E�x0H�c�D���:��Q+���Ȓ���ٽ�v���ڔ�����μ��nH��0��66F��ɗ��征O)�@�q��   �   mɨ�6߿W���0� �W�3��͖�[����(��%���/.������������H�X�`2��X�p��l��
�w�%�-��d뾿���$K���-v���k���䀽�g�����@Ƚ�$��
�����h)�u�1��4�l:1��;(��b���������ý����↽��x��χ������[�'�G�}͙�#��,���u��   �   �+����ۿx,��.��S�Ra}�S����ѥ�U���c������ܥ��ѓ�~�d�T��/��35ݿj��Ѵs���*����\��� 6I�������U��A=��<n��*���6޽������ -���;��2E�}0H�f�D���:��Q+���ʒ�u�ٽ�v��fڔ�f���f����G�����j5F�?ɗ��~��N)�D�q��   �   |���1�ѿ���P�%��>I�67o�����}<������l���_����T����yo���I�ڣ&����� ӿ䒟�&h���"�3lݾ`����2D����LfŽZ���"����xĽ'T8��{-��+I���a�2%u�-���R����M���s�:�_�b�F��+�J��vn�����PZ��`��ٽ��"?�heA�2 ��]۾�t!���f��   �   �����?¿S���z��9�<Z��z�a����1����������=��pPz���Y�� 9��������ÿ�J��V�I�Zt;=���G=�F����ٽ$�ͽ7+⽉��|l'�M�?Ru��P��Dԟ�����$\���4���ൾ����֣���򌾱sr�^@J���$�n"��hݽ�Zɽ�mս�V���:��6��Y�˾_A���T��   �   �<���H����޿,�	�2Z%��QA��\���r�z	��6���߿��B�q�L"[��@��$��	�?߿������y??�3��Q����p��O5�������������[?���o�O���}���;3U�&����'��?����|S�����E�˾�:��䑾�xl���<����`� ������	�D13�n$}�`Q����u>��   �   0�c��f��A ¿������&� N<���M���Y�l�]��Y���L��E;�V&���Vh�����y^��z�c��%�O��գ��oh���.�6g����_)��kR�v#��
� �Ҿ�6���c�.�%�vi4�6�=���@� .=��3�r�$��=�Y���Uoо���������O��,'�n�����+B-���f�4���8w��.%��   �   L?��~�B���6�ʿ��򿦄�ҧ�4Z+�</4��7�Э3�&*������HO�+�ɿ���g�}�C�>�<�&�ƾ�����R��+�e."��3�a\�/A���Ǹ��+�����1�D'N���g��|��k��R�����2�z��f�ҟL��/������T���錾iDZ��b1�X� �E�*�8�Q�֢���kƾO��   �   �o�f�N�J��ଥ�*�ƿ6�*� ����}����X�,�
�3 ���_Xſ0������N����<��=�s���@��-�9u6���[�S���`��ɴ��7��g<G�6p������Μ��3��ڟ��a[���0���l��q֛�����](n���E��������{���|���p|Z�<w5�rc,�v^@�Q�s�W��گ��   �   p����"�V�Q�d���P,��;g���|̿�ݿ�k�7�����ܿ�2˿���B���ρ��P�7�!��c��x(���Æ��CQ���3���3��Q�,;����z���&�"�7�Q�8����.���i���̿r�ݿWo���������ܿ�5˿����Rҁ��P�\�!��h���+���ņ��FQ�m�3��3��Q�:���ﵾ�   �   ���������09G�C�o�>����˜��0������!X���-���i��uӛ�Ӓ���#n���E�E��������������zxZ��t5�3b,�f^@�~�s������jq���N��K��Ԯ����ƿ
��� �ҧ�����l�0�
� �f��u[ſ۲��I����N����@�����s���@�l-��t6���[������   �   ?���ĸ��'�+����0�^#N��g��|�(i���|�������z� ~f�S�L��/�U��L����挾�?Z��_1�[� �Z�*�[�Q�|���
mƾl��?�҄~�˜��+�ʿ�������2\+�p14��7�$�3�^�*�������R� �ɿ��B�}�>�>�p�:�ƾ���)�R���+�6."��3�Z^\��   �   �hR�!���驾��Ҿa1���`���%��e4��=�W�@��)=��3���$�0:�F���:jо���K�����O�)'����g��{A-���f�����yx��/%���c��g���!¿��:���&��O<���M�^�Y� �]�,
Y�NM��G;�F	&�P�5k�S���s`����c�g�%�UR�أ�krh���.�]g�&���])��   �   �yX?�ݐo�A���������;P�j{���$��<�r��`M��<��#�˾t6��@����rl��<����� ��{��R�	��03��$}��Q�����Qv>�.=��`I����޿��	�:[%�0SA��\���r��
������?�����q��$[���@���$�~�	��߿���������A?�֜�����Ns�BQ5�Q�����B���   �   (�'��:i'��M�Mu��M���П�Ǚ���W��^0��rܵ�{���🞾v�mr�";J�0�$���Lcݽ�Vɽ�jս�U��:��6����˾�A�	�T�ꓒ��@¿)��B{��9�:=Z���z�[����2�� ���]����>���Rz���Y�H"9�P�������ÿ@L��$V��J�tv;�����=�����ٽt�ͽ�   �   b���vĽ?P�6��x-�/(I�X�a�e u���������?K��ܲs�^�_���F��
+����h�P����V��p
������<>��dA������\۾�t!�πf�����k�ѿ�����%�l?I��7o�����2=�������m���`��!��E���R{o�<�I��&����+ӿ����'h�%�"�nݾ����X4D�o���fŽ�����   �   �<��Gm������4޽B�����,�h�;�Z0E��-H�ԆD�"�:��O+���ʐ��ٽ�s���ה�-���x����E��ʁ��4F��ȗ�~�qN)���q��+��x�ۿd,��.�&�S�~a}������ѥ����<d��H��Yݥ�Jғ�(~�P�T��/���D6ݿ�j��8�s���*���g���|7I�������U���   �   P�h��*|���!k��;�ڽ�G�����F�+�"�.D%��!�w��p�\/��u�ӽ����a��!�l�X%Y��in����`��5�8r���վ�}�+8a�?��bJͿ���X"�N�D�@Ii�������������T��v8��LX��nNj�,�E�t�#�t<��VϿ����v�c����iؾ-'��y:����r���~��   �   ��{�B��������ʽ<�8�����L,�x�4��b7���3�l*���
��콪�ý����)g���cl�MX{��z���f�0?4�X���z�Ѿ����]�&���,ʿ������UA�	e��V���������I��i���?��䍄�D�e��iB�  !�T(��̿�7���(`����$վ�<��S�8�0���e��o���   �   �g�������ٽ|�6���8�_gO��a��<l���o��k�K_���L��O5�Tp��(���ѽ`:��ԫ�������7��`����/�zT����Ⱦ����US�����B���������>8���X�2�y��݊�ꀔ��ߗ�-^�����oy��GY�f�8��^��D��ܔ¿vU�i����˾𾇾�&4�W���4䳽�2���   �   ~�ν������o<��a�YՂ�璾<���s��r���dǦ��@��3��T׀��=]��8�Jg��^�>�ƽsM��������0�)�ףz��o��ӱ��+C�P���T²���vR�>�)���F��c��+{�^���.���(~���nz��vb���F�0�)�x���~���������D�F
��ϼ���~�:{-��F��n�ƽ�����   �   43���/�N@\�*���&Ȣ�D$��ߚԾ�
羧��e��7��r徠yҾ���>@���B����W�9u+��K	���ݽ���#�>g�b���dL���.�>q�CU���nͿ�	��v.��61�̣H�<5\��@i���m�Ȝh�"1[�P�G�Bo0�|��e����Ϳſ��Rr�֩/��@��삪���j��N&��+ �C�}O��   �   �@A�1�v�UE��x�����辒{��q��%��'.���0�n�-���$������徏���N����r��Q=�����D������R�=:����վz�o�P�97���Ҳ��sݿ���:��h�,�X`<�F���I���E��I;�R�+�������ܿ�v��.��X1Q����)׾�p��}VU��\ �����M�eP��   �   ����Yߩ�2 پ�U�"�G�=�,JU�Q�g�U�s��;w��r�Phf��sS���;�� ��S�l.־�s���Ā�7'G�i�!��X�)p��?�,���쵾���9Z/���i����2����߿:���O������%�(�r�$�^��j*�ؘ �zG޿i͹�h畿n2i��/�\,���Y��@^���UA�M����90$�JUJ��   �   �������F��/7��\��|��-f���Ĝ������������X̛��-���i~�jgZ�$5�zF�-⾨ͫ� ���b�G�#�%�!_�W�/�yU_��j��(�о����>�1u������3���UԿV��B� �*�		�:��� �����iҿ����1\��U}s��=���$Xоn;��Ѝ_���0�os��('��I��삾�   �   _�ᾁ����@���p�!Đ�('��k����x̿�aֿ{�ٿ%�տ�-˿:��5����T��=n�/?�e�S�߾������v�0w?��_$���$�.@��$x������ᾜ����@�"�p�����7$��6���[u̿�^ֿ�ٿڣտ�*˿t��ƈ���R���9n�n,?�c��߾�����v�Mv?�D`$�#�$��0@�<)x�'���   �   ��>�:5u�&����6��YԿ���� ���
	���� ����zlҿܕ��^��4�s��	=�@�6Zо�<����_���0�Tr�]&'�R�I�VꂾT���̈�,��L+7���\�hz��dc��������������
����ɛ�m+���e~��cZ�%!5�+D���<˫�������G���%��_�(�/��X_�hm����о�   �   �\/�|�i�6��������߿���Q������%�(�f�$�&���+�0� ��I޿>Ϲ��蕿�4i�Z/�y.���Z���^���UA�OL����J-$�QJ�����s۩�6پ���"��=��EU�j�g�I|s��6w�<�r��cf�|oS���;�� �8Q��*־ q�����$G��!��X�q�:�?� ��������   �   B�P�9���Բ�$vݿx�����^�,�~b<�L�F���I���E��K;��+�:��,����ܿ%x��/���2Q����\׾�q���VU�V\ �&��WK�M�*<A�"�v�{A������P��Vx�n�8�%��#.���0���-��$������2��ū��\���@r��N=�����C�3���p�R�4<����վ2|��   �    q� W���pͿ���/��81�ʥH�r7\��Bi���m��h��2[�ڜG�|p0�r������+�Ϳ�����r���/��A��`����j�N&�m* �d?�NJｴ/�
�/��:\�����Ģ������Ծ*�ө��_������l��tҾ����<��@��>�W��q+��I	�o���ݽ����j#��@g�^���XO��*�.��   �   �����ò�ۜ俘S���)�|�F��c��-{�y���C���$��ppz��wb���F���)���u忖���&�����D��
��ϼ���~��z-��D����ƽ켻�f�νy�����j<�1}a�҂�y㒾^~��o��v𩾉æ��<���/���Ԁ�9]�8�Ld�|Z�B�ƽ�K��В����𽑩)�I�z��q��6���-C��   �   ͥ�����P������\8�*�X�ăy��ފ�́��a����^�������oy�ZHY�ڠ8�._�JE���¿04vU�g����˾����)&4�����⳽�/��Kd��R����ٽX�l2�ݺ8��bO��a��7l�Ψo�(k��_�ɁL�L5�nm�D&�D�ѽ�7��4�������8�����;�/��U��H�Ⱦ����WS��   �   ����x-ʿR�v��dVA��	e�]W����,����I��Ɂ��������p�e��iB� !�F(��̿7���(`�����վp<��y�8����d��*m��y�{����������ʽx��5����YJ,��4��`7���3��i*����
�N콸�ý\���Af��1cl��X{�H{��h�o@4�I�����Ѿ���]��   �   ����JͿ��"Y"���D��Ii�J������������>��O8��X��Nj���E��#� <�VϿ�����c�[���hؾr&��x:���2���~���h�)|�򕽅j����ڽfG������F��"�,D%�!�!�Aw��p��/��
�ӽa��Zb����l�'Y��kn�����)�5��r��� վZ~�9a��   �   Y����,ʿ������UA��e��V��K��H����H��„����\���R�e��hB�r� ��'��̿�6���'`�����վ�;����8����nc���l����{����������ʽd��5����[J,��4��`7���3�j*����
�P콬�ýK���!f���bl��W{��z��*g뽱?4�������ѾC���]��   �   ������g���P���8�2�X�L�y�C݊�-����ޗ�I]��9���nmy�PFY�B�8��]�MC����¿�쒿ltU�'��߅˾�����$4������೽/���c�����Z�ٽE�`2�׺8��bO��a��7l�֨o�2k��_�ЁL�L5�mm�>&�"�ѽ�7��Ʃ��F����6�������/��T����Ⱦ����US��   �   񝆿����0���Q���)���F��c�$*{�e������}���lz��tb��F���)�R���|�h���y���!�D��
�`ͼ���~��x-�8B����ƽǻ����ν�x�����j<�}a�҂�x㒾_~���o��z𩾐æ��<���/���Ԁ�9]�
8�6d�#Z��ƽ�J��6���a�𽢧)�I�z�;o�����~+C��   �    q�rT���mͿ,���-��51�J�H�b3\�f>i�^�m�r�h��.[�R�G��m0���������Ϳ ����r���/��=������4�j��K&��( �T=��H�F/�µ/�j:\������â������Ծ.�ة��_������l��tҾ����<��	@��,�W��q+�8I	�B�
�ݽ����#� =g�����TK��J�.��   �   ��P�:6��CѲ��qݿ������,�|^<��|F���I�n�E��G;�^�+�*�����X�ܿ�t��<,��v.Q�����׾�n���RU��Y �l��5J�LL��;A�Ԛv�bA������D��Rx�n�9�%��#.��0���-���$������5��«��P���r�wN=�<���B��������R�D9��p�վy��   �   �X/���i�����`���߿��jN�2����%��(�`�$�^���(�&� �xD޿�ʹ�4啿�.i��/�((���V���[���QA��I���$,$�GPJ�����K۩�پ����"��=��EU�l�g�M|s��6w�B�r��cf��oS���;�� �7Q��*־�p����$G��!�W�}n�L�?�����굾T���   �   ����>�:.u�ؕ���1��8SԿR��� �Z�2	�V��' �U�뿭fҿː���Y��8ys�\=�$�ETо�8��B�_���0��o��$'�<�I��邾������!��B+7���\�fz��dc�����������������ɛ�p+���e~��cZ�&!5�)D���˫�>�����G���%�A]�h�/�S_�Ii����о�   �   �ᾕ��N�@���p�q����!��j���Hr̿6[ֿ�}ٿm�տD'˿K��߅��P��L5n��(?�#`���߾��E�v�	r?�~\$�^�$�},@��#x����͕ᾍ����@��p�����7$��5���]u̿�^ֿ�ٿ�տ�*˿w��Ɉ���R���9n�n,?�c�^�߾������v��t?�^$���$��+@��!x��	���   �   ����>�����L(7���\�>x���`��۾��~����������ƛ��(���`~�^_Z�b5�A����mǫ�������G���%�\�R�/�&T_�zj����оz���>�1u������3���UԿU��B� �,�		�<��  �����iҿ����4\��V}s��=����Wо;����_���0�op�2$'���I�r肾�   �   ����ة�Tپ�	���"��=�sAU���g�pws��1w�:�r��^f��jS�؈;�v� �,N��%־m��ֿ���G��!�9U��m�f�?������뵾]��(Z/���i�����/����߿:���O������%�(�t�$�`��l*�ژ �}G޿l͹�i畿m2i��/�4,��XY���]���SA��J�̅��*$��MJ��   �   �8A�{�v�o>��܏����辄u��j���%��.��0���-�(�$�U��������������r��I=����E@�������R��9����վz�d�P�67���Ҳ�sݿ���8��h�,�Z`<�F���I���E��I;�V�+�������ܿ�v��.��S1Q�����׾�p��5UU��Z ����aI�pJ��   �   -���/�6\�ε������_��ݐԾ���4��Z�����<g徶oҾR����8���<����W�Km+��E	��`~ݽ�����#�=g����4L���.�8q�@U���nͿ�	��t.��61�̣H�<5\��@i���m�ʜh�$1[�T�G�Do0�~��g���
�Ϳƿ��Rr�Щ/��@������ȝj�M&�C) �r<�dF��   �   ��ν7t�����f<�^xa�<ς�8����z���k��쩾����$9��M,��Iр�l3]�28�5`��S��ƽ�F��^���q���)�!�z�fo��ñ��+C�N���R²���vR�>�)���F��c��+{�_���.���)~���nz��vb���F�0�)�x���~���������D�9
�Qϼ��~�z-�qC����ƽ>����   �   ,b��k����ٽ��{/�c�8��^O�ea��2l��o�Gk�$�^�V}L�H5��i� #���ѽ13��J���~����4��?��&�/�BT��t�Ⱦ����US�����@���������>8���X�2�y��݊�途��ߗ�-^�����oy��GY�f�8��^��D��ݔ¿vU�b����˾����&4�3���᳽n.���   �   8�{����.�����ʽ��^4���SH,���4�D^7�T�3��g*����
���i�ýp����c���^l�/T{�y���e��>4�>���j�Ѿ����]�&���~,ʿ������UA�	e��V���������I��j���@��䍄�F�e��iB�  !�T(��̿�7���(`����վ�<����8���Cd���l���   �   ƷJ�Z\�ڡ������%��:��d��Dt	��$����?��z������
�׽ޭ��pM��Ko�TvC��1���D�P}��(�ʽ��_�w��M��NS���G�����⶿S�����-��HL�t�i��ȁ��������U���c���xj��2M��/�����,�A���񃋿xJ�b��A\����~���%�j�׽8����]��   �   l\�n�s�����9��?׽E8����v��/ ��-"�����h����� ̽����R���S�Z��C��P������?˽۽��Dt�m{��q$	�
kD������JK�ta�z/+���H�T�e��x~�뼇�P���*�����~�� f�n�I��.,�L}�yu�]	��C���,G�!p�tf��;{��6$�Y�׽.��r~i��   �   =���d֝��������M��$��,8���G���Q��`T�hP� �D�]24�<1�*��x)�P���y���gx��t�Nu����̽A����j��W��|���A;�RX���򫿥ܿ�
��L#�f�>��zY��p��w��j���:���o�LhY��;?���#����v�ݿ�|������M�=�q���ߴ��bq������ؽRl��Ty���   �   <s��eܽ6f�9'�.�H�
�h�-�������ꢔ�ּ��ɓ�I���V���Qc�ڢB�KT!�x*�x�ϽSw���ۙ��!����н2����\�Fˤ����
�,��o�F���˿O9��b�� 0�ZSG�\�Z���g��el�~g�T2Z���F��/�<(�e�����̿Z���p�0�.�`0��%���,rb����ߚ۽jT���q���   �   �T��5��C��q��Ɛ��#��j伾)(;n_׾шھ�X־�;˾aH����h����j��l=�9�����,�Ƚtc��VٽP����K�4)��G&پɹ���U�Z����&��D�����z��0r1�L�A��\L���O��K�t�@��}0�6���T�����V���	����V�����x۾Yp���UP��l�T��ȑɽ��ӽ�   �   ң+�N[�����n&���ξ��`a��&�������i�����a��N�"˾z��F���U�p&�L��k�%+轆O
�'�9�*����z���;� L9��mw��D��ќſ���.	����b'���/��c2��/�|&���D�5=���Ŀ枿�Zw���9����t߾������9=�>���?� [��	��   �   %Xh��������k ���>c(��|=���M�8SX��[��yW��iL�Ys;�R#&��T�p�뾜X��{瓾�c�"(/���\2 �mx��)�g�e��/���"�����O�w���b�����ǿ+��r����w�&��,��Ҧ�Ŝ ����_9ƿgr���;��\�N�;@��9�۵��.g�8+�n��W��l�<�3��   �   �K���˾�|���"�p5D�րd��y��9����u��H����呿܄��Y~��a��A��d ��� ���Ǿ6旾f�d���/�5���r
��#���E�c8��X��5����(�V�Y��͇�gM��T����fԿ�$濥8񿒯���I�3��lҿ1���S������X�$�'�#�������#�����E���������
�2�Xzh��   �   fEȾ���TW+�t�U��Ѐ�;˕��+��Vh���H��L¿b������L������W�~��ES�T`)��e�?<ƾ�Ⓘ�;Z�)����E�Q*��\��B���AȾB��T+�x�U�F΀��ȕ�)��Ke���E��8¿l���#��΅��_����~��BS��])�4d��9ƾ����:Z�H)����_F��*��\��E���   �   �9����(��Y��χ��O��:����iԿ&(�<����M�1�俿nҿ����Q�������W
X��'���������<�����E�����������2��uh�qH��y˾�y�[�"�q1D�I|d�pw������s������㑿o����T~�>�a���A�b ��� ���Ǿ䗾��d�c�/����Rs
�j%�ٙE��:��<[���   �   w��ԷO�o���������ǿ8��������x������`��(� �E��d;ƿt��=��T�N��A��;�����$/g�58+���TV��i�j�3��Rh�����������ߍ��_(��x=�B�M��NX���[�=uW��eL��o;�& &�R�!��DU���䓾hc��%/�۰�*2 �:y��)���e�I2���&��   �   �N9�qw��F��0�ſ��쿶	�n��6'���/�fe2��
/�&�J��l� ?뿁�Ŀ@瞿v\w��9�����྾����9=����=��V�
�	���+��H[����;"���ξ³�1^�B#�3��D����������\��˾$w������$U��&����~i�T+轎P
�E�9�����D}��n=��   �   N�U�ꛎ��(�����D������s1��A��^L�l�O���K���@��~0�D���U�
���W���
����V�����y۾�p���UP� l�N�⽆�ɽJ�ӽqN��$���C��|q�PÐ�����߼�)#;DZ׾��ھ�S־67˾0D��\��W|����j��h=�R�����ɼȽ�b��ٽ���K��*���(پ����   �   �o������˿N;����>0��TG��Z�d�g�~gl��g��3Z���F��/��(�c�����̿�����p���.��0��Q���rb���)�۽�Q��En���n���ܽ�b��z'��H�6�h�����P���^���J����œ���T���Lc���B��P!��'���Ͻ�t��:ڙ�r!����нp���\��̤�0���,��   �   FY�����	ܿ~��M#���>��{Y��p�y��k��<���o�iY�(<?�4�#�8��Ьݿ�|�����b�=�o���ߴ�-bq���1�ؽTj���v����rҝ�D����뽕J�;
$��(8�\�G�D�Q�R\T�.	P��D��.4�(.����L%�|��dw���dx���t��u����̽~����j�5Y�����3C;��   �   �������LL�b�"0+�v�H�*�e��y~�W�������w���&�~�Bf���I��.,�H}�_u�8	���B��R,G��o��e��0:{�$6$���׽���{i��\���s����6���׽�4��ڡ�W�� �m+"����D��������|̽毧������Z�� C�7�P�H���A˽����Ft��|��K%	�+lD��   �   ����@㶿���R��Z�-�TIL���i��ȁ�������E���E��hxj�v2M�z/����,쿺���{���VwJ�˷�_[��9�~���%��׽���]�.�J��X\�0�������t$����� ��!t	��$����O��������}�׽d����M���o��wC�w�1���D�l~����ʽ����w��N���S�^�G��   �   3���C��iK�za�r/+���H��e�nx~�����������؊~�" f���I��-,��|�pt�{��DB��{+G�?o�%e�� 9{�p5$���׽��Czi�\���s�褒��5���׽u4��ա�X�� �m+"����G��������|̽௧�������Z�k C���P�����<@˽O���Et��{���$	�^kD��   �   :X����Uܿp
�8L#���>��yY��p�zv�6j��n9�~�o�gY�x:?���#����ݿ�{�����ʛ=�P��޴�%`q����l�ؽ$i��
v���~��ҝ������뽂J�2
$��(8�Z�G�E�Q�V\T�4	P��D��.4�-.����:%��{��&w��dx�T�t��t��L�̽;����j��W��z���A;��   �   �o����p�˿_8���� 0�JRG��Z��g�
dl�@|g��0Z�.�F���/�'�\���!�̿�����p�l�.��-��9���Gob�D����۽8P��/m���m��ܽhb��z'���H�'�h�����N���`���M����œ���"T���Lc���B��P!��'�5�Ͻt��Rٙ����l�н���`�\��ʤ�0���,��   �   ��U������%�����&��t���p1�ȱA�[L���O�4�K���@�|0�����S�o���T��D���V����"v۾Dn���RP��i�Z�⽏�ɽ��ӽ�M������C��|q�BÐ�����߼�)#;GZ׾��ھ�S־>7˾6D��`��Y|����j��h=�$����Ƚ�`��Rٽg����K��(��R%پ���   �   �J9� lw�oC��L�ſ��	�^���'��/��a2�/��&�8����y:뿑�Ŀ䞿YWw�/�9�����ܾ�i���46=�H���9��T�V�	�:�+�TH[�����%"����ξ���.^�B#�4��G��
��������b��˾!w�������U�^&����g�Z(�BN
���9�J���gy���:��   �   �����O�-���������ǿǙ������Nu�\��`����� ��快6ƿp���9��-�N��=�+6�����)g��4+�@��T��h���3�jRh�����s������֍��_(��x=�A�M��NX���[�AuW��eL��o;�* &�R� ��:U���䓾c�G%/����0 ��v�&)�^�e�h.��� ��   �   92����(���Y��ˇ�gK���}���cԿ�!�l5�6����F��}��hҿS���Ě���|��X�0�'�����H���������E�A����X����2��th�7H��R˾�y�O�"�h1D�D|d�nw������s������㑿r����T~�C�a���A�b ��� ���Ǿ�㗾�d�{�/�C��q
�"�ДE��6���U���   �   �>Ⱦt���Q+�l�U�h̀�cƕ��&���b���B��%
¿X���$����������~��>S��Z)��a��5ƾ�ݒ�F5Z�j)�x���B��*��\��B��QAȾ2��T+�m�U�B΀��ȕ�)��Me���E��;¿q���(��҅��b����~��BS��])�-d��9ƾ����<9Z��)����DC�2*� \�A���   �   F��N�ʾ�w���"�*.D�hxd�8u��"���ip��㜔�]�������O~���a���A��^ �Ƌ ���Ǿ����G�d�+�/�$��p
��!���E��7���W���4����(�K�Y��͇�cM��Q����fԿ�$濩8񿓯���I�9��lҿ5���V������X� �'�	�������������E���5�����E�2�6rh��   �   �Nh�l���������)��P\(��t=�2�M�^JX��[��pW��aL��k;�|&��N�����P��pᓾ�c�l!/�8���. �v�4)�`�e�y/���"������O�s���]�����ǿ)��r����w�(��0��Ԧ�Ȝ ���c9ƿjr���;��\�N�2@��9⾔���-g��6+�&��T��g���3��   �   ��+�zD[�]��������ξ���R[� �φ�������f��d����˾�r��:����U�A&����Xc潭%车M
���9�����gz��;�L9��mw��D��Ϝſ���,	����d'���/��c2��/�~&���F�8=���Ŀ	枿�Zw���9����?߾�6���n8=�f��@:�ZSｰ�	��   �   �I������C��wq�.�������ۼ�~;FU׾�~ھ}N־F2˾�?��2���x��Z�j��c=���Ķ��Ƚ�]��'ٽ�����K��(��&پ�����U�X����&��A�����|��0r1�L�A��\L���O��K�x�@��}0�8���T�����V���	����V�����x۾p���TP�.k�*��͋ɽ��ӽ�   �   Ik��#ܽ�_�Gw'��|H��h�����������ĵ��*�����P��Gc���B�L!�$�`�Ͻ�o���ՙ�b����н*��6�\�ˤ���� �,��o�D���˿M9��b�� 0�XSG�Z�Z���g��el�~g�V2Z���F��/�>(�i�����̿Z����p�,�.�I0�������qb����ڗ۽P���k���   �   '}���ϝ�ȯ������G�$�2%8�n�G��Q��WT��P���D��*4��*�T����<w��8s���]x�J�t��r����̽�����j��W��r���A;�PX���򫿣ܿ�
��L#�f�>��zY��p��w��j���:���o�NhY��;?���#����y�ݿ�|������L�=�i���ߴ�7bq����Ħؽ�i��~u���   �   t\��s�����84���׽�1��:����� �X)"���.����*��~y̽鬧�h����Z���B�)�P�6����>˽����Dt�_{��m$	�kD������IK�ta�x/+���H�T�e��x~�뼇�P���+�����~�� f�n�I��.,�L}�{u�_	��C���,G�p�ef���:{��6$�d�׽����zi��   �   ��-��!=�-b���bҥ�J�����ؽ�����Í���?��㽶	ν�8��������o���:�g��&���,�R��X���z��R�����b���*��l�����o�ɿ^�����(w.���E�xNY�>�f�HFk�ڗf��vY�`!F�<-/�­������̿#v��_�o�t�-�?l󾀁���[�����W{�8z>��   �   ��<��Q�QH|�U*��฽��ֽ�@��������Q
����`��Zk�uɽ������5U��(��������X����dV��QO��2��)e��"(���h�Z����ƿ#��@w���+��eB��qU��Kb�~�f�&Bb��~U���B��E,�JE�����`�ȿ�圿=�k�&�*�r���*�X��������.���bH��   �   1�j�C燽��Re˽o�,�O��+�۟3���5���1���'�!��8�X2�fc��U쒽F+h�V�B�5�?�HAj�ML���%�PmG��G����߾�J ���]�������{9�����#���8�8zJ�h4V�\EZ��V��BJ�<�8�l�#�S��~쿵r��Wr��֢`���"�6#�G�����O���	��v��t����f��   �   ���ҽ�mu�]����,�"^H�n�`�vs��'��8���}�0ko�f�Z��3A��$�����ؽ̪��,��%�w������F���u;������ξ�� M�Q݈����
ڿ&���w��~*�t :�*1D�$�G�d�C��|9��	*�,;�����ڿ���gʉ���N����v�Ҿ6?����B��n�3���ti��~���   �   X�׽���g)�NP��wy�!���b���2���ϸ�N_������񭾱=��C㌾��p�AQG�����K��h"ƽ�"���3���ܳ�����,�w�~�|����v��X7��u��ם���ÿu��f �~���%��.�:[1��.��9%�����d���W�ÿR��"�u�r8�����d��#���3�����@½��������   �   ���|=��o��<������0�ξ-�c���_���|����c�����侉�ʾvs��������f���4������ݽ˿�����������Sa�$����御��iT����z��s�̿��N�����-�<u�į�v:�0���U�<H˿��������UT�w'�%�+ţ��>e�bO"�!+�$�ͽͽ����   �   ��G��������HξV��ϑ�3�"� �0�6�9��i<�q�8�6/�Њ �*��`��ɾ☡�(|�=�@�* �h�c׽�%���!�C�h��\����P�x/2�"<f��~��뀬��"ȿ,R࿌�s����J������|��f޿Jƿ����Yc��#�d��g1�W����������F��w�����vར4��O��   �   o���|��0(�h���v(�6DD���\���o���{�����z�.�m��DZ�LxA���%�-2	���۾�Ԫ�۟����B�<I����@�{��?�(�+�e���0,پ!���;��xi�E���yo���g��j�ƿ'�пb�ӿ�Ͽ$nſd������)����f�c*9�|x�P�׾q��xJe�b)�&������89���G��   �   �󫾆
侬�˖7��i]��‿9ې��?��N����e��Q����ST��t�~��eZ���4�v����ྯ���{�R':�X���0�����,��<�t�~�x���
�]�7��e]�t����ؐ�=������c��N�����'R����~�MbZ�A�4�n����ྈ���$
{��%:����d1��T��/�p�<�I�~��   �   �/پ����
;�h|i����� r��wj��P�ƿ�пO�ӿ�Ͽ�pſ����!����	��o�f��,9�#z���׾��\Le�F)�&�Q����k6���G������x��z#ྂ��Cs(�K@D�8�\��o���{�R��v�z���m�AZ��tA��%��/	�h�۾Ҫ� ���U�B��G� ~���A������(��e������   �   S�022��?f�����K���d%ȿU࿕����L�o�����>i޿�Lƿ�����d��d�d��i1���=��������F��w�`��#t�0���K�L�G�����@ ���CξyP�������"�=�0�R�9��e<���8��2/��� �d'�@\�|ɾ����|�4�@�.�Y~�6c׽2'潙����C����f����   �   ����kT�����|��Ӊ̿X����^�H/��v�:���;�\���W��I˿�������WT��(��&�ƣ��?e��O"�/*��ͽpͽF������=�*�o��8��x���D�ξ�y辌���Z���y�����������L�ʾ�o�����@�f�E�4�\����ݽ�ɿ����w�����|Va�\&�����   �   �Z7�ku�wٝ���ÿ��꿨�ީ���%�x�.��\1�&.�;%����fe�=꿀�ÿ7��u�u�
s8�#���e��b#��3�$���>½��������׽���	)��HP�xqy�����^��{.���˸��Z�������:��#�����p��LG�<���F���ƽ� ���2��Iݳ�����,���~������x��   �   M��ވ������ڿ$���x�*�*��:��2D�x�G���C��}9��
*��;�8���ڿ�����ʉ�8�N����݅Ҿ^?����B�Xn�����8g��t
������̽�"o뽒����,�YH��`��ys��!��5���}��eo�q�Z��/A�m�$���شؽ�Ȫ��*����w��d�� I���w;�������ξk��   �   ��]�������:뿰����#���8�F{J�|5V�bFZ��V��CJ���8���#�fS�'�s���r���`���"�2#�*�����O��	��u�����
�f���j��ㇽ���_`˽Vi�w)��K�f�+�	�3�ض5��1���'���u5��-��_���钽@'h���B��?��Aj�oM���&�oG�I��֠߾�K ��   �   ��h�����ƿ$���w���+�(fB�lrU�JLb��f��Bb��~U���B��E,�VE�����I�ȿ�圿��k���*��~�a�h�X�������G-��|_H�P�<��{Q��C|��'��#ݸ�`�ֽ_=��������O
�B��8���h�ɽ����� ���2U���(���-���X�D���`W� SO��3���f��#(��   �   d�l������ɿ����&��nw.��E��NY�Z�f�JFk���f��vY�$!F��,/�~��,���	̿�u����o���-�;k󾼀��ɏ[�����~U{��x>�H�-�� =��+b�����ѥ�������ؽ�뽝������ @�8��
νD9��<����o��:���X(���-�R��Y���{��R�W���d�*��   �   ��h�����ƿ#��<w��+�ReB�tqU�8Kb���f��Ab��}U��B�E,��D�����y�ȿ圿��k�$�*��}ﾯ�z�X�L�������,���^H���<�t{Q�`C|��'��ݸ�P�ֽN=��������O
�@��;���h�ɽ����� ���2U�o�(���������X������V�RO�&3���e�2#(��   �   ��]�w�����9뿘����#��8�~yJ��3V�XDZ��V��AJ�<�8���#�BR�B}�uq��Kq��%�`�V�"�C!�ד����O���	��s�������f���j�oㇽ���!`˽$i�h)��K�^�+��3�ض5��1���'���u5��-㽲_��e钽�&h��B���?��?j��K���%�WmG��G����߾�J ��   �   ��L��܈�y���N	ڿ����v�~*�j�9��/D�СG��C�,{9�n*�
:����B�ڿ����&ɉ���N���2�Ҿ�=��/�B��l�p����e��Z	��� ��q̽��n�i��k�,�YH�Ӝ`��ys��!��5���}��eo�t�Z��/A�k�$�����ؽTȪ�*���w�:d��F��zu;�ʛ��Z�ξ���   �   �W7�pu��֝�}�ÿ�꿈��r����%���.��Y1�@.�L8%�f��>c�� �[�ÿ���_�u��o8����b��6!��3�,��<½׻��������׽����	)��HP�Qqy�v���^��w.���˸��Z�������:��'�����p��LG�)��:F��Sƽ���,1���ڳ�j�� �,�P�~�����Uv��   �   ����gT���Xy��υ̿��&����D,��s�4���8�����R��E˿����G���"ST�?%��!羫£��:e�_L"��%���ͽeͽ��t��{=��o��8��c���6�ξ�y辉���Y���y�����������N�ʾ�o�����+�f��4�����ݽ�ǿ�p���j�轿���Qa�#��M���   �   �O��-2��9f�|}��*��� ȿ�O������I�q����y��c޿�Gƿp���La����d�"e1�3�d���7���#F��t���q� .��K���G����� ���CξbP�������"�<�0�S�9� f<���8��2/��� �g'�C\�|ɾ�����|���@����|`׽#���V�C�. �������   �   �)پt��u;��ui�����gm��Ze����ƿX�пw�ӿ)�ϿEkſ�������������f�4'9��u�_�׾q���Ee��)�	�����n5���G�j����x��Y#�u��8s(�B@D�2�\��o���{�X��|�z���m�"AZ� uA��%��/	�a�۾�Ѫ�ڝ����B�
G��{���=����X�(���e���   �   -�����7��b]��ހ��֐��:�����m`���K�����O��"�~�N^Z���4����,������{�o!:�6��A+��+���+�1�<�ۇ~�D����
�P�7��e]�p����ؐ�=������c���N�����+R����~�RbZ�C�4�m�����h����	{��$:�x���-�����+���<� �~��   �   ����v����6��np(��<D�_�\���o�h�{������z�m�m��<Z�qA���%�
-	���۾KΪ�
�����B�"D��w���;�����(�b�e���,پ���;��xi�@���vo���g��j�ƿ)�пd�ӿ�Ͽ)nſh������+����f�c*9�wx�8�׾C���Ie�^
)��
�4�����,4���G��   �   ��G�����D���+@ξ�K��܋���"���0���9�b<���8��./�2� �=$��V�vwɾ/�����{�S�@�H��w�]׽�!潃��'�C���'����P�j/2�<f��~��瀬��"ȿ*R࿍�u����J������|��f޿�Jƿ����[c��$�d��g1�N����h���F�iv�����p�*,��9I��   �   *��0=�p�o��5������ξ�t����p���v����/������m�ʾ�k������J�f�n�4�p��C�ݽ8Ŀ����C��ӽ��Ra��#����従��iT����z��q�̿��N�����-�>u�Ư�x:�2���U�?H˿·��	����UT�r'��$��ģ�
>e�RN"��'�R�ͽ;
ͽ���   �   ��׽>��n)�@DP�ly�S���zZ��x*��FǸ�wV��Q����譾$6���܌�n�p��GG����%?���ƽ���4.���س�q���,��~�L����v��X7��u��ם���ÿs��f �~��
�%���.�:[1��.��9%�����d���Y�ÿT��$�u�r8�����d���"��3�p���<½?���Ե���   �   ����ɽ�j�t����,��TH���`�ts����2����|��_o���Z��*A��$�=��b�ؽ4ê�&���yw��넽���E��Pu;�䛌���ξ�� M�O݈����
ڿ&���w��~*�t :�,1D�&�G�d�C��|9��	*�.;����
�ڿ	���hʉ���N����^�Ҿ?��,�B��m������e��C���   �   :�j��ᇽ����\˽�d��&�zH���+�h�3��5��1��'����D2�)(��Z��@咽�h�x�B�j�?�C<j��J��%��lG��G���߾�J ���]�������{9�����#���8�8zJ�j4V�\EZ��V��BJ�>�8�l�#�S��~쿷r��Xr��բ`���"�*#�.�����O��	�'u�������f��   �   J�<�"zQ�GA|�&��#۸���ֽ�:�Z�����N
�k��� ��e��ɽ��������%.U�r�(�%�����2�X�+���V�^QO��2��e��"(���h�Y����ƿ#��@w���+��eB��qU��Kb���f�(Bb��~U���B��E,�LE�����`�ȿ�圿>�k�$�*�l�����X�O��&���f-��6_H��   �   ����h&�-�D�i4m��Ќ�a��H���!ýU ˽��˽�LŽ�շ��n��t����Ge��`1�!7�V�¼b"��8Sļ�Y����Rսf8+��
��Zsľj:��D����A���Cѿ9���6{��#���2���<���?���<�@�2�
$�������N�ҿmf��ѹ��F3G�J�1�ʾ�Q��C�8��C����Y�i~'��   �   �&��R7��vZ����ʜ�QŴ���ɽ�Qٽ�B⽝r�P�ܽν���z<��Fق���L����������T�ּ�b�z:��6|ӽ��(���g����
�B�@�]�� ��οc����B�T.!�&�/�|[9���<�4T9���/�Z_!���k"��_�Ͽ����6�����C�����CǾE+��f6����@䞽A�]��~/��   �   	�K��k���� 2����ͽUJ�Db��������&��*�HI	��t��
0ؽ~���J}���^�Ͽ)�ʾ	�XE�C,��؁��fν�"���x�������T�7�v�D���B�Ŀ��������f'�nQ0��`3�x00�?'�����]��e�ſ������x�np:�i�}̽������.�B��
����j�\+H��   �   +���D���OȽR���6��(�w�;��J���S��1V�0Q��UE��3�ֺ��c�$@ٽ	۪�^���l�O�e�7���G�␅��Qǽ[��4Tg�z̪�z����)��Zc������M��ܣڿ�|���?�r����"�:%��O"��9�����!��¯ڿk���\R��� e�ץ+�[�����8�p��V#���޽x���V8���os��   �   *�.�:���J/�0Q���q��b��:����{�� a�����m̏�^��8�g��iE�oU"����JȽg]���,�|ar�^֌�7��x���Q��p���+۾Z���^K��[������=cĿK���g����
������D,�
�mC������ÿ�`��􀃿L�����ݾ�����X�{��&Խ�`����������   �   ���!��#I�4x������R���T��ԹѾ��۾��޾kھ��ξ~0���=���ݎ�d�k���<�/������i���J���V���ܺ��� �=u9�����U�� ��1 0���c����
Ԫ��Lƿ&e޿�+�����vf �7E���￧�ܿ*�Ŀ�Щ�mb���#c�0�|��谿� ����>����ʽ)��������
ǽ�   �   ��'���Y�Ⰺ�y�#�ξ�:���W��l���0���H�B��1�꾗�Ⱦ"�������N�h����/���Ơ��D���'�/U!�6^d�ɔ����ܾ����?���n�ٽ��$�������s˿�eտ�ؿ{�Կ�0ʿ�
������s����l�Ⱥ=����`OܾҦ��'�e��/$����^�Ľ�n��^�ϽV'��   �   O_]�&u������A6辦����"�$N7��:G�^4Q��LT��;P�:iE���4��" �E	���vl���Ԍ�L;U�r��/��ǽ����[׽�
�Or>�H냾(@��4+�#'���A���i��������Q���9���̰�M���"ޤ��z��8�����f�r?��H��g�^W��������=��c�R�ڽ�eĽ�н����%�&��   �   {
��񇽾�3���_�v�7��*V�k�p�4タ�g��r���ֈ��ׁ��9n�6S��4�ѿ�Y��Aƹ����Y�N�����d�'"ɽ҂ʽ�|��]�ӭS����O���/���\��7��&V�4�p������e���o���Ԉ��Ձ�Q6n��2S�e�4������ﾺù�� ����N�I���c�v"ɽ��ʽ����`�ԱS��   �   LC��X/��)�&�A���i�	��������<��ϰ�����Wि�|��������f�vt?��J�yj�TY��
Â�P�=�Xd�[�ڽTdĽ#�нV���Ǆ&��Z]�r��ٌ��w1������"��J7�7G�l0Q��HT�+8P��eE�_�4�*  �� 	�U�⾍i���Ҍ�-8U�b���,���ǽ��� ^׽-�
�u>��탾�   �   $ݾ���?���n�ۿ��b��𓻿Kv˿uhտ|�ؿ�Կ�2ʿ��������t����l���=����bQܾ)�����e�{0$���[�Ľ�l����Ͻ�$�Ǆ'���Y������﫾��ξ>5���7��2��]-���d���������Ⱦ���L���z�N�we����j���r���f����)꽄W!��ad�M����   �   Ɍ��"0���c�a	��֪��Nƿ�g޿�.����g ��G��N�￞�ܿ��Ŀҩ��c���%c�p0�k��&��������>�.�šʽT��������ǽ����F�I�".x�����N��P����Ѿ��۾��޾Nfھ0�ξt,��P:���ڎ���k�5�<�\�����Mg���I��W��޺�F� ��w9����$X���   �   ��?aK�b]������"eĿe��.j��
������`-�
�0E��?�⿻�ÿ�a������2 L������ݾE�����X�����Խl_��l���@���-(佋��SF/��*Q���q�X_�������w��T]��,��ɏ�[���g��eE��Q"���VFȽrZ��)�1`r��֌������p�Q�]r��x.۾�   �   ��)��\c�𩒿O����ڿ�~���@�|��Ȏ"�;%��P"�p:�����"����ڿ%����R��Oe�Y�+�����r��{�p��V#�J�޽@����6��|js�Ѡ���?��~JȽ��������(�خ;��J���S��,V�!+Q�QE�ܦ3�:���`�;ٽת�l���k�O�1�7�>�G������Sǽ����Vg�8Ϊ������   �   ��7��v�M���u�Ŀ]��������hg'�<R0��a3�&10��?'�b��d������ſ�G�x��p:�y�z̽�~�����.�e��轞�� j��'H�Z�K��k������-����ͽ�D�V_��������#��'�nF	��o���+ؽ����8z��\�^�b�)���	�kD��,��ف�Xhν��"���x�8������   �   N�@���� ���οN���0C��.!���/��[9� �<��T9��/��_!� ��~"��]�Ͽ���������C�p��(CǾ�*��� 6����'㞽��]�E|/��&�#O7��rZ�����ǜ��´�ȝɽ�Nٽ�?⽎o�h�ܽ\ν<��x:���ׂ�>�L������������ּ�c��;���}ӽ��(����Nh��w ��   �   \D�D�������Cѿ����l{�D�#��2���<���?��<��2��	$����6����ҿf��n����2G��I�X�ʾIQ��J�8�bB���T�Y��|'�c��^g&��D�k3m�9Ќ��`������!ý/ ˽��˽�LŽ�շ��n��ή��XHe��a1�%8���¼�$��Vļ�[����}SսY9+�)��0tľ�:��   �   ��@�{��. �� οY����B�..!��/�*[9�N�<��S9�P�/��^!�j��}!����Ͽꪧ�������C����OBǾR*����5����_➽��]�r{/�_&��N7�OrZ�t��lǜ�n´���ɽ�Nٽ�?⽉o�c�ܽXν7��t:���ׂ�$�L����"��P�����ּ�b��:���|ӽ�(�g��g����
��   �   0�7��v�
�����Ŀ��뿲��~��f'��P0�(`3��/0�L>'���J�� ��,�ſ����2�x�o:�S��ʽ�`����.�E��o�����i�&H�0�K��k�;����-��z�ͽ�D�B_��������#��'�lF	��o���+ؽ����"z���^���)���	�fC�
,�v؁�xfν�"���x�����ԅ��   �   ��)��Yc�,����L����ڿ�{��J?����̌"�9%��N"��8��������ڿ볶�Q��n�d�,�+�����7��e�p��T#�U�޽(���5��Jhs�����?���IȽ����T���(���;��J���S��,V�+Q�QE�ۦ3�6���`�;ٽ�֪�*�����O�Ƶ7���G�菅��Pǽ����Sg�̪������   �   ����]K�A[�����
bĿ׽�/f����
��~����+��	
�&A����⿔�ÿ2_������L�N��6�ݾ�����X�
���Խ�\���������h'�=��F/��*Q���q�H_�������w��R]��,�� ɏ�[���g��eE��Q"���FȽ�Y��N'�u]r��Ԍ��������~Q��o���*۾�   �   ���0���c�����Ҫ�Kƿ5c޿�)����2e ��B�����=�ܿ��Ŀ�Ω��`��� c��	0���������}�>�b���ʽ�������� ǽ�������I��-x�ꖔ��N��P����Ѿ��۾��޾Ofھ4�ξw,��P:���ڎ���k��<�0�����[f��/H���T���ں��� ��s9��
��2T���   �   ��ܾ<���?�%�n�^���_��x���xq˿gcտ[�ؿ�Կ.ʿy������q���l��=�3���Kܾ����e�k,$�@��`�Ľ�i����Ͻ�#�:�'�,�Y�����y﫾o�ξ(5���3��0��^-���g���������Ⱦ���A���N�N�,e����᣿����ڟ���$꽡S!�\d�U����   �   >��f(�F%���A��i�*����	��:7��ʰ�я���ۤ��x�������f��n?�>F�yc�T��2����|=�p`���ڽ}`Ľt�нj����&�/Z]��q������T1������"��J7�7G�j0Q��HT�-8P��eE�d�4�,  �� 	�Q�⾃i���Ҍ��7U���6+��ǽ���X׽o�
�"p>��郾�   �   ��������+���Z�b�7��#V���p��ނ�lc���m��U҈��Ӂ�%2n�/S��4�ͺ�K����������h�N�����]�ɽIʽ�z�]�6�S����$����.���\��7��&V�0�p������e���o���Ԉ��Ձ�V6n��2S�h�4������ﾭù�� ����N����}a�Qɽ�ʽ�y��[���S��   �   >W]��o��։���-�s����"�VG7��3G��,Q��DT�<4P��aE���4�� � ����⾙e���ό�03U�m��=&�H�ǽ\���X׽�
��q>�냾�?��+�'���A���i��������P���9���̰�Q���%ޤ��z��;�����f�r?��H��g�GW������(�=��b���ڽ�aĽ�нn���6�&��   �   ց'���Y�>���r쫾��ξ�0�=��L����%*�c�I����p��:�Ⱦ�����K�N�Pa����̟��n���{���u$�ET!��]d�������ܾ����?���n�ս��������s˿�eտ�ؿ�Կ�0ʿ�
������s����l�Ⱥ=�~��QOܾ������e��.$�X����Ľ�i��#�Ͻ\"��   �   ����(
�I�)x�����AK���K��w�Ѿ�۾��޾Qaھc�ξ�'��D6��׎���k�.�<�>������a���D���R��~ٺ��� ��t9����VU�����# 0���c����Ԫ��Lƿ&e޿�+�����xf �<E���￫�ܿ-�Ŀ�Щ�ob���#c�0�v��а�����%�>����ʽ��������ǽ�   �   �궽c#佁���B/�7&Q�|�q�N\��U���Ut���Y������ŏ��W���g�=`E�OM"����?Ƚ-U��# �;Xr�ӌ�������[Q�Rp���+۾O���^K��[��󌣿;cĿL���g����
������F,�
�qC����⿁�ÿ�`������L�����ݾ������X�Ȧ��Խ�]��B�r���   �   :���b<��3FȽ����R��0�'���;�v�J���S��'V�&Q�'LE�A�3����\��4ٽ�Ѫ�������O�T�7���G�t����Oǽ����Sg�X̪�b����)��Zc������M��ۣڿ�|���?�r����"�:%��O"��9�����!��¯ڿl���]R��� e�֥+�R�������p�eV#�i�޽$���
5���fs��   �   T�K��k������*����ͽX@�\�������^ ��$�TC	��i��'&ؽ�{���u���^���)��	�r?��,�.ׁ�qeν��"�Q�x�����څ�N�7�v�C���B�Ŀ��������f'�nQ0��`3�z00�?'�����^��f�ſ������x�np:�f�p̽�������.�@�轌���e�i��%H��   �   &��M7��pZ�@���Ŝ�|���`�ɽ4Lٽ�<⽃l�P�ܽKνG	���7��Ղ���L����L��N���f�ּm`��9���{ӽg�(���g����
�@�@�[�� ��οc����B�T.!�&�/�~[9���<�6T9���/�\_!���l"��c�Ͽ����7�����C�����CǾ:+��B6�Z�ｃ㞽 �]��{/��   �   9��/"�p�8�3oV�14v��&��w������X��R����5�� L���dw��UM�9��v������:���
� �;����~�2��w���K���P�_���v�o���hR�����uT���b˿�������r3�n��B-������X̿����OQ���LU�����J�_���ib�
x��Kν�z���?J��#��   �   ��!��`/�PJ��k���������`^�������H����|C������������k���:���	�ȗ��4v� 8�4O[��i����3�a��Ї���M����e�ݾnY��O�ۅ�U����HȿUu�ڄ�\��z6����D1�`��B������ɿ�ɧ������Q��N��z� f���^�F:�f�˽*���2�L���(��   �   ��>�L�W��~�Ζ��N����ƽlڽ:��Ȁ�<��罙�׽{���,ߤ�Vl��2�O������ּ�$��Ό��x�ۼTf7�NQ��=���g�D�q���N�Ӿ�!�LjE�BT�����<����ݿ;��Na��L����6��F��(��'1޿����ڟ�-�����G����mپ�����T����x^ŽҊ��T��:��   �   �q�0:#����Ͻ��'�
�	��q�$�(+���+��'���Y���0��0eͽD��Q�z���9����3�V>�h�>�$9�����7������þ1��C6�s�k����������Ϳ���E���v�����"i�1���F�+LͿ0��lo��f�l���7�K�	�9Ⱦ������D����һ�R���G~c���Z��   �   㝽ܯ½h����,��F�~H\��Hm��jw�*�y�'�s���e���P�S7�
�CH��ǜŽ��b��4��%+���L��H��l�۽'�%���t��B���
��"���R�/��������m���Ͽ����!����k࿍Dοw����>��љ��L:S���#�QV���{��aM}�|�0��J�� ��p ��FS|��х��   �   �Xѽ8����&��K���r�-싾Q�����̰�~۲��OW������V��(�b��!:�^����������)�^�y�c�
-��ȎȽ����#V�m����Ҿ"�8�6�_d�ɰ��67������lÿE"Ϳ�Gп]�̿k�¿����t7��^∿oEc�Z#6����{Ӿ��W�[�_��Q�ܽhO��l������!���   �   rb
��2���b�ً��K������BTپ��v
��dZ���6���辵:Ծ�����������R���"������Ҹ�=瑽���؋��#*��_ �V�6�r怾ie��!�쾌A���?��.g�b����f��t��禬��F��f��i���V9��m���d��=���,6�t���p퀾��8��S�NFĽX��>��`�����ս�   �   �4�u�l��6������6Qᾐ��q0�/����'��;*��&���~��������ھ�����u��+�_�y�(������v���њ�o��� n��zݽK����T��0���)���9��3����;�T�Z�.1v��ǅ�Y|������a����Մ�J�s��X�� 9��5�q"��mѽ�����*Q��t� �޽����ԝ��:���Ͻ?��   �   ��g��"��G�ľ2�����+�nA��QR���\��)`���[��|P��?��!)�����E�/[���:��%$_��$��"򽵁�������Ơ����ɨ����+�I�g������ľ���9����+�|A��MR���\�B&`��[��yP��?�>)����5B�zX���8��;!_��}$�6 򽪀��⋞�Ƞ����0�����+��   �   C3���,���=��Ǚ���;���Z��4v��Ʌ�g~��ʝ��S����ׄ���s�b X�9#9��7�i%���ӽ�?���8,Q�v�N�޽6����ӝ�[8��T�Ͻ��Z�4���l��3��ȅ���L�����-���_�'��8*��&���������8�ھ�����s����_��(�O����t���К������o��Z}ݽ���5�T��   �   #h�����C�f�?��1g�8����h��v������H��l ��J���;���n����d���=����n8�������8�vT��FĽLW��E<��f�o�սz_
�6�2���b�֋�H�������Oپ��L��<U���1��E辊6Ծ|�����u����R���"�h����ϸ��命|������R,��; �$�6�s耾�   �   ]�Ҿ�#���6��ad�n���9������nÿ`$Ϳ�IпV�̿;�¿g����8���㈿LGc��$6��	�S}Ӿ����[�	����ܽ�N��������,��,Tѽ'���~&�H�K��r��苾�M��� ��Ȱ��ײ�
뮾�S��j󖾄��d�b��:�H��������얃��^���c�7.��4�Ƚ����&V�/o���   �   ����"���R���������yo���Ͽ�����	����
��Eο�����?�������;S���#��W���|��]N}���0�#K�����b����O|��΅�|ߝ�,�½����
���,��F�-C\�HCm�ew�E�y�s~s�Q�e���P��N7�v��iB�� �Ž4핽b��4��$+�?�L��I����۽,�%���t��D���   �   |���D6���k�!�����<�Ϳ[������J��p���i����H�!MͿ���p��I�l���7���	��9Ⱦڽ���D��һ�j���y{c���Z�@q��ꎽ���p�Ͻ�����
�P��y�$�$+���+��'�S������*��,`ͽ$	����z���9�Y��P/�>���>��:��n��7������þ�   �   �"��kE��U����>��޿Q<���a�0M����:7��F��)���1޿����&۟�b����G���mپ����T�u���]Ž+ъ���T���:�,�>���W�{�~��ʖ��J��b�ƽ@gڽ.�轓{�7������׽C���ۤ�7i���O����8�ּR!��J���,�ۼ�g7��R��� ��!�D�������Ӿ�   �   FZ��O��ۅ����EIȿv�@������6����1����b�� ��ɿɧ�s����Q�TN�6z��e��p�^��9�z�˽L���J�L�v�(���!�^/�,J�O�k�������[��0���$F��A������ʧ��R�k��:���	�Ĕ��T0v��8��O[�Vk��f�3����Ј�A�M������ݾ�   �   ���@iR�M����T���b˿��&��8���t3�`��(-������gX̿�����P��LU�k���I辰���hb�?w�bJν	z��>J�x#����-"���8�_nV�d3v�B&��.����~���X��J����5��DL��>ew�.VM����� �����\:�4�
�D<����]�2��x���L���P��_��|w��   �   �Y��O� ۅ�_���}Hȿ5u迾��.��<6�F���0����ܣ�!��ɿ�ȧ������Q��M�=y�e��v�^�9�{�˽����)�L���(���!�v]/��J���k��t����[�����F����A������ç��D�k���:���	�z����/v�l8�N[��i��R�3����2��Z�M�]�����ݾ�   �   �!�jE��S�h���<��\�ݿ\:���`�L�|��6��E��'���/޿񸿿�ٟ�P���=�G����Ckپj����T� ���[Ž�ϊ�k~T���:���>���W�z�~�Nʖ��J���ƽ�fڽ���o{�h7����׽9���sۤ�$i����O������ּ  ��l���l�ۼ�e7�4Q��4���g�D�i���4�Ӿ�   �   ����B6���k�D������όͿ����������֮�Nh����>E濥JͿ���1n��N�l�<�7��	��6Ⱦ���U�D���dϻ�p���cxc�L�Z�Rq��鎽H����Ͻw���
�$��V�$��#+���+��'�M�����*��`ͽ
	��y�z�"�9�����,�<���>�g8��)��7�,���þ�   �   �	�.�"���R�f�������l��xϿr��R��;��%��z࿮Bο����R=��q����7S�ѧ#�cS��zy���I}��0��F��m�������K|�zͅ�Rޝ�.�½���
�]�,��F��B\�$Cm��dw�6�y�j~s�K�e���P��N7�o��LB����Ž�약 b���4�%"+���L�PG���۽J�%�_�t��A���   �   ��Ҿ!�ζ6�F]d������5��/ ���jÿO Ϳ�EпC�̿W�¿�󲿛5�������Bc�� 6����xӾ���ۇ[������ܽZK��n����������Rѽ���f~&���K���r��苾eM��� ��Ȱ�wײ�뮾�S��h󖾀��Y�b��:�0�����>�����{�^���c�D+��܌Ƚ���"V�l���   �   �c�����@���?�4,g���d��%r��夬�mD��D��S��W7��Ik����d�7�=����r2뾌~��6뀾*�8� Q��AĽ�S���9��Z���ս�^
���2���b��Ջ��G��_����Oپ���B��7U���1��F辋6Ծ|�����n����R�{�"�����ϸ�g䑽u�������'�� ���6�>倾�   �   /��M'���6��F��S�;�|�Z��-v��Ņ�fz������U����ӄ���s�X��9�_3�%���ͽ������%Q�jq���޽c���%Н��5��]�Ͻ����4��l��3�������L�����-���Z�'��8*��&���������8�ھ����vs��}�_���(�����xs���Κ�����k��)wݽp���T��   �   �g������ľ
����d�+�
yA��JR�W�\��"`�V�[��uP�l?�*)�֫��=ﾱT���5��s_��y$�$�{��@���hà���� ���ف+���g����i�ľ���(����+��{A��MR���\�B&`��[��yP��?�B)����3B�qX��y8��!_�g}$���~��8���Ġ���$���$�+��   �   u�4�խl�S1�������Hᾴ���*�<��N�'��5*���&�����L�����ھѵ��Mp��w�_�ϡ(�����Jo��̚�w��� k���wݽ�����T��0��c)��h9��"����;�I�Z�(1v��ǅ�Y|��Û��b����Մ�N�s��X�� 9��5�k"��_ѽ������)Q�4t�r�޽����4ѝ��5���Ͻa��   �   �\
���2�ٿb�jӋ��D������^Kپ`��K ��P���,��H��1Ծ�w��	��Q���h�R�]�"�z|��Bʸ�����(��u����'��z ���6�4怾7e�����{A���?��.g�^����f��t��馬��F��i��n���W9��"m���d��=���$6�a���Q퀾3�8�S�UDĽU���9��]﫽��ս�   �   Pѽ����{&�'�K��r�拾/J�����1İ�|Ӳ�箾�O���=����b��:�$����	��3�����^��c�J*��ŌȽ(��#V��l��\�Ҿ"�,�6�_d�Ű��47������lÿF"Ϳ�Gпa�̿m�¿����v7��_∿qEc�[#6���{Ӿ����[�ݪ���ܽM��􌏽,������   �   Mܝ��½j�����,�jF�=>\��=m�M_w�W�y��xs��e�m�P��I7�$���:��őŽ�畽*�a�o�4��+���L�vF��ޏ۽��%�(�t��B���
��"���R�,��������m���Ͽ����#����l࿏Dοy����>��ҙ��L:S���#�JV���{��%M}��0��I��8�������K|�u̅��   �   �q��玽V����Ͻ����
�ڹ���$� +���+�n�&�P��3���#���Yͽ�����z���9�����#�}8��>��7�����,7�\��x�þ&��C6�m�k����������Ϳ���H���v�����$i�3���F�,LͿ2��mo��g�l���7�H�	��8Ⱦ~���m�D��>ѻ�`����xc�D�Z��   �   v�>�(�W���~��ǖ��G����ƽ�bڽr�轊v�L2���֊׽l���פ�.e����O����Z�ּ���������ۼ�c7�HP������%�D�X���;�Ӿ�!�FjE�>T�����<����ݿ;��Pa��L����6��F��(��'1޿����ڟ�.�����G�����lپ������T�n���]Ž�Њ�KT���:��   �   ��!��\/�]J�
�k��퇽�����Y������C���봽�>��&���W�����k���:���	�ʍ���#v�8��D[��e��5�3���������M�����Z�ݾkY��O�ۅ�T����HȿSu�܄�\��|6����D1�`��B������ɿ�ɧ������Q��N��z�f����^�$:���˽����_�L�%�(��   �   �6��<��J���[���l��{���9��f���$O|�5:i�C_N�b�,�0��쾽�x�`�h곻 ��9@?<;���9���ռ,^��[Ľ0���o�:����G�F�"��BS����"4���@��	Hп@k�4�u��~���п����៿e���f�U�ս%��M��z�����æ8����hʸ�~�����X��=��   �   �<�,F��`W�,�k�:���6��֏��(���z���_��@����kk�FH��T3�������`�(� �:����e��ؼW\�c������y/l�R���v�VS ���O��������nb���Ϳ��޿�U�5AN�}�޿�7Ϳ1���P���̂�
R�} #��.���y������%�5�����L_��0���kY���@��   �   i�O���b���}�|������0���\��@T�����f��>���G3�������j���6���4��A���ӻ8˻��M�0�߼�W�Ip��7���a�8���a�g���0F���w�=~������ÿ�Կ��߿�?�Pr߿�Կ+�ÿ'���ו��	y�s�G���2;龝Ū���t��-��?������4ׄ�9�[��YK��   �   �q��.���s��`#��yҽO
齴)�����������7��a�D\ս�>���_����d���%� 5�N+����p�.m��x�ＧbQ��r��G�
�2Q���� Ҿ����6���d��!���ᠿ:�����Ŀ��ο�	ҿ�wο�XĿ)��������%��6fe���7������־�5���a���Z��n����i����a� �^��   �   m����k��RJҽ=l�������!��B1�G�<���B��C���<���0����H�
�����������M�I���o޼�Ѽ٠��TL�(l��<@��0�<�@���f9��v��'�#��L��-w����k��D.�����$���и����~�������}v��mL�{�#�����z������!I�����'ͽL���gt}�0n�D�}��   �   ��O�w�d�'�^�D��`���w�R��9a��FU��к�����bqh�q�K�ri,��E��d۽���sr�<4�ʇ��j��K��A���pཐ�%���l����3۾���6G1��V��y�T����Ƙ�󇠿F��*���!��g���	x��T�v50���ڹھX���_q���-����\ϵ�z���|��݁�ೕ��   �   ��h��3�8���`�\*�����r����!��\��k¾{���}��Σ��^����u�	�I����(p������6%���EP��;��$P�։�pŽ~>�|[I�C{������'L�����3��[Q�<�k��*�������È�tC����~���i�<O��|1������6�� ��c?I�1H��lҽ����h!���ꁽ�ǒ��n���   �   ����>�PKq��o���0����̾���f���J����X>����Z�߾��ž$���������]���*������I��?����e�Z�]�����L������̘'���d��t��,�¾�_�:��7*�bN?�(�O��yZ�)�]�?�Y�TN�8=�Za'��1���쾅l��KĒ�c�\�."����n5������f�~���*̪���޽�   �   ��8��r��������G}�X���e�)S#�Kl+�P�-�vy*��~!�Z�����Hp߾����D���dGd�+��!��V��P�#�t��6|�����4Aʽ�D	�y�8���r������)y����Zc�[P#�fi+�n�-��v*�|!�
������l߾񔸾'���3Dd��|+����T��U����t�o8|��Ø�xDʽ"G	��   �   f�d�Iw��_�¾�c����*�XQ?�Q�O�}Z�\�]�R�Y��VN��=��c'�Z3�����n��ƒ���\��/"���뽞6��@���'�~�|}���ɪ���޽V���>��Fq��l��4-����̾#�徧����G�Z���;�����c�߾2�žB��������]��*������F���󌽇�e��]�(�����t�𽎛'��   �   V}��c����O�4��3�3�z^Q�c�k�n,��p���=ň�E����~�4�i�]>O��~1����&뾲8��W!��&AI�RI��mҽR���!��h遽�Œ��k�����z��p�8���`��'�����╪�'��$X��g¾�����y���ʣ��[��Ȧu�(�I����tk��L����"��CP��;��%P��׉�:Ž�@��^I��   �   G���۾���iI1�]V�ʣy�邌��Ș���������+��5#������Hx��T��60�����ھ�����`q���-�6����ϵ��y��e�|��ہ�j���� ���	�t�ȸ'��D��`�	�w�\��&^��2R��Է��,��Ulh��K��e,�qB��_۽���r��4�����j�.K��C���s�ԍ%��l��   �   �;��My���#�6�L�o0w�]	������/�� ������Ѹ�^���9������Xv��nL�p�#�`���u��@���"I�_���'ͽ(���$s}��n�{�}�Ϡ��9h���Eҽ�f��k��ٶ!��>1��<�c�B�^C�F�<���0������
���J�� ��C�M�C���j޼�ѼE���VL�n��WC��u�<�ך���   �   Ҿ��6���d��"��㠿����H�Ŀ�οҿ�xο�YĿ�������q&��%ge�T�7�����־�5����a�J��z��6���i����a�_�^�D�q�R,���p�������ѽ��#����x��P��p4��[��Vս(:���[���d��~%�-��%����p��l�� ���dQ��t����
�@4Q����   �   �c�|���1F�x�w�������ÿ�Կ��߿�@�!s߿ÏԿ��ÿ�'���ו�d
y���G��g;龳Ū���t��-�f?��G����ք���[��WK���O��b���}�xy�����{-���X��NP�����V
��L����/��D���9�j���6�w{������@���ӻ�˻��M���߼h�W�r��p8���a�d9���   �   5x�%T ���O���������c���Ϳ_�޿@V꿱A��N���޿�7ͿN���P���̂��	R�Z #�j.��{y��j�����5������^�������iY��@�<�<�*F�]^W�T�k�}8���4��6ԏ��&���x���]��Z���Mhk�4H��|�/鼚������@�(�@�:����4i��ؼ^Y\���������0l�V���   �   �H���"�hCS����l4���@��CHпkk�K�s����}�ƃп˳���៿���؋U�Y�%��L��py�������8�B��jɸ�����a�X��=� �6�%�<�F�J���[��l�t�{�����H���O|�N:i��_N���,����&���<�`��� ,�9p0<;�u�9@��D�ռ.^�]Ľ�0���o�龭��   �   6w�{S ��O��������Vb���Ϳ|�޿PU꿼@��M���޿�6Ϳ����oO��ĵ�	R���"�]-���x��ژ���5������]��Ѝ��^hY���@�W�<�)F��]W���k�.8���4���ӏ��&���x���]��E���1hk�H�_|��.�f���`��p�(���: x���f�ؼ�W\��������/l�����   �   �a�8��D0F�r�w��}��\��U�ÿg�Կ�߿�>�Wq߿�Կ,�ÿ&���֕�Ny��G���h9�:Ī�t�t�-�=��x���8Մ�Q�[��UK���O�}�b�M�}��x����� -���X���O�����!
��*���|/��0����j���6�?{�L��\�@�@�ӻ�˻ܰM��߼ՁW�6p��7���a�8���   �   zҾT���6���d�!��ᠿU��Ŀu�ο�ҿZvο�WĿ࠴������$��Bde���7�/��՛־�3����a���2�⽲���g��o�a�s�^���q�2+���o������ѽp�c#��ʼ�L��0��X4��[��Vս:���[��֥d�+~%�
,�`$���p�i��N��CaQ�r����
��1Q�!���   �   e8��u��5�#�װL�f,w���K���,��'�����ϸ������|��$���={v�kL���#�	���,�����"I����$ͽݙ�Dn}��n��}�J����f���Dҽ�e����t�!�g>1���<�3�B�<C�,�<���0������
�˶� �������M�`��2h޼��ѼO��?RL��j���>��.�<������   �   ݲ���۾۽��E1��V���y�����Ř�c������\(�� ��е��$x�w�T�430���ضھ����o[q�۩-�q���}˵�xv���|��ف��������B�ss�1�'���D��`���w�<��^��R��ȷ����Glh���K��e,�\B��_۽���r�=4�����g�ZK�@���n�>�%��l��   �   �y��ҙ���I����3�OYQ���k�G)��"��������A��j�~�d�i�+9O�mz1����#�4������;I�ZE�hҽ��������恽HÒ��i��֧罸���8�I�`�U'�����������X���f¾�����y���ʣ��[����u��I����'k��̣��,"���@P���:�� P��Ӊ�Ž�<�}YI��   �   ݄d��r��ʪ¾�\�[����)��K?�M�O��vZ���]��Y��PN�>=��^'�/����&i�������\��*"����0��鱊�q�~��z��OǪ��޽���j�>�Fq�ml���,���̾��後����G�U���;�����`�߾-�ž<�������͐]���*����F��x�I�e��]���������n�𽷖'��   �   Ρ8��r�����A����u����a��M#��f+���-��s*�Fy!�d��V���h߾\���.}��b?d��x+�s��B���덽
�t�P0|����0?ʽ�C	���8��r���������x����Jc�OP#�_i+�j�-��v*�|!�������l߾씸����Dd��|+����V�����t��1|�𾘽>ʽ�B	��   �   �����>��Bq�<j��5*��%�̾��0���*E�����9�܏���߾~ž��������Ӌ]���*�ڹ��LA���j�e�#�]����������'���d��t���¾^_�%��(*�VN?�$�O��yZ�(�]�>�Y�TN�9=�[a'��1����|l��=Ē�5�\��-"����4�������~��z��zƪ�&�޽�   �   @��Ǐ�}8���`�%�����������>T�� c¾����v��3ǣ�|X����u�.�I�����d������4���:P���:�WP��Ӊ��Ž�=��ZI��z��j����K������3��[Q�3�k��*�������È�uC����~���i�<O��|1� �����6��  ��-?I��G��kҽA������災��Uh���   �   ���?�Zq�j�'��D�P`���w�~��[��O���������fh���K� a,�|>�$Y۽x����q��4��~�?d�tK��?��Do���%�3�l�泣�۾��(G1��V�ܠy�R����Ƙ�􇠿G��*���!��h���	x��T�v50���ѹھK����^q�o�-�&���ε�x��s�|��ف������   �    ����d���Aҽ�a��Y��S�!��:1���<���B��C���<��0�z���
����8�����s�M�ȳ��]޼6�Ѽ����PL��j��?����<����=9��^v���#��L��-w����k��F.�����&���и����~�������}v��mL�y�#�����r������!I�����&ͽ�ޙ�p}�n���}��   �   .�q��)���m�������ѽ �V�����@���� 1�wU��Pս�4���V��N�d��v%��ἂ����p�c��ҒＺ_Q��q����
��1Q�m��Ҿ��x�6���d��!���ᠿ;�����Ŀ��ο�	ҿ�wο�XĿ-��������%��6fe���7�����־�5���a�������Z���h��:�a�(�^��   �   A�O�	�b���}�w�����V*��wU��vL����� �����w+��Z�����j�8�6��u�r��p�@��sӻ��ʻP�M��߼4�W��o���6���a�8���a�_���0F���w�;~������ÿ�Կ��߿�?�Qr߿�Կ,�ÿ'���ו��	y�s�G���.;龖Ū�z�t��-�>?������3ք�]�[��UK��   �   |�<��(F��\W�h�k�M7��x3���ҏ�0%���v���[��I���0dk�4
H��x� (�.���<�� �(��d:�9��l_�vؼ5V\�
������^/l�F���v�RS ���O��������mb���Ϳ��޿�U�7AN��޿�7Ϳ0���P���̂�
R�~ #��.���y�������5������^�������iY���@��   �   (��*?��
���9���߅�!�����u0r���`�ʴJ��0�t�Dݼ��������@>�;l4<,]U<T�3< Mm;@�*�9���x����㽆�0�+��z´�P��[4��TF���o�8��^˝�H̫�S���Yշ�m����׫�o󝿦T��i�p�'�G�k� �?O��,#������eQ��1�:��r)��4嚽҈��{���   �   �<������ 爽�p��L����ˋ��ۈ��|��w�l�a��G�<h'������d[\�(����C;�)<6<<��4;8�0�;���˄�\�཈.�Sl~�����������,C��l�
ʉ�xM�����9屿R괿�߱�f���g��b��m���D�����(������>h��B�M�i����2g��l��^���h����   �   �F��bm������~���|��Q���Д��}a��&����#��>φ��k���C�\0��QּDG��X˻ -�:`��;Xɰ; ��8��B�l��\���o׽��&�	s��ܩ�X�侂j��:�g a��W�����k0��D����m��������x���n����a�&;��;�v꾜ٱ����7�C��1�>ܽ�����
��Hl��#Z���   �   �"��Ɗ��ƹ����,(ŽTнF�׽/�ڽ��ؽ�Wѽ��ýl簽�N��@�|�0VD�������8�=���Y�p#��8tf�`���or��[ɽ'��z�a�HJ��OYӾ�	�z�+�4�O�{r�W���:Δ�7���>"���a��-����m��n*r���O��3,�6
�@\׾.���j�s��4�Ւ��%˽v���~֌��ʄ�⨆��   �   �b��Ҷ����ɽF��i%��o�8�_��L{����g�H�����Ƚ ����{�.
6�tP��j\����H�0
=�����u�i	c��=���u��K�:��������������9�7�X�Qt�k���ዿ�*��&�������$as���W� �8��H������������X�� ��������������TG�����   �   ~갽$ҽug��.p��#�8G5�j�D�T�O��U��LT���L�"Z?��,�����=��xȽ����S�]�
0���׼����b=�� R��U��:���a���D3���w�[m���վJ�B� �F�;�kS�8f�5�q�,�u�gWq�e�� R�:��[�����Ӿ�٤��Cz��J:��g	��̽۞�FЅ��2|�֋��.S���   �   ouνq��\�>b7�'�T�X�p��?��aE��{f�����&�Bl���Ct�L:V�&5��z�
�潞����#|��=5�y%
��u��P���LK�l��-ڽ����'T�L����������"C�;x�n31�t�@��yJ�R�M��I�KE?�T?/�l'�s����۾�(��L��6�O�wX�܏㽘��������p��s��'�����   �   :���-�}�A�kYj�D�+՝��E��ѱ����ľb�ƾR���p�������+���z���M�3#������m���E��2�I�&�&��%�6H�������MU2�:Kj��P�����+ݾ�L ���YV��$�Ug&�>#����+r��8����վV㰾ؚ����[�5!&������i�������e�[�D6s��O��P���   �   �I��@�7r��N��om����˾���V8��r� �}�"s�����I�ܾ�*þ����|��w[���)�����w��������X�7=A�!OM��C|�읦��߽�G��@�8r�L��mj���˾�+4��H� ��z��n�������ܾ�'þ�����z���s[�@�)����jt��᪊�v�X��<A��OM��E|�	����߽�   �   �W2��Nj�AS��䙸�~.ݾ�N ����X�J$��i&��!#�ψ�t�2<��O�վ�尾����3�[�-#&�u���xk�������e��[��4s��M���M��D6��p+�/�A�FUj��Fҝ��B��P�����ľ��ƾ����%������5)���{z�	�M�A0#�+���Lj��xC��*�I���&���%�y7H�����,����   �   �*T�I���.�����E�az��51���@�0|J��M���I��G?�UA/�')�����۾�*�����1�O��Y�ב�ަ������7�p�.�s�j&�����rνm��}Y��^7�'�T��|p�=���B���c�����J񎾔i���>t�
6V�n"5��w�D��ꔭ�O|��95�#
��s������NK��m���/ڽú��   �   �w�ro����վ�K�2� �x�;��mS��f���q���u��Yq�Le��R��:�]�9��T�Ӿ�ڤ�ZEz�<L:�oh	�7�̽�۞��Ѕ�22|�����Q��R谽ҽjc���m��#��C5�b�D���O�U�
HT��L��U?�?�,�x���7���Ƚ&���Y�]��+�z�׼�~���<���R�	U��<���d���F3��   �   ̀��Ĥ����������9�P�X�MSt�����8⋿�+��A��������bs�k�W�Z�8��I�D�����������X�� ���	��3��������F����Xa��������ɽ���� ��Tl�8����w�������.���Ƚ����L�{�L6�>G���U���H��=�̿��cv�"c��?��xw�9�K��   �   �K��8[Ӿ�	��+�ްO��|r�T���>ϔ�;���9#���b������qn���+r���O�V4,��6
��\׾�����s�4���&˽����f֌�:ʄ�0����!��1������������$Ž�н�׽��ڽ�ؽ�Rѽ��ý�ⰽ�J����|��OD�^��>��p�=��ݓ�`-� ��8vf����Zrr��]ɽ�����a��   �   ީ���侂k�
:��a�]X��M��21������n��]���|�����o��I�a��;��;����ٱ�0���I�C��1�6ܽ�����
���k���Y��F��Sl����������Z��ޣ������^������ ��:̆�g�k���C��+�Jּ�:��D˻�g�:���;�Ͱ; ��8d�B�(������q׽��&��s��   �   �����ﾤ���-C��l��ʉ��M��B���屿�괿B౿����g��w��m���D����f(������h����M���H��f���������A<�����*戽�o�����Aʋ�ڈ�X{���w�[�a��G��e'�����	���T\�`��0�C;�+<�6<D<�4;̉0�����̄��ཬ.��m~��   �   ô����4��TF�T�o�l���˝�i̫�d���Zշ�]����׫�C�sT����p���G� � ��N���"��F���FdQ��0�>�꽫(���䚽T����z������>�����L9��`߅�ڵ��<�0r�O�`���J��0����Dݼꊔ����@���8�;(i4<ZU<��3<�;m;t�*�Й��y��-��Z�0��+���   �   ����������,C��l��ɉ�SM������䱿�鴿�߱����?g�����m���D����W'������pg����M�i����e��8��7���<����;��r����刽^o�������ɋ��و�{���w�	�a�YG�Ze'�h���	��<T\������C;�,<�6<�<��4;Ć0�׽�7̄����.��l~��   �   �ܩ���Ej�:���`�JW�����/������+m���~��)��� ���m��c�a��;��:���@ر������C�h0�ܽ�������~j��AX���D�� k��x�������v�����r���^������� ���ˆ��k�g�C��+��Iּ\9��B˻�r�:���;HӰ; ��8��B���9���o׽|�&��s��   �   �I���XӾ=	�Ʒ+�L�O��yr�����l͔�Q���E!���`��&����l���(r���O�$2,��4
�8Z׾������s��4�8���"˽���(Ԍ�2Ȅ�L����������%���r����#Ž�н$�׽��ڽ��ؽCRѽ��ý�ⰽ`J����|��OD���x����=��ד� � ��Xnf���,nr��Zɽ�����a��   �   l~������~�������9���X�HOt�l����ߋ��)�����������^s���W�:�8�=G������'���)�X�� �L��������.�\D�����>_��������ɽ���Z���k�������w�N���������꽢Ƚ�����{��6�4F��FT��t�H�h�<�����r�c�G<���t���K��   �   ��w�l��'�վ�H��� ���;�%iS�f���q���u��Tq���d�6�Q��:��Y�j��ʮӾFפ��?z�H:�1e	�(�̽�מ�ͅ�=,|�]���HO�� 氽��ѽna���l��#��B5�ԔD���O��U��GT���L��U?�$�,�\���7��{Ƚ鞘���]��*���׼�z��07��O�rU��8��l_��C3��   �   T%T�ٰ��ð����ྪA�{v�h11�.�@�$wJ�M���I��B?��</�8%����l�۾&������O��U�.�㽥�������%�p�	�s��#������,pν�j���X�
^7�\�T�|p��<��ZB��bc�����3񎾃i���>t��5V�V"5��w��潘���q|��85�2!
�Vn�����IK��i��U*ڽ���   �   S2�HHj�O������.(ݾ%K ���,T��$��d&��#�D���o��4����վ?ాF���X�[��&�&��� e��������d��	[��.s�MK��K��4��f*�<�A�iTj�f�ѝ�KB�������ľ��ƾ����������*)���{z���M�%0#������i���B��W�I��&��%��1H������뽽L���   �   mE��
@��r��I���g����˾2��70��,� ��x��j��q����ܾ$þ]���,x��Qo[�}�)�ß��`o�������X�|5A��HM�	>|�s�����߽�F��@�_r��K��j��Ԋ˾���4��:� ��z��n�������ܾ�'þ�����z���s[� �)������s������X��8A��JM��>|�����I�߽�   �   	2���(���A�ZQj�o퉾�ϝ�u?��몼�D�ľ��ƾ������R���&��Avz�W�M�R,#������d���>��b�I��|&�&�%�R0H�����g콽��kT2�kJj��P�������*ݾ�L ���JV��$�Pg&�:#����(r��8����վN㰾͚��i�[�!&�����h��������d��[��/s�%K��J���   �   �nνrh���V��[7�0�T�$xp�v:���?���`�����<�f��k9t��0V��5�t����`���|�25�0
�g��R���GK��i��'+ڽƷ��&T�����X������C�&x�`31�k�@��yJ�P�M��I�IE?�S?/�k'�q����۾�(��?���O�FX�B�㽱���¶��*�p���s��#�������   �   
尽2�ѽ�^���j�V#��?5�K�D���O�VU�8CT�>�L�JQ?��{,�x���0��{Ƚљ��R{]��#�H�׼�r�� 1��M��U��8��<`���C3�C�w�m����վ�I�0� �8�;�kS�3f�4�q�,�u�iWq�e�� R�:��[�����Ӿ�٤�hCz��J:�Ig	�R�̽�ٞ��΅�;.|�Ĉ��O���   �   �^��p����ɽ"������i�����Vt����n
�����}꽲Ƚ:�����{���5��8���I��0�H���<����8q�:c�L<��<u�g�K� ������ˉ��v���9�/�X�Qt�j���ዿ�*��)�������%as���W� �8��H���������㆑���X�� �a��2��Đ��J����D������   �   �������촩�����B!Žtн��׽��ڽ�ؽ�Mѽ��ý�ݰ��E��"�|��GD�Q}��	��Ċ=�ط�����  ��ff����?mr��Zɽ����a�J��/YӾ�	�m�+�,�O�{r�V���9Δ�8���?"���a��/����m��o*r���O��3,�6
�:\׾'���S�s�p4����*%˽����BՌ��Ȅ������   �   �D���j��Ԯ������
��D���:���v[��֝������Ȇ��k���C��%�`?ּp'�#˻ �:�Ю;��; ��8��B�������5o׽R�&��s��ܩ�C��yj��:�c a��W�����l0��E����m��������y���n����a�$;��;�r꾘ٱ�����C��1��ܽ����	��0k���X���   �   �;��~���t刽o�� ���ɋ��؈��y����v�%�a�TG�Ib'�a�����hI\������D;�4<L&6<<<��4;؀0�Z��f˄�
��c.�4l~�����������,C��l�	ʉ�xM�����:屿R괿�߱�g���g��b��m���D�����(������:h��5�M�[�����f����ԫ�������   �   ��ʽ��ɽCEŽ%)��̟��^M���璽F��K�\��y6�m��(_м�R�� mۻ@��:��<d�<8{�<:!�<=�<�1c<0�/;��t��L%�Z��������8�_L��.�{�������-��zK���e�c�z�����B������:�z��f��L��/�����.�_���	D��Mw_�*./�!��\��ؽ�̽?]ɽ��ɽ�   �   F�ɽ8�ɽ�\ƽPx��{6���&��L꘽����Jl���F�T5 �tM�\ơ���'��������;L~X<<O�<8�<h|�<@�U< �;Lu���#�L0���;��V6��b��C��o?�;N��-+��8H��b���v��ց�C���ҁ�Γv��Gb�0�H��4,��$�aE羷����܍���[��8,�y:��S��Խ�ɽ��ƽ�
Ƚ�   �   =Dǽ�ʽRʽL�ƽ�|��/9���|������獽y��MS���*��� �����<�4� ��(,�;��B<8cx<��u<x�,< W:�Az�O��Ⓗ��*�.�4�u������־i���(#�s�>�gfW���j�QLw���{�a-w�Q�j��PW�s�>�E�#�z"�Y�۾܎��f�����P�	�#�o<�L���ʽ�:�����0ý�   �   ڛĽ$:̽�ѽ��Խ-�Խ=ҽG>̽�Xý�R���'��敽�Ԁ�(S�k1"�jV�$���P�ͻ`U�:P��; W<�;`��󃼖��+���fݽ�e#�G�d�T��� (Ǿ<�����0��F�ӊX���c�8�g���c��X��3F��/����Nm���Bʾϔ��?�w���?�����_ν�.�����R(�������   �   ʶý&ҽ��߽P{�����k��!���������������&׽J���P���2B���~S�@��ü@Q��`�� $c� m�кƻXy������t���>̽c�#�O�n���8Y��v�߾� ��z�n�1�9RA�_aK�ĲN���J�6�@�"�0��f���~�޾�޳��֍�g\�1�)�`���ֽA]���1���>��䪽��   �   ��ƽ�8޽u)��_��.w�+���f!��%���$�Ƹ ��'�.��|!��vҽ�����̈́�w|A�L��j��x�I�����G�4��	!���t���*_��9�u�3u���}þ8����-��]3'���/��j2��/��%���Ϋ���澧���l�����s�7�<�~6�|O⽂���������r��PW��͑���   �   нԯ����0���1���A�a�O���X�1�\�U�Z��KR�ٷC�R0����sW��ĵ̽���&
f���!�<⼞m������`�Ӽh�&4i��p��p��Z�"��!U�[���¦��?Ǿ���P�A����'��,��t
�����`Y྘���S���Y����I�(��`J����������,�~�E���y�� q���   �   %���/�"�i�>��gZ�\]t�RI����������K������Sq���S�3��(��彾���Tۀ��<��V���������(���d����~�ֽ�=��7��He����-D�������Ӿ��侑��񾯉�v�߾=�̾ӿ��<���#��SRM��s ����)��� C����k�x�U�:tZ���w��锽d(���   �   �����J��@�Hg��冾�Z��Ew���ǵ����Jr��I���"��U����ǌ��o�N�E�������;��R��y[T��81���)��)=��zi�0���ܜý���I�t�@��g��ㆾOX���t���ĵ�n
��6o��O���K��Ӳ���Ō�T�o�B�E�?�����8����XT�961�\�)��(=�B{i������ý�   �   @?�6!7��Ke������F�������Ӿ��
�y���쾑�߾�̾=´�C���p���TM��u �(��������D��;l�b�U�LuZ�ӏw�锽8'��%�b���"���>�XdZ�fYt�G��}���L��š��Q����Oq���S��3��%����R����؀��<�	T���������(���d������ֽ�   �   J�"�h$U��\��Ŧ�hBǾ��澾Q��B����)��.�=v
������[ྴ��`U��H[����I�����L���\�������~�����y��qp���н���8����31�t�A�̅O���X��\�"�Z��GR���C��0����R��E�̽B���Of�r�!�v��h��ȡ��p�Ӽ�h�
6i�Lr��$���   �   �9���u�	w��B�þ�뾘�����35'���/�kl2��/���%�)������G��������s���<��7�6Q���1���[���Bs��zW��������ƽ7޽.'��ո�4u�Ǚ�:d!��%�M�$�~� �e$� �����
qҽ2�� ʄ��vA��	�rc��ȩI����LG�Z��&"�^�t�����`��   �   H�O�����[����߾(�p|��1��SA�#cK��N�;�J���@�o�0��g�����޾�߳��׍�� \� *���@�ֽ7^���2�� ?��d䪽�R�ý%ҽ�߽y�!���������n���)�������!׽�~��	���e>��xS�����ü�Q� K�� 7a����8�ƻnz��C��"v��A̽�d��   �   P�d������)Ǿ>�����0���F�S�X�,�c���g�P�c��X��4F�Ƶ/�H��Zn���Cʾa����w�@�?���،�~`ν/������(��у����Ľ�9̽��ѽ]�Խ/�Խ�ҽj;̽�UýXO��$���╽�р�"S�,"�
M������ͻ@��:8��;�[<0!�;`��J���W��v,��
iݽ@g#��   �   ��u������ ׾B���)#���>��gW���j�oMw���{�S.w�"�j�kQW���>���#��"���۾���������P�4�#��<����7�ʽ�:����0ýDǽ�ʽ�ʽW�ƽ�{���7���z�������䍽�y�vIS���*��� �▬�X�4��Q��;�;��B<gx<��u<��,<��V:HFz�+��r㒽�뽄�.��   �   ^c���C��}@��N�_.+�r9H�Xb�:�v�)ׁ�����ҁ�$�v��Gb�R�H��4,��$�IE羘���f܍�^�[�]8,�R:��S�ɉԽ�ɽt�ƽr
Ƚ�ɽ�ɽ#\ƽ�w���5���%��Q阽���`Hl���F�(3 �|I��¡���'� z����;4�X<$P�<r8�<&|�<��U<��;`�u���#��1��a=��W6��   �   �L������N���-��zK���e���z�,����B�������z�Hf�kL��/�S���-�ؚ���C���v_��-/����`[�Vؽz�̽�\ɽE�ɽ��ʽi�ɽ�DŽ�(������M���璽���\�{y6�j��T_мtS��Poۻ���:�<X�<(z�<��<�;�<<.c<p�/;��t�]N%�\�������8��   �   �b��-C���?�@N��-+��8H�gb�4�v��ց����Fҁ��v��Fb�w�H�4,�H$�ID�̓���ۍ�d�[��7,��9��R콺�Խ��ɽs�ƽs	Ƚ#�ɽ�ɽK[ƽ�v��5��%���蘽d���Gl��F��2 ��H�F¡���'��t����;�X<�P�<�8�<�|�<0�U<��;�u���#��0��4<��NV6��   �   ��u�Z�����־"��@(#���>��eW��j�aKw�}�{�B,w�*�j��OW�\�>�E�#��!���۾����`߆�!�P���#�M;�U��"�ʽ�8�� ��'.ýFBǽ�ʽʽ��ƽDz��n6���y��Ĝ��H䍽�y��HS��*��� �"����4��G�8>�;��B<�hx<�u<��,<�BW:�?z�ը��ᒽε���.��   �   d�d�����2'Ǿ�:��9���0��F���X�T�c���g�s�c�X�f2F���/�Z��k��AʾM�����w���?�r�K��V]ν6,��X}���%��,����Ľ7̽��ѽD�ԽN�Խ1ҽ:̽�TýsN��b#��
╽р�Z!S�|+"�&L�V���0�ͻ ��:���;$_<�*�;�g������.*���eݽe#��   �   ��O�����X���߾����y� �1��PA��_K�
�N���J�s�@�r~0�e�^��޾�ܳ�5Ս��\���)�����ֽfZ��+/���;��&᪽�뵽E�ý."ҽ`�߽�v��������n������������F!׽.~������>���wS�3���ü�Q�HE�� 7`��,�بƻ�t��P��is��6=̽b��   �   9���u��s��C|þ��Ƭ�����1'��/��h2��/�-�%���+�����%���Q�����s�b�<�*4��K������~����o���S�������ƽ�3޽0$��t���s����Xc!��%���$�� �$�ވ�{���pҽ�~���Ʉ��uA����a��t�I����xG�>����X�t��|���]��   �   m�"�^U��Y������=Ǿ�澋N�^?���%�+��r
�}��'V����:Q���W��"�I�X���E�����p���������~����$v���l��:н_��������1�i�A��O��X�z�\���Z�)GR���C��0�����Q����̽�����f���!�>⼾e��f���B�Ӽ=d��/i��m��X���   �   �;�g7��Ee�+����A����	�Ӿ����j������߾�~̾Ҽ��������tNM�up ���������@?����k�׎U�{mZ�{�w��唽�#����ҙ���"�b�>�.cZ�hXt��F���|����������6���dOq���S��3��%���� ���C؀��<��R�Z�������(���d����%�ֽ�   �   ����F���@�qg��ᆾ�U���q������O���k�����(��௟�����o�%�E�������3������PT��/1���)�>"=��si�橖���ý�����G�%�@��
g�Uㆾ�W��4t��Mĵ�7
��o��0���5��²��tŌ�;�o�'�E�!��v��C8������VT�D41���)� %=��ui�D���o�ý�   �   -���]�"�~�>��`Z�.Ut��D���z��W�
�������턾�Jq�$�S��3�^"����&���LԀ�v�<�MM�������M(���d������ֽA<��7�sGe������C��������Ӿ���h���񾗉�f�߾0�̾ʿ��0���	��8RM��s ����������B����k��U��pZ���w�4攽�#���   �   �н_�����B���1���A�ӁO���X���\���Z��BR���C��0����BK��N�̽���y�e���!�P��\��T�����Ӽwb��.i�n����<�"�� U��Z���¦�n?Ǿ`���O��@����'��,��t
�����YYྑ���S���Y��o�I���J�:���:��򆃽0�~�2��w��Hm���   �   ��ƽU3޽�"��n���r�і��`!�?%���$�ѱ �� ����6���jҽ�y��"ń�nA�C��V��L�I������F����a���t�}��4^��9���u��t���}þ�������N3'���/��j2��/��%���˫���澠���c����s��<�X6�O��ﶽN���Z���q��U�������   �   ��ý"ҽ��߽>u�����@��������������N׽>y����9���oS��t�üh�P�("�� �\����h�ƻNq����s��L=̽Xb�v�O�����X��<�߾� ��z�`�1�2RA�]aK�²N���J�6�@�$�0��f���y�޾�޳��֍�S\��)�7����ֽ�\��1��G=��O⪽U쵽�   �   ��Ľ?7̽d�ѽ{�Խ
�Խ`ҽ�7̽�QýTK�� ���ޕ��̀��S�%"�j@��x��Hxͻ 5�:���;`j<0=�;�)�탼���)���eݽ7e#���d�����'Ǿ�;��ٲ�~0��F�ΊX���c�9�g���c��X��3F��/����Jm���Bʾʔ��0�w���?����b_ν�-���~��'������   �   �Bǽʽ�ʽz�ƽ�y��i5���x�����Z⍽fy�7DS���*�� �����`�4����W�;��B< rx<l�u< �,<@�W::z����Hᒽ`����.���u�w�����־]���(#�n�>�dfW���j�QLw���{�b-w�R�j��PW�t�>�F�#�x"�W�۾ڎ��`�����P���#�V<��ག�ʽ
:�����.ý�   �   ��ɽL�ɽp[ƽ�v���4���$��:蘽����El��F��0 �hD�̽����'��0��x�;�X<�S�<�;�<��<H�U<� ;�{u�&�#��/��b;���U6��b���B��b?�6N��-+��8H��b���v��ց�C���ҁ�Гv��Gb�2�H��4,��$�`E羶����܍���[��8,�l:��S콿�ԽӴɽ!�ƽ
Ƚ�   �   ��!�/��Rn��V�`&���n�Ľ�^��JĂ�լG��� ���,t"���:8<@Y�<�)�<��<��<�l�<��<L>R<��n��f���?���o��Ą5��'v�H0���Ⱦ�w�q�3� �n�/��9��W<��9��/��C!��7�x�����ξLϩ�"≾�`���:���!�z�������R��������   �   O���%��j����+O��=�1�ǽT&���`���R����iȼ(�N����ȁ�;��u<��<���<BD�<��<R�<�.H< ʩ�(E���>��e�������@3���r��坾�ž>��y3�f���,�t6��B9�
6�p�,����������O]˾��������i�\���7�L��]$��=����<��#������   �   �u�������|�����{��Iн����ﮕ�/r�\5;�\��Q��$!� f�8 �<�|<�x�<���<*�<���<l^(<�c'�h٫���;��1�����W�,��Ji��M���U��X��{�����К$�&Z-�"R0�69-�pi$�4�������澺]��J���
ـ���Q�A.������	�K2���������|��   �   ���������6F�b������TȽ<���C��ޘv���B�Y���V���DG�@D��!�;�0F<���<<��<0
a<���; 1������<{9��n�����c#�~�Z�):����
=Ծ/m���l�Y������g"�/y�!N�,�
��c���!ԾǱ�䑾ٮl��j@����
��C��U��x����V�4��Z��   �   X�	�|��r�����(
����+����_�Z�սvw��dY�������4e��.�x�������������9 ��;��<���; O�:��� hƼ��9�<�����ڽI���BI�>܀�ؠ��}{���b޾����	��
�����h��������4۾�������a�����Q��N*����h�=�޽XGؽR�ܽb������yx��   �   �
�\h�������\F�S�z��>q�*����������ɽ$;��T����[���l�Ҽ(�t���P,���� [Ż@�m�j�伬�>�FĐ�(νz����6��!g�����������¾.�پ���N��l`���D���J���Ծ䧼�]8�������%^��t3�y�&Xｑν�����������jt̽��ݽ����   �   |j��t����j�	""�.N(�c,��,�w<*�\�#�̛�D���t�� cѽ�ڪ��K���F�����C�����	b���*�����	��bK�b����Ľ���r%�2ZM��x� ����Ȧ��*���`Ǿ��Ͼ
Ҿ�<;m����g������ˆ�.�`�6r7��n����'½h���^!��ԗ�Ei��X���Ž~rܽ�   �   ĸ����V�� X(���7�6�E�2XP��W���X�xU�K�Ō<�c()�N��Ɩ��Sƽ���Wj��q/�8���\�����k��(*���a�����<����9��{�h�6�A�W�<�y�u���Y[��O���C����h��	Ȧ����(9����|�U!X��s3�bN�`�"ʷ� ����~�6al��=p�N����������x�̽�   �   ���*��L�$��=�4!U�Yak��~���D������3僾&�v��_�tXD���&�,		��	۽�m��vv��H�T�`�4��L+�	n6�b@T�z=���j����ý��S����$��=��U�U^k��~�����6������)ヾM�v���_�YUD���&��	��۽|j���s���T���4��I+�Xk6�1>T��<��j����ý�   �   ?;����%�6���W�8�y�>���c]����������k��Wʦ����;����|�:$X�v3�ZP�Pc��̷�C����~��dl�Ap�����Ƿ��뺯���̽���Z��h���V(���7�ВE�YUP�|W���X��U��{K�z�<�_%)�������Oƽƥ���Qj�0m/�n���V会���i�2'*�!�a����������   �   ��Tt%�H\M�jx��ᑾ�ʦ�:-��KcǾ��ϾҾL?;�¾�i�����͆���`�7t7�$p����`)½`���*#���՗��j���Y��!ŽDsܽ�j��K��V��v�� "�[L(�-,���,��9*���#��������o���^ѽת�`H���E���<���~����a�����*���Ҥ	��bK��b����Ľ�   �   ���c�6� $g�m���������¾��پL�����c��rG���L���Ծ�����9������e'^�iv3���>Z�nνͫ����������u̽E�ݽ����nh�������hE�����Xo���T��B�㽼�ɽ,7������C�Z�7�4�ҼԄt�|���+����`OŻ��m����E�>�Ő��ν�   �   ����DI�j݀�S���D}���d޾#���>��D��+��������
��6۾֧�����.���C�Q��O*���?j�޽�Hؽ��ܽ��� ���
y�Ƭ	����k������'
����۲�� ]�F�ս.t��V��d���}.e���.�����\���h��� F�9к�;�<���; k�:@���hƼ��9�R���a�ڽ�   �   �#�7�Z�D;��s���>Ծo���m�e������h"�#z��N���
��d���"Ծ�Ǳ��䑾įl��k@�����
�E��0V������@W���B[���>�����E�>���`���RȽ���A��4�v���B���,O��7G����5�;�8F<���<���<La<��;�1������|9� p��s���   �   ��,�uLi��N���V�����8��p����$��Z-��R0��9-�j$�������P��$^������Dـ��Q�SA.���D�	��2���P��Z�p|��u����֭�l�����z��Hн��������,,r�T2;�h���K��D!� ��8��<|<L{�<6��<T�<f�<�](<0l'�Z۫�2�;�3��A���   �   �A3���r�=松��ž+���3��f��,��6�C9�Z6���,������Ζ�O]˾��������F�\�p�7�@��`$��=���`��K����l��&��j����O�=罡�ǽ�%���_��kR���fȼ��N����0��;t�u<"��<N��<�D�<���<��<�,H<�㩺hG��>��f�������   �   r�5�Q(v��0����Ⱦx��q�b� ���/��9��W<��9��/��C!��7����,�ξ�Ω��ቾF�`��:�I�!�(��C�����+�����_��ڝ!���1n�eV�;&�׭�9�Ľ�^��(Ă���G����*����t"� �: <�X�<�(�<���<��<pk�<�<�:R<��n�li��k�?��諒q���   �   �@3���r��坾�ž*��a3��e�]�,�#6�LB9��6���,�;��9���m\˾���ꐇ�I�\���7�����#�I=�_��������(�����M%�?j���wN�*<�Նǽ%��q_���R�z�fȼx�N���� ��;L�u<n��<���<E�<|��<x�<�.H<�ͩ��E��t�>�f��ј���   �   ��,�{Ji��M��!U�������*��<�$�xY-�cQ0�i8-��h$�d�����S��u\��4��� ؀��Q��?.�����	�X1���������
{��t�������A����/y�OGн{��������*r�1;�y��,J��$!� ��8��<x|<|�<��<^�<��<�a(<�W'��׫���;�i1������   �   �#�x�Z��9��B��<Ծ�k��8l�{������f"�x�M� �
��a��  Ծ�ű��⑾��l��h@�s���
�QA���R��
���cU���RY�
��c�N����jD�����B��#QȽ�	���@����v���B����M���4G�P��9�;�:F<о�<Ç<(a<0��;�#�����My9��m��K���   �   ��_AI�Rۀ�����z���`޾�������ߨ����$�f��k��P2۾������厁�x�Q��L*��pe�H�޽}Dؽq�ܽf�轒����v�|�	�}��R��̹�.&
�<��V���[齢�ս�r��U������\-e���.�V������0��� ��9P��;d�<���;@��:����bƼ��9�������ڽ�   �   �����6��g�����[�����¾
�پg�뾼���]��BB��H�n�Ծ����G6������h"^�Er3�:�HT�νڦ��Л��H�q̽C�ݽ����f�F�����C�g�z��<n�.�����.���ɽ�6��A�����Z�|���ҼD�t�v��+�����AŻ(�m�R�伿�>� ��ν�   �   #���p%��WM��x�gޑ��Ʀ��(��h^Ǿ`�Ͼ�Ҿ:;����e���
���Ɇ���`�$o7��k�^��4#½ڜ�����З��e��yT��Ž nܽ�e�����
�V��"��J(��,�g�,��8*���#�s��*���n��^ѽ�֪�H��^�E�Z���:���|����a����v���n�	�.^K��_����Ľ�   �   �5��7�Ɲ6�9�W�ǁy�����*Y��ﶤ�����f��sŦ�&���6��:�|�xX�Lp3�wK�[��ŷ�0����~��Zl�R7p�׎��貖�������̽��� ��4���T(���7�D�E�TP�mW���X�PU�{K��<�%)�d�������Nƽv����Pj�tl/����T�<��rg��#*���a����������   �   �{���V�$��=�eU��Zk��~�s������M��������v���_�qQD�{�&��	�� ۽�e���o��ޟT�#�4�BC+��d6�W7T��8���e����ýs{�.����$�=�U��\k��~�.������^����⃾��v���_�)UD�Ϣ&��	��۽2j���s��!�T���4�H+�;i6�-;T��:��Dg���ý�   �   r��������S(���7�g�E��QP��W�t�X��
U��wK���<��!)�6�� ����Iƽ���_Ij��e/����NJ伨�⼤c�� *��a�����9����5������6���W�׃y�ޞ���Z��븤�����sh���Ǧ����9��h�|�2!X��s3�@N��_��ɷ������~��_l�<p�����Ҵ������+�̽�   �   �f��"���~����"�]I(��,�+�,�M6*��#����B��ci���Xѽ�Ѫ��C����E����b/��.s����a�����𪶼��	��[K�
_��Z�ĽJ��Eq%��XM�fx��ߑ�fȦ��*���`Ǿ��ϾS
Ҿ�<;T���~g������ˆ��`�r7�gn�����&½����� ��<ӗ�-h���V���Ž�oܽ�   �   5	�}f�x�����C�z�,���l�@��������_�ɽ2�����Z�����Ҽ�lt��P�P�+� Z�)Ż��m�����>�r���bν&��o�6�� g�r�������5�¾��پ���"��O`���D���J���Ծڧ��R8������m%^��t3�]��W�<ν����Z�������2s̽F�ݽ\���   �   =�	������ڹ��%
���������X�؄ս�o���Q��<����&e�9�.�r���`x������ ��9���;<�<h��;��:z��^Ƽ"�9����~�ڽB���AI��ۀ�y���){��Db޾�������������c��������4۾�������X�����Q��N*���hh��޽�Fؽ��ܽ{�轃����w��   �   �������% �^D�'���4�ཤOȽ���n>��эv���B�7��dD��8#G����XV�;hGF<^ā<�Ǉ<�a< ��;��������w9�Pm���罩#���Z��9������<Ծ m���l�M������g"�,y� N�*�
��c���!ԾǱ�䑾ͮl��j@�����
��C���T�����PV���"Z��   �   $u�����x�����x��Fн����n����'r�6.;�l��D���� � f�8��<(|<���<���<��< �<�g(<0@'�
ի�v�;��0�������,��Ji��M��hU��6��m�����ʚ$�!Z-� R0�59-�oi$�4�������澷]��H���ـ���Q��@.�����	�.2�e��������{��   �   ���%��j�2���N�6<罱�ǽ�$�� _��kR� ��bȼ$�N� �����;0v<H��<8��<xG�<ܱ�<��<P3H<����C���>�Te������@3�r�r�n坾��ž-��r3�f���,�r6��B9�6�o�,����������N]˾��������c�\���7�E��T$��=���� �� ������   �   4\��k{�1�o��O]���E��'+�l6�43�����Y��V�1���ϼ��!� �G;��]<�Y�<���<���<�=��<���<���<��<��Ȼ:yԼ�RQ�(V�������I'��Z�̙��-,��������پ�o�����l�����̥��ھ�Tþ'&��7�����w� �T�v <���.�͝+�,�1�1�>��\O��"a�i�p��v{��   �   ՠ{�G�w���l�o�Z�D��(*������p���~Ѕ�v�7��Dݼ��>� �:@B<̈�<�8�<�I�<Xh�<,�<x��<�a�<�<�޻/ؼ�Q�ħ�:��%�ŉW�L݆��墾��uq־�������K�����׻�#׾����N���(��kos� Q�=�8�#�+�q�(���.��G;���K�Yw]���l��w��   �   ��p�0n�|Rd�d<T�Ud?�H�'�rA��&���N�����J�����-��e�����;�~{<�б<M�<�}�<P��<&e�<2Ѓ<�з;Pt�(6伕IT��i��Ȁ�N3!�P�䁾�\��r����̾��޾���\��!꾅c޾��̾,���=��T��kEg��xF�#v/���"�F �J�%�?�1���A���R���a�T|l��   �   d�`�]T_��W�.`J���8�)$�$������Ľ����l��(�B׼�dW��*��P �;�Lk<:��<���<�<:�<��8<`��:�O��Q���+Z��d���8轑��#
F�|�t��h������`:��]qξ��ؾK�۾�׾��̾�6��h����3����y�:T���5��� �����r�����B#�SK2��UB�]�P�#t[��   �   �L�4dM�E�H��+?���1�L�!���������@ֽ����T^��\`���#�2ټ �m�Ս��Qw;�<�jO<ȖT<�L'<�[�;�	��Z:������Mf�vy��$����m�9�d�b��N��F\������ڹ�:`¾��ľD���s���ד��Eh���⁾Ȼ]��;�>� �g���8�"���Ҕ����ܖ-�"�;�<bF��   �   ?)7��:�ߣ9�ܲ4�"r,���!��(R�|���ӽ*���v���p�Ci6�� �T1��d((�p|R� ��:��; �88���ql��?ۼ�-�0�{�����<d����/.��jP���r��퉾C��e;������M���া>����p��Ā��&�^��=�?D �����ټݽ�=ڽ���D���kH�)|�$�l/��   �   �i"�E)��,���,���*�*&�hX������Ѫ �Wz潡ɽ(�����EX��� ���|n��8]�:���Q�h����׼�7���V���������n�㽨�
�7�$���?�-�Z�s�s����q���YҐ�kߐ�珌��4��
-q��U�K�8��>�� ���ݽ���������	���Ѹ�y�ʽH�������w�y���   �   )���V!#�J�)���-��0�Q�/��-��_'�)�����t���\�Ľpw������GH�y���"���-Ἲ��R�U�'�j=U��������i�ɽ�3｜&��+�i!3�*AF�fyW���e�Lo�b�r��.p���f�jsW��C���+���d��wg̽ƪ�wp���;����>���8^�� F��1�н`�����   �   ����z������+�G7�)�@��QG��J��I���C�]�9���*������,�߽xY������Wt��N�|�;�?<�_�M���n��č���*ƽ��佑���z����h�+�77���@��OG���J�g�I��C���9��*�7����^�߽'V�� ����Rt�}�N��;��<��M�5�n���ԟ��)ƽV���   �    3ｴ&�h,�f"3��BF�Z{W��e�o�S�r��1p���f�EvW�bC���+����g���j̽�Ȫ��r��2>��<􅽔����`���H����н���#���)�����!#��)��-��0���/�-��]'��������q��罠�Ľt������BH�������%�4�O���'��9U�k���C���g�ɽ�   �   ����
��$���?��Z���s�n��������Ӑ�ᐾ����B6���/q�o�U�e�8�N@�J"�b�ݽ���]�����Ը�	�ʽ��⽑���Gy�����j"�$)���,���,�N�*��&�fW�������� ��v�ɽ�	�����s?X��� �伐f���)]��:���Q�^�׼"5�N�V�ر��p����   �   �dཬ��$0.�(lP��s���D���<��Q�������⦾�����q��󁀾-�^���=��E �d��R���ݽ�?ڽ�������I��}�n$�mm/�{*7�#�:���9�M�4�4r,�V�!�t�@Q�6��|�ӽm��t��czp�Gd6�� �4)���(��HR����:@&; �8��\il��;ۼ��-�w�{������   �   2������9��b��O���]��c��ܹ��a¾1�ľǡ��ڈ�����Ui��~まF�]�S�;�Q� �h���9�������6��4�-��;��cF�%�L�AeM��H�,?�$�1�=�!���������>ֽ����S\��6`���#��ټ(�m�(���@~w;��<�sO<ԞT<0T'< i�;����8��;���Mf��y���   �   ):�~��dF��t��i�������;���rξa�ؾ��۾G�׾��̾�7��=����4����y�	;T���5�S� ����~s�l���C#�^L2��VB���P�Iu[�t�`�OU_�êW��`J��8�&)$��#�B�ｷ�Ľc��l�*�(�V<׼�YW�@��� 2�;�Tk<���<���<��<j�<��8< �:�O��Q���,Z�Fe���   �   ��/4!�C�P��䁾m]��d����̾
�޾���]��"�Nd޾��̾�����������Eg�6yF��v/�a�"�� ���%���1���A���R���a�(}l�g�p��0n�Sd��<T��d?�\�'�[A�U&�q��������J����6*���W����;\�{<�ұ<O�<~�<ƴ�<0f�<�Ѓ<�ѷ;�t�47伝JT��j���   �   4;�ױ%���W��݆�y梾���r־U�龊��RL��n���*��\׾����N���(��kos�Q�A�8�3�+���(�/�.�-H;�!�K��w]���l�x�w�6�{���w��l���Z�+D��(*����7�����Ѕ���7��BݼL�>��-�:�BB<���<�9�<�J�<�h�<^�<���<va�<��<P�޻�0ؼX�Q��ħ��   �   ����~J'��Z����,��B����پ�o�����l���������ھ=Tþ�%��ꙑ��w���T� <���.���+���1��>��\O��"a�S�p��v{�\��k{��o��O]���E��'+�N6��2罟���Y��.�1�`�ϼ�!��G;��]<PY�<��<��<��= ��<��<P��<��<�Ȼ�{Լ%TQ��V���   �   :��%�W�E݆��墾���6q־W��}��@K��`���(��n׾#��N��<(��Tns�.Q�g�8�g�+�Ȧ(�b�.�MG;�2�K��v]���l�`�w��{���w�	�l���Z�XD��'*�8��?��D���pυ���7��Aݼ,>�`;�: DB<r��<:�<�J�<8i�<��<���< b�<��<��޻�.ؼ�Q�ħ��   �   ���2!��~P��ま \�������̾'�޾ �꾶[ �cb޾��̾���A��p���Cg�hwF��t/���"�@ �J�%�?�1���A���R���a�{l�N�p��.n�Qd�;T��b?��'�6@�t$����T�����J����0(��PQ�����;\�{<�ӱ<�O�<6��<���<Pg�<X҃<�ٷ;�o��3�7HT�i���   �   -7轕���F��t�#h������I9�� pξ��ؾ��۾��׾A�̾t5������2��X�y�)8T�D�5�� ����dq�B���A#��I2�TB���P�er[���`�xR_��W�A^J�ֵ8�B'$�D"���｢�Ľ���l�?�(�x9׼�UW�@���87�;�Vk<���<���<��<�<��8<�4�:��N��L��G)Z�c���   �   ��⽖����9��b��M��[������ع��^¾ܷľ}�������*����f��2ၾG�]���;�K� ����@7��	�1�7��@��	�-�'�;�`F���L��aM��H�')?���1���!��������w<ֽЇ���Z���`�	�#�
ټd�m������w;��<DvO<�T<�W'<0r�;򮻾3��=���If�6w���   �   a�.���,.�FhP�2�r�쉾yA���9��θ��i��ߦ�_����n�� ��*�^�[�=��A ���H��d�ݽ\:ڽ)�㽾����F�z��$��i/��&7�z�:�)�9��4�]o,��!�b��O�}��\�ӽ����r���xp��b6�� �\'���(� >R���: 4; �8�賻8bl�7ۼo�-���{������   �   ��㽌�
��$���?�Q�Z�U�s�`�������tА�yݐ������2��z)q���U�R�8��;�f���ݽި��w~��9��θ�͙ʽT�⽉����u����f"�n)�(�,���,�r�*�&�SU����,��� �u��ɽ���M���Z>X��� ���0e���&]�`:�ĭQ��푼v׼�2���V�����j����   �   S/�F$�])��3�2>F�7vW�=~e��o���r�+p�2�f��oW�cC��+�8���^���b̽ª��l��b8��������Z��-B����н���~��>&�'��?#�
�)�S�-�/0���/�g-�o\'�������Kq�����Ľ�s������BH�-�����P$�&��M���'�}7U�ʘ�����x�ɽ�   �   B��nx�����+�?7���@��LG�Q�J��I���C�E�9���*�����1�߽}Q��򬕽�Jt���N���;�r<�r�M�&yn�ξ������`$ƽH��>���w�~����+��7���@�2NG�G�J�?�I�+�C��9���*���������߽�U��Ȱ���Qt�ͮN�S�;�<��M��~n�����X����&ƽ����   �   �'�*���#�X�)�-�-��0���/��
-��Z'�ٜ�����n�~�罏�Ľ�o��퍀�Q;H��������$��H� �'��2U�z���㢦���ɽ�-��#�?)��3�?F��wW��e�o�c�r�.p�W�f��rW�pC�^�+�����c��*g̽�Ū�*p���;���񅽵����]��.E����н�������   �   ih"��)��,��,���*��&��T����ƍ�c� �~q�ɽ�������7X�i� �伲Z���]���9���Q�N呼.׼�.��V�ʭ���������M�
��$���?�d�Z���s�p��������ѐ�ߐ������4���,q�ͯU� �8�Z>�� �n�ݽb�������V	��.Ѹ��ʽ�������2w�����   �   =(7�Җ:�C�9��4��o,��!���N�����ӽ
���o���rp�]6�e� �<��(���Q�@��:�o; < 8@ͳ��Tl��0ۼS�-�1�{�����L`���@-.��hP�`�r��쉾�B���:��V������া����p�������^��=�$D �����｜�ݽp=ڽ7������H��{�q$�Mk/��   �   )�L�9cM��H�*?��1�@�!��������8;ֽ)����X���`���#�,ټP�m�蕍���w;,�<,�O<�T<tc'<興;�ۮ�n.�����wGf�\v���⽓���9�.�b�`N���[�����;ڹ�`¾q�ľ%���^���Ǔ��9h���⁾��]���;�)� �U���8������������-���;��aF��   �   ٗ`��S_�#�W�_J�s�8��'$�\"�\���Ľ���l�T�(�@3׼�HW��\���N�;�ak<���<�Ư<��<��<L�8<�z�:�N��H��w'Z�Jb���6轌��-	F���t��h��?���!:��-qξ׭ؾ1�۾�׾��̾�6��`����3����y�:T���5��� �����r�y���B#�+K2�jUB��P��s[��   �   H�p��/n��Qd��;T��c?�W�'�a@�p$꽞������j�J�ľ�2$���@��x �;�{<\ױ<jS�<���<и�<�j�<�Ճ<��;�h�T0伤FT�\h��^2!��~P��ま[\��@��Z�̾��޾��꾲\��!�~c޾��̾(���8��O��cEg��xF�v/���"�8 �7�%�-�1���A���R���a�|l��   �   ��{��w���l��Z��D�/(*�a��\��;���>υ���7��?ݼ8{>��]�:hHB<���<2<�<M�<Fk�<��<��<vd�<d�<��޻F,ؼ��Q�Qç�Z9�ư%�z�W�,݆��墾��bq־�������K������ӻ�!׾����N���(��ios�Q�9�8��+�i�(���.��G;���K�Hw]�i�l���w��   �   ��ž�2¾X����n��b]��������U���*�F��!C������)�l#�� ��9$�X<��<��<�=�=�=���<�Z�<�7k<�%;%M����N�Y������޽�E�<{5��Z��(~��玾d���a��Y��`d��Sś��`��ς���i���P�9�=��K3���2�:�<�o�P���l��l��񁙾򨪾0Ӹ�c4¾�   �   �]¾~.��mµ�����`���~��zS�LC)���x��8Y��U�������N�xwF<`�<���<3�=Vd=�U=��<jӳ<�U<��:XXa��j��!]�� ����޽���k4�3QX��({����E0��$�����Ǡ��<������j�����e�U2M�m�:��-0���/��r9�`M���h��%���򖾢֧��˵�����   �   ^J���~��Э�|������0v��LM��w%�[] �@��P���%��ҥ�����l<���<���<���<���<ک�<^B�<��<��<�6��Տ�^-���g�����޽���q30�!R�>�r������ے��噾���v?���瑾o��ҕt�XZ�j�B�*�0��'�!�&���/�ܤB��-]��}�m���ͧ���������   �   �L��%�����Ύ��$����h��DD��4 �����cw���|��%6� ^ϼ����A;4[K<N�<B�<tj�<(̵< 3�<0�:<И;�A���Ƽ1�)�*�{�Η�������<�*�+I���e��^7��l!�����̡��������x���`��kH�2�2��"�$��1\�'!��R2���J��ih�(��뒾i���姾�   �   &ڙ�픘�z���ʮ���_w�B�Y�:%:����t���B:Ľ�v���TQ�������'�� l};��+<�ci<��x<t3[<d}<�`�:�������c�H�O�
���W��r��F���%��?�>�V�/}k��z�B߁�v���F~���p���]���G���1����v��ˌ������s��3��%N��j��؂��K��:I���   �   �����w��Ri����u�Y�a�@J� �0��k�/U��}�ν�ӣ���y�P�4����I���n����Q�p�G; �}; ��:��\��97�P���5�:�E�*%��6��$�˽���0��]I"�t6�54H��CW�d�a�Zg�]�e��I^�*�P�Zb?�+����x2�B��i%�E����A���	��k0��|I�[�a��tv����   �   �f���h�o�d���[��N��H=��*��G���.=��Y���[��Ԏq�i�6�����y��<mu��d3�D�'�S�Jr��$Q����i�T�>a��P觽�/ȽW��K�A��f�"��:0���;���D��J�B�J���F�J>��0��D ��U�6|��էڽ�zý����7���7^����ؽ�X��|d�[;'��<��oO���]��   �   �BB�X�G�.gH�NE�S#>�,�4�I�(�������m���R޽𰾽�l��TɁ��N�׹"����:0��;ݼ����U��nOA��2u�m3������J׽70��qj�)��Q��#(��/���3�J'6���5��1��s*�3���
�H\�H��Y�Ľj��t:�����q��7ђ������7ýh��e��E��o *�cD8��   �   ��"��9+���0��3�ܝ3��B1�Ӭ,���%���%���R2�`ν"���8*��Y&v�j�R���>���<�W�L�`n��Y���)���^ν�r��r�|��a�"�!;+���0���3��3�qB1�9�,���%�����-�2/�]νA����'��H!v���R��>��<�B�L��Zn��V���&��h[ν�n�q�����   �   (i�"��`P�`#(��/�z�3�C(6�
�5���1��u*������]�r��H�Ľ�l�� =�������
���Ӓ������:ý��e��g���"*��F8��DB�,�G��hH�hE��#>�c�4��(���.���k���P޽X���bj���Ɓ�[�N�\�"�����'�`3ݼ������1JA��,u�j0��ݟ��4׽M-���   �   ���fJ������"�*;0���;�0�D��J��J���F�A>�̶0��F ��W�3����ڽL}ý6���ƶ���`���ؽ\��ff�z='�i�<��qO��]�W�f���h�;e���[��N�+I=� �*��G�����;��W���Y����q�N�6����Br��T^u�LV3���'���R�2j��pH�U����T��^���姽�-Ƚ�   �   �˽M��B���I"�D6�^5H�EW�(�a�Kg�c�e��K^��P�"d?�^�+�'���3�����'㽈G⽦�ｼ�����m0�I���a��vv�(Ă�0����x��Jj��Y�u���a��@J�]�0��k��T��t�ν:ң���y��4���B��XV�� �P�`�G;0�}; a�:�\��+7� � ���E�#���4���   �   0W���潗����%��?���V��~k���z�4���w��cH~�t�p�%�]��G��1�������ԍ���:���t���3�R'N��j��ق�M��fJ��Lۙ�����m��������`w��Y��%:����F����9Ľv��PRQ�������8��0�};��+<�li<��x<�<[<�<`��:���p���a��O�:���   �   ח��|��y����*�-I� �e���-8��D"��㥐�����P���мx���`��lH��2��"����]�!��S2�)�J�kh����쒾j���槾�M���%��ޤ��}������i�h�iED��4 �����
w��6|���6��Zϼ����A;�aK<@Q�<b�<�m�<nϵ<h6�<�:<��;�:���Ƽ�)���{��   �   \��n�޽~��*40��!R�Q�r�����6ܒ��晾4��
@��?葾�����t��XZ���B���0�+'���&�y�/���B��.]�}����z������>���K��`���Э���������v�=MM�$x%�`] �������%%��Х�Ȃ���p<���<���<���<���<ޫ�<0D�<��<�<`�6��ԏ�-���g��   �   I��g�޽,��4��QX��){�S���0���ڄ��Ƞ��<������������e�k2M���:��-0���/�<s9��M�Y�h�&�����֧�&̵� ��&^¾�.���µ�����`��L�~� {S�VC)���M���X����������N�\yF<�`�<F��<z�=�d=�U=���<�ӳ<`�U< �:Ya�7k�h"]��   �   2����޽=F��{5�t�Z�
)~��玾�d���a��Z��Rd��7ś��`���΂���i�j�P���=�8K3�J�2��<�P�P���l��l���𨪾.Ӹ�]4¾��ž�2¾F����n��M]��������U�y�*�'���B�������(�^#�� ~�9��X<̆�<���<F=��=�=ֶ�<�Y�<�5k<�%;\(M����u�Y��   �   � ��l�޽���C4��PX��({����0���%���bǠ�<��U���򟀾��e�1M���:�,-0��/�`r9��M�M�h�p%��>�@֧�Y˵�+��N]¾ .������>��Y`��8�~�zS��B)��l��NX��� �"�����N��zF<�a�<Ԡ�<��=�d=V=��<^Գ<ԝU<���:TVa�Uj�7!]��   �   �����޽P���20�7 R�J�r�p����ڒ�8噾����>���摾���\�t��VZ�!�B��0��'��&���/�ףB��,]��}������@������|I���}��<ϭ����ǭ���v��KM��v%�E\ �V������,%��ͥ�z���s<Ύ�<���<Z��<r��<���<$E�<���<�<�6�ҏ�b+���g��   �   ƕ����������*��I�T�e�^�s6��p ����� ��������x���`��iH���2�z"�����Z��!�_Q2�c�J��gh�:����꒾�g���䧾pK���#��Ӣ����������h�
CD��2 ������t��az���6��Vϼ����/A;$eK<�R�<��<�n�<�е<�7�< �:<0�;�5�>�Ƽ��)�j�{��   �   �T��Z�潞��A�%�?�1�V� {k���z�
ށ��t��D~�9�p�5�]�x�G���1�������2���y���q�@�3��#N��j��ׂ��J���G���ؙ�m��� ���X����\w���Y��":���������6Ľ�s��OQ�<��V ���	���};�+<|oi<\�x<�?[<�<���:��B���_�C�O�V���   �   i�˽�����'G"�!6��1H��@W���a��g���e�G^���P��_?�k�+����y0�����!㽶A⽗��p�����i0�szI���a��qv�\���\���v���g����u�B�a�,=J�J�0�Ui��P��R�ν�ϣ���y�l�4���?���L��@�P���G;��};�y�:��\��'7�z민��
�?�E��!���2���   �   ѐ轩H����ץ"� 80���;��D�J�]�J���F�w�=�+�0�YB ��S��w��̣ڽ�vý,��������Z��4�ؽ�T��8b��8'�W�<��lO�d�]��f�?�h���d�(�[�� N�wE=��*�1E����h8�kU���W���q�G�6�����o���Zu�,S3���'���R�vh��NF�	����T��]��W䧽�+Ƚ�   �   �g�y��LN�� (��/��3�\$6�˔5�!�1��p*�l��,��Y����}Ľ.f���6���������͒������3ý���������v*�1A8�D?B��G��cH���D��>�݈4��(����?��~h��*N޽����i���Ł��N�@�"����J&��1ݼ�������0IA��+u��/�������׽J+���   �   ��"�-8+���0���3��3�y?1�H�,���%��
�����4*��Xν��#���v�ƠR���>���<���L��Sn�,S��"���Vν�i�Bn����|"�Z6+�q�0�x�3�i�3�@?1���,���%���S���-�n\ν^����&��L v�ԦR�]�>�j�<���L��Yn��V�� &���Zν�m�bp�����   �   �AB��G��eH�N E�� >�p�4�3�(�I�����sf���K޽Ω��$f����5zN���"�k���⼆'ݼ�����6CA�,%u�(,��&���	׽�'��0f���%M� (��/��3��$6�ӕ5���1��r*�J��"
��[����ĀĽ�i��:������&���В�\���G7ý���������*��C8��   �   4�f���h��d��[��N�[F=�q�*�,E� ��
7὚S���U��F�q���6�F���f��pHu�DA3���'�L�R��^��<Ἄ���T��Z��T᧽�(Ƚ.�轎G����c�"��70�g�;���D�VJ���J���F�� >�Q�0�|D ��U��{��t�ڽhzýp��������]����ؽQX��Ed�;'�Û<�oO���]��   �   ����Ww���h��t�u���a�G>J���0��i�nP����ν�Σ���y���4���� 8��0/��@�O���G;@~;���:Pc\��7�p⯼�
�g}E����=0��f�˽>�����F"�P6�\2H��AW�#�a�\g���e�*I^���P�	b?���+����R2���0%��D����"���	��k0��|I��a�+tv����   �   �ٙ��������L���s^w��Y��#:����ϣ��v6Ľ%s���LQ��������p�`�};��+<X{i<4�x<�K[<�<�=�:l���{��%[�}�O����3S��,��D��2�%�W?���V�|k�&�z��ށ��u��F~�Z�p�L�]�}�G���1����]����������ns��3�r%N���j��؂��K��I���   �   �L���$��ǣ��v��������h��CD�u3 ������t���y���6�XSϼ��QA;�mK<�V�<��<<s�<$յ<�<�<\�:<��;d*�R�Ƽ��)���{�������ཎ����*��I���e�<�
7��+!��ڤ������z���\�x���`��kH��2��"���"\�!��R2���J��ih���뒾�h���姾�   �   FJ���~���ϭ�D��U����v�/LM�.w%��\ �~������w%��˥�p���y<���<���<v��<���<���<�H�<^��<��< q6��͏�0)���g������޽���20�N R���r�����_ے��噾w��a?���瑾f��Õt��WZ�[�B�"�0��'��&���/�ҤB��-]��}�d���ħ�����r����   �   �]¾m.��Zµ�����`����~��zS��B)�D����TX��� �$�����N��}F< c�<~��<��=�e=W=��<�ֳ<��U<@$�:�Pa��h��]�������޽=��4��PX��({����,0��u����Ǡ��<������f�����e�N2M�k�:��-0���/��r9�YM���h��%���򖾜֧��˵�����   �   P��Y���
�z��������%Z��0�{���@�p��m"���p��:��D��L<Rc�<�C�<�>=ڎ
=�O=,q�<���<`�}<�Ϻ;��ǻ�����1��[�'ɕ�P�����sN���#���6�E�E���N�K�Q�l�N�S�F�P];�//�j�$��Z��w!��J-��ND��g�4w���量5-ľ�⾒�����
����   �   x@�ʾ��l�����Nݾ�*��#$��1�x�Yq>�{I����e�o�|�������<��<���<�� =�=�2�<0n�<�+�<`B^<оn;8��'���?�b� ���q1ý������#��S5�{C��PL�OO���K��C��H8�,�h�!���0��4A*�.�@�
c����#��|���/�޾����o����   �   �/�k�����u���dӾ����ɕ�lKo�q8�pQ�ƨ��a�m������"��\�;}�<6�<���<��<���<x&�<�3�<`��;0@,�p�p����4"3��,x�����>Yɽys�	��� ��1��=�m�D���F���B�;�:��`/���#���Jo��W��g!�6�6�ޑW�LG��%���Q��M�Ӿ�=������   �   �8 �#u���"𾂼ܾ�&ľȐ��*���%a�"s.�+���[���l��
�8N�P�;\�U</�<jU�<Z}�<��<�m<"�;�_�3[���Ӽj1"��^��̏��屽;ս������]����*�
�4���9��:�"e5���,��!�#�ױ�@���Q	��}�k'���E��/m��Q��j����¾]۾v��0����   �   k��J��pI׾��ƾ�@���8���R��6P�UY#�����ꩱ�M?o��J���� �B���;��L<<Qp<�]< �<@�6;�Ȼj�����8-�=f��K������F�˽��л�������8�$���*���,���*���$�v��R�f4��Z����9�T��|��t.� �Q�[g|�j�������¾��Ծ[K��   �   ])ƾiľ�λ�K2��
���/�����g��>�;��V콢�����x��[#��"���-�������:;@7�;�.�:������O�����wV��%M�������2���ؽ�l�'��F������)��C ���!����������ҟ�c���r�H�ҽc_ɽf�ʽ�`ڽZV��6$�c3���W�{:��ɹ��^����-������   �   
Φ������V(����p�#�O�E�.�i�����ܩ��K���o@�j�2+��|�U��7�|���_�<��Na�{a:�D�x�z�������޽����K	�$����H��Y� ��!�B0�������3�����뽷�ӽ�f�������#��jv������M�ȽԴ� ����1��(T�p�v�����#���`���   �   �g�� 텾�~�\�j��+T���;���"�&B
�M�/��
ە��)i��2��5��Sڼ��ļzFҼ�Q�_*���b�Zt��|����eὠ���a�w�#��{.��5��7�-�6�{2���+���"�͏�g�� �F��!wɽ� ��Z���v�v�N5t�����J���h`�����]S�b�(���E�wa��x��_���   �   �5\���_�$�]�ÝV�a4K���<��d,�j��{8	�J$�j�̽�m���	���l���E��(.���'���4��HU�p愽����nҽ`� �����n/�a9C��}R�9\���_���]���V� 6K��<�te,����O8	�\#��̽l�����#l���E��$.�1�'��4��CU�Pㄽ����jҽ�� �؜��k/�G6C��zR��   �   #y.�s5��7���6��y2�J�+�y�"�������� �
 �yɽ�"��-�}�����v��9t�����/����c����佮U��(���E��a�
x��a��J����h��b
~�g�j�-T�Ú;�+�"�BB
��~�J���ٕ�'i��2�n2��Lڼ��ļ>Ҽ�L�}Y*���b��p��U����`� ��_���#��   �   �I	�g�����.���� ��!�[0�^�����4���������ӽ+i�������%���x������E�ȽT����R�1��+T���v�j���	���b���Ϧ�|������]����)����p�g�O��.�ƪ����d���v���m@����%��l�U�d*����`	_�����[�M[:�T�x���������}޽߮���   �   +�ؽBj�2���������)�ZD �6�!�������������Fe��u�n�ҽ�aɽ��ʽxcڽ:Y���%�j3���W��;��f���(���}/�����T+ƾLľ�л��3��H���'�����g��>�Â��콀�����x�Z#���� w-�@��� ;;�N�;���:8�����O�����Q��M����陡����   �   ������˽r齆����������$�P�*���,���*���$�)w��S�h5��\����;�q��^}�Bv.���Q��i|��������7�¾T�Ծ9M�F����K׾�ƾ�A���9��cS��7P��Y#��������>o��I����B� �;�L<dZp<��]<��<�6;��ǻF�6��-��f��I���   �   fˏ��䱽�:ս������ȡ�w�*�ι4�j�9��:�f5���,�ܗ!��#���� ���R	�t~�)l'��E��1m��R��.k��.�¾�۾���İ��q9 ��v��$𾸽ܾ�'ľ�������s&a��s.�s���[��ҽl��	��N���;��U<�1�<�X�<���<��<�&m<7�;�1��&[�|�Ӽs."�H�^��   �   w+x�:���8Yɽ�s�T��y� ��1���=��D�m�F�D�B�ٚ:�"a/��#�����o�oX�2h!���6�˒W��G������R��>�Ӿ�>�@����40����q �R�eӾe��ʕ�Lo��8��Q�꨻�E�m�D��p�"�(b�;�~�<��<���<
�<��<:)�<7�<���;$,�|�p�J��� 3��   �   b�+����1ý>��#�#�T5��C�)QL��O��K�\�C��H8�E,���!�@��_��tA*���@��c�,��g#��������޾H���io�R���@���<m�_���Nݾ�*��P$��o�x�wq>��I����A�o��������<<�<v��<�� =v�=�3�<Bo�<�,�<�D^<��n;(��>&��l?��   �   �[��ɕ��P��7�N���#�&�6�p�E���N�R�Q�^�N�5�F�$];��/�2�$��Z��w!�dJ-��ND�ug�4w���量>-ľ�⾘�����
���L��R���
�b��������
Z���{�x�@�N��:"����p��:����<&c�<PC�<�>=��
=dO=�p�<<��}<�˺;��ǻ�����2��   �   b�~����0ý7�ｊ�f#�;S5�C�BPL��O�0�K�t�C�H8�x,���!��������@*���@�zc�����"�������޾1����n����!@�s���l�N���Mݾ*���#��_�x��p>��H�$�����o���������<�<���<� =��=�3�<�o�<4-�<�E^<`�n;<�� %���>��   �   p)x������Wɽ�q�.��"� �1��=�e�D���F���B�$�:��_/�y�#� ��Vn� W��f!�B�6�ՐW��F��w���P��f�Ӿ�<� ����/����V��L���cӾ����ȕ��Io�98�jP�����m�2{��t�"��j�;6��< �<���<��<ʫ�<*�<8�<���;,��p����I3��   �   �ɏ�㱽S8սU���,����f�*���4��9�i:��c5�G�,���!��!���� ���P	�U|��i'�-�E�N.m��P���h����¾�۾�����7 �is��� ��ܾH%ľz������#a�rq.����hY����l���N� �;��U<p3�<�Y�<��<
��<)m<�;�;&��"[��Ӽ�,"�!�^��   �   N󭽔�˽�������Ǝ�K�$���*���,���*���$�Lt��P��2��W������6�ޢ��z��r.��Q�e|����}����¾��Ծ\I�[��8��qG׾��ƾ�>��7��LQ���3P�CW#�����榱�:o�NF�$����B��&�;��L<p]p<��]<4�<P�6;0�ǻ���(
-��f�{H���   �   X�ؽ�g����ޓ����b'��A �L�!����������ڝ�N_��co���ҽ6\ɽD�ʽ�]ڽ�R��Q"�6	3��W�9����������+������'ƾ,ľ�̻�80�����r���y�g�_�>���>������x�QV#�x��Lo-�@X��p#;;�U�;@��:������O�
���P��M����Ԙ������   �   �H	�?��+��h���� �!��-�j�t���1�������ܘӽRc��[���V ��0s��������Ƚ�𽿋�P�1��%T��v��������^���˦�_����ɻ��V&���p���O�^�.�է�Q��䥲������i@�)��!����U�&�4��P_�t��0[�Z:�j�x��������|޽u����   �   Gx.�Z5���7��6��w2���+���"�������	 �����rɽ���ꗽ����v��.t�����ȡ���\��D���P���(�J�E��a��x��]��P숾�d���ꅾ�~�e�j��'T�k�;���"�r?
��z��
��Oו�Q#i��2�l0��Iڼ��ļH<ҼL��X*�܊b�Np��ݟ��L`὿���^�/�#��   �   /5\���_���]�@�V��2K���<�wb,�����5	��ｱ�̽h��:��Jl�[�E��.�*�'��y4��<U��߄�����eҽH� �љ��h/��2C��vR��1\���_��]�ǙV��0K�n�<��a,�h���5	�[��̽�i��>���l���E��#.�<�'� 4��BU��ℽ���@jҽ�� �����k/��5C�?zR��   �   0�f��x셾�~���j��)T���;�i�"��?
�Xz�&
��֕�+ i�Y2��,�4Aڼ��ļ�2Ҽ�F��R*��b�rl������w[����[�[�#�~u.��5�_�7��6�\v2��+�N�"���)��P
 ����uɽj��헽����O�v�t4t���������`��^��4S�4�(�Y�E�/a�4x��_���   �   �ͦ�R󥾨��e����'��:�p�r�O�h�.�j����彚�������g@�Y�B��|�U��������^�"��_U��S:��x�����c���+x޽Ҩ��~F	�$��U���~�r� �m!�g-������t2�ɱ��뽀�ӽf�����"#��v�������Ƚ���ߍ���1��(T�E�v���������`���   �   +)ƾ,ľ�λ��1����������9�g���>������0�����x��T#�>��Le-�` ��@U;;8q�;`+�:0i��P�O�>���J�M�\��*���	����ؽ�d�^��ƒ����'��A ���!�O��������'��b��+r���ҽ_ɽ�ʽ�`ڽ&V��$�I3�l�W�l:������J���w-�������   �   J����6I׾M�ƾZ@��;8��.R���4P�X#����D����9o�YE�B��ЗB��7�;��L<Xhp<��]<��<�7;��ǻ�剼���-���e��E����$�˽�
�#��@�����w�$��*�q�,���*���$��u�CR�&4�^Z��^��j9�<���{��t.���Q�Hg|�_������{�¾v�ԾBK��   �   �8 �u���"�N�ܾ~&ľ|�������$a�Er.�A���Y��"�l���� N�P�;�U<7�<�]�<���<��<�4m<pU�;����[���Ӽ�("���^��Ǐ�Bᱽ�6ս>�����������*��4���9�L:��d5�j�,�Ö!��"����&���Q	�~}�k'���E��/m��Q��j����¾T۾j�� ����   �   �/�b�����V���dӾ���zɕ��Jo��8��P�������m��z��X�"��p�;��<`"�<b��<� �<Z��<.�<x<�<��; �+���p����M3��&x������Vɽ�p���� �.1�A�=���D�U�F�J�B��:�h`/�c�#���9o��W��g!�,�6�֑W�HG�� ���Q��G�Ӿ�=������   �   t@�Ǿ��l�����Nݾ�*��	$����x�q>�4I�����-�o��������<�<B��<�� =��=6�<�q�<�/�<�K^<�n;`��`!���<�'b�����0ý���E�=#�1S5�*C�~PL�O���K���C��H8�,�[�!���,��0A*�'�@�c����#��y���,�޾����o����   �   �X���T���I�9���#�&��N���������L�ξ��丽��S��^����㹜|q<�z�< R�<n��<P��<���<У<$�M<��w;��ƻX���<N缓�$��bX�3����3��3غ�xPҽ�0潓��� ��Y �&���������}��e��˫���@�<q�������r������:$�*E9�J�*�T��   �   �U�~jQ�ֳF��6��� ��T	�P;�*Ƴ������J������zTQ�
���@�1� �h<���<�A�<z.�<�S�<X��<Y�<4�!<�;Z:���7��� ���1�Xd������@��ʼ��v�ӽ����c���K��V*������~�����d������{�`��~s=�X�l�Ņ��<r����p�
��{!�2/6�g�F��bQ��   �   ��J��MG�o(=��R-��Q������׾̫�H�����A�fz�PQ���~K��N�� @Ǻ��L<,"�<J��<�0�<x��<ۏ<ț*< ��:F��������K�)���X�����]���챽b�ƽ��ٽ�x�j��������k��܃�t��S��"'齢���v��R�3��`�_������Y۾ش�	��v;-���<��/G��   �   ��:�ދ7��M.����������Ǿ���upu�M5�����(&����C��G��`�T�\�<���<p�<���<�*d<�s�; D�[G�vV��:x�O�@�xp���������"��H�ȽQ	ؽ�p�G����t��q
�~��+�ڽ�ҽx'Ͻ1�Խ�^轫���N$��	N�D�����zɾ<���G���-�nG7��   �   �=&���#�'�����kv���Tپ`'��8Z���Q_�C"&���8֜�$�<��F�� �˻@�;L%<А3<ȡ�;�ġ:|)�4D����5j;�5�r�����`-�� O��'ӽdI὚�&Q�#���h��B��'��P_�i�ս`Ƚ�a��BԷ��^���˽$�����H�5�S�f������ղ���־;����������"#��   �   �Z��L�5������&�ܾ;𽾡V��%���{G�Q��WؽBT���9�P}̼��0�P���<�: ع���ǻp�~��弌n/�_�q�6�������ڽ~��/����
�(V��W�����A
����*
������ٽ��ƽ�!������@�������G��Zǽ�t����N�D�x��P��͇���x׾��� �ك��   �   ���Z�쾻)⾐Ѿx��~@��Jw����^��K0�v	��Fǽ䎌���;�h�� ���D�7�l*�(Ro����������Y�<1��N���_Z齢��<v�4V(��1��J6�.6�e�1�*�ڻ����X��4��ս�N���������`*��D󀽳H���e���Žg���<!��lL���}�4�����>�ʾ`�ݾ�d��   �   tN¾����(���:���s��E���Uh�r�@�3������fʺ��'��]�F�E���
Լ⬷�v�Ǽ��آ5�L!}� ת��ݽ��	��$�B�=��S���b�C�k�z	n�,bi�k�^�ϒO��=��(�,�����9ؽ<���\ו��8z�F5X��I�V�O�p,p�t�½^?��1�!��I�l�t�
����梾𳲾`���   �   3I�����"+��|J����~���b��5E�
�'��C�Ћ�4g��7)��N�[���.�պ�lM�W@&��R��苽�+��L�򽂙�~�;�5^��F}�����г���K�����B-��[L��!�~�^�b��7E�W�'��D����Ng���(����[�h�.����I��;&�|�R�{勽v'��`�򽑖�
�;�F�]�LB}�Z���e����   �   =�k��n��^i�_�^�G�O��=���(�<����i9ؽ����ؕ��:z��7X�I�I P�91p�\����½�C���!�\�I�D�t�>���A颾�������2Q¾��������<��_u���F���Wh��@�C��$����ʺ��'��]�F�~���Լ������ǼV���5�3}��Ҫ��ݽ��	���$���=��S�}�b��   �   ˴1��G6�S+6��1�'*�d������W�e4��սpO��~���`����+������J��Sh���Ž�j���>!��oL��}�=���-���ߍʾ6�ݾ�g꾯��2��^,��Ѿw��B���x����^��L0�?
�|Gǽ���~�;���4���(�7�_*�Bo��v�����̱Y��,��b����T齛��s��R(��   �   �����
�T��U�)���@
�_���	����뽢�ٽ��ƽ�"��������B����I���ǽ�w�������D��x��R��؉��<{׾^��l�U��
\�BN����S���/�ܾ���W�����|G�3��Xؽ�T���9��{̼��0��s����:�9��`|ǻ�~�p�弸g/���q����������ڽr���   �   �K���ӽ�F�?�`O�Q"���g��2�����`�a�սBaȽc���շ�V`����˽T������5�q�f�N���2ײ���־t���ҟ�I��b$#�U?&�L�#�f�����Vx��eVپ�(��&[��S_�!#&��뽷֜�X�<�F��x�˻'�;(%<��3<p��; =�:���9������c;��r������)���   �   :���ݟ��� ��нȽLؽIp��F������.�h��1�ڽ��ҽ�(Ͻ��Խ/`轐���O$�<N��D��뀣�s{ɾ�	���H���-��H7�դ:���7��N.����܉�����Ǿኟ��qu��M5������&��2�C�ZG���T�t�<f��<�<V��<�5d< ��;��ﺰJG�M��Ls�;�@�ip��   �   8�X�����\���뱽��ƽ��ٽ�x���򽚳��`�� 򽘄�1�����'齠����� �3��`�������Z۾s�����=<-���<��0G���J��NG�/)=�|S-��R�����׾�̫������A��z��Q��K��N���3Ǻ�L<�#�<���<p3�<ʌ�<ߏ<(�*< S�:�:������z��S�)��   �   ��1��d�`���d@��ϼ����ӽΟ�*d��&L���*����������ｴ��.���{�����s=���l�$����r�����ȑ
�|!��/6�صF� cQ�U��jQ�4�F��6�&� ��T	��;�eƳ�ݘ��J�-�����sTQ�斴�@�1� �h<\��<�B�<�/�<bU�<&��<([�<��!<@�Z:���T5���� ��   �   5�$��cX�����4���غ��Pҽ1����� ��Y �
&�����b�r�}��J�������@�Cq����-���������:$�2E9�J�*�T��X���T���I�9���#���*��슶�������L�����丽o�S��^�� �㹔|q<�z�<�Q�<.��<��<&��<�ϣ<(�M<p�w;��ƻF���\O��   �   ߯1��d�г���?�������ӽƞ�c���J��)�����������������&{����s=���l�{����q�����-�
�_{!��.6���F�;bQ�2U�jQ�\�F�6�x� �%T	��:⾡ų�E��� J����$���SQ�ޔ����1��h<��<C�<&0�<�U�<f��<l[�<T�!<��Z:����4��[� ��   �   ��X�����[���걽r�ƽ�~ٽw轡��^��������?�������὜%�������q�3���`�� ��*���X۾N��g���:-���<��.G���J��LG��'=�R-�8Q������׾˫�����]�A�jy��O��V|K��J���Ǻ(�L<L%�<���<J4�<���<�ߏ<|�*<``�:�8������x��H�)��   �   N����������
�Ƚ2ؽ�m�BD�������� ����ڽ��ҽc%Ͻ'�Խ�\轎��tM$�gN�+C���~���xɾ��6��F�j�-�@F7�s�:���7�kL.��������F�Ǿ܈��knu�jK5�����#��]�C��A�� �T��<b��<x�<r��<t7d<X��;�ﺜHG��K��nr��@��p��   �   rJ��yӽ�D�#��L�s���d��������+\�p�սM]Ƚ*_���ѷ�M\����˽y��D����5�=�f�����Բ�
�־���b������!#��<&���#�ċ�D��t���Rپ�%���X��UO_�A &�Ƚ뽊Ӝ���<�t?����˻(4�;�%<,�3<(��;�O�:x��8��Y���b;�)�r�V����(���   �   #���
�/S��T����)?
����������f�ٽR�ƽ���ė��q��ŕ��&E��jǽGq������D�Fx�#O��΅���v׾���S���X�DK����!�����ܾ���T�����xG��(Tؽ/Q���9�lt̼l�0� U�`��:�����uǻP�~�*��g/�ܶq�d���O����ڽ���   �   4�1��F6�c*6���1��*�и�ؐ��U�C0�ΫսK�����􀐽h'��b����E���b��oŽc��1:!�jL��}�-���{ﲾ��ʾ}�ݾ�a꾔��6�쾳&⾶Ѿ���1>��Ju��[�^��H0���Bǽ����G�;�\��̣��|�7��Y*�>o�8u��6��&�Y��,�����jT�[���r�{R(��   �   ��k��n��]i�B�^���O�{=���(�^����A5ؽL����ӕ�@2z�F/X���H���O�S&p�$½�:��k~!�κI���t�ͅ��H䢾1���v|��rK¾����C���7��
q���B���Qh��@�N�����:ƺ�P$��E�F����� Լ����Ǽ]��A�5��}�fҪ���ݽ��	�u�$�N�=�SS��b��   �   �H��R���*���I��ұ~�~�b�V4E�Y�'�.B���Lc��@%��P�[���.�M��9D�6&��R��ዽ!#��9�򽇓���;�3�]��=}�ڌ������zF�����}(���G��X�~���b�'2E�ˊ'�.A���
c���%��	�[�	�.����(H��:&���R�"勽*'����n����;��]�B}�6���7����   �   BN¾�������>:��s��rD��[Th���@���������ƺ�X$��=�F����t�ӼB�����Ǽg��S�5�]}�Ϊ��{ݽ��	��$���=�NS���b�}�k�� n�Zi���^��O�/=�>�(�4 �)���4ؽ{����ԕ��4z�U2X��I���O�i+p���½?���!���I�L�t������梾ճ��<���   �   ���)��{)�<Ѿ��@���v����^�?J0���Cǽ苌��;���Ɵ��t�7��K*�4-o��j����ΩY�[(������N�?��`o�O(�ǰ1��C6�W'6�0�1��*�������T��/�ʫս�K��$���d���&)��j�H��le���Ž�f��q<!��lL�h�}�&�����-�ʾM�ݾ�d��   �   �Z��L�������؍ܾ�ｾ4V��.���zG�0��Uؽ�Q���9��r̼��0� 3� �: ��� Tǻ$�~�*��`/�Ѯq���T����ڽz�r��^~
��P��R����=
���������뽿�ٽ4�ƽ���^���@��З��rG��ǽNt��͐�7�D��x��P�����x׾�����Ѓ��   �   �=&��#���{��5v���Tپ'���Y���P_�i!&�=��SԜ�8�<��>����˻ A�;p %<��3<���;`Ϣ:h��-�����[;�t�r�J����$��ZF���ӽ>A��^J����c��'������\�l�ս�^Ƚ�`���ӷ�:^����˽�콧��6�5�B�f������ղ���־6���������"#��   �   ��:�؋7��M.�������`��Ǿ݉���ou�yL5�~����$���C��A��p�T�@�<���<Z!�<V��<HCd<x��;�9� 6G�pA���l�8�@��p�R���⛣����ڹȽrؽ�l�C���������$�ڽ$�ҽ�&Ͻ��Խr^轒���N$��	N� D�����zɾ7���G���-�kG7��   �   ��J��MG�j(=��R-��Q������׾�˫����5�A��y�oP���|K�K����ƺ��L<.'�<D��<�7�<���<��<��*<���:�*�����p��/�)���X���� Z��*鱽>�ƽ�}ٽ�v轄�򽒱��������7���������&�p���h��F�3���`�[������Y۾ִ���t;-���<��/G��   �   �U�~jQ�ԳF��6��� �~T	�@;�Ƴ������J���������SQ�0����~1�h�h<��<|D�<�1�<�W�<���<�^�<$�!< [:|��0��� ���1�wd�̲���>��<����ӽh���b��K���)�����,�����>�����{�Z��xs=�P�l�Å��:r����o�
��{!�1/6�d�F��bQ��   �   	�[���ύ�����0f��D���!�� � �ľ����L��������*�8�]��W�;є<,��<к�<���<V�<�Q`<��;@/1�`a?�������Q�}f8�K�T���n�gg��*s���'��.M��������{-���㚽B���ں��SQٽ���92�Qul��͜�I;�y���#�u�E���f�X*���ٍ�<[���   �   �}��/�
���T���zb��pA��`�y?������������H�p��4���w�(�ȧ\�pw�;��<�r�<���<dU�<v�<�[-<��;�ۻ�6��X�μ��F,�<�J�ͣe��J}������H�����C������\��<���%��".��b����pս�)�E/�jah�B!��j�ɾ�A��	!��hB���b����w����풿�   �   |W��T���nℿW�s���W��?8�0��fZ�㸾�7����?�2]��nϛ��U"�@\�0��;\gr<'�<T��<$҂<LI<`��:����t���Ｐp ���E�Vf�0
��!f��"7������7K��򞠽p���9~���S��fȔ��Q���=������|2ʽ�+��E&�&�\��]��綿�b���J��8�/�W��s��̄�����   �   �'��R�����t�7�`���F���)���"�޾����L_|��(2�
��⍑�Ӵ���`�@t�:�4)<U<|2<H�;�h����t���ݼ��"�_�T�H����������|^��J	������z뼽����\q���Ȭ�����l����>���j���J�S���� 轚��&�I�->��f������R����)�9�F�3`���t�/׀��   �   ��i��f�O�Z�FxH��1�_������%�ǾӔ���Xc�L!�%�׽mw���	�LXr��*���n;��c; _���4�pt��86��']��r��ᜮ��ʽhG���D�����Z���"D�)���5ӽ�½
C��=!��Lv����������4��:Т���˽���>^2� �m�	���<Ⱦ���<���0���G���Y��e��   �   h�I��sF�4�<��6-�ٕ����Ǩپ ��xQ��V�G�j�ŏ��	�r���
����I����LL�����6J��u��@k��/8㽾z��k��?#�g0+���-��+�%���%����}���Ľ[z���B������Ap���t����������ὰ����J����������f־��p��ð+���;�f�E��   �   �-(��%����X��� �nݾ\񷾘Γ��e��*,�����|n��T+^���	����v݀������Ѽ�"�q�p�v����ݽzh�<{'��1A�K�V�2�e��4n���n�K\h���[�ͺI�۰4���m4���⽊���&���}��T\��/R���c����u������gS&�8#\���������U׾�O��Y���#���$��   �   t��`���������\ҾC���>ؗ��v�cA�Ԇ�s�ֽĝ��r5P������ۼH�Ӽx��8����5���i���/ ��E�8j�D˅�#r���䜾fY�����������c��uւ��gf��eE���$�� ��Oս����j���8O��4���5�LV�@9���J���h��*.���a�V���4���7�ʾğ�6h������   �   WyԾ�VҾJfɾ`���o���Dő��-v���I�A� �����^��|���e�J�c�l��#�]I�"7��-���P�DV,��4Z�X:���1f����þ�~Ͼ�|ԾZZҾviɾ:���凧�NǑ�01v�0�I�� �L���������Y�J�.�� �@XI��3���}��mM��R,��0Z��7��0휾c��r�þ?{Ͼ�   �   rV��ȁ������sa��jԂ�]df�:cE���$�4��Mս����"��+9O���4���5��OV��;��N�� k��-.�vb����劬�T�ʾ@���k�����o��L�����뾎_Ҿ����ڗ�Yv�qA�<��;�ֽ�����5P�	��,�ۼZ�Ӽ@�t�8�T�����9d��9, ��}E�g3j��ȅ�Po���᜾�   �   0n���n�	Xh�}[���I�1�4����2����L��E&���}��U\��1R��c�
��H��������U&�Q&\�r������{X׾�R��6���%���$��/(��%�����V� ��pݾ[�"Г�Y�e�P,,������o��H,^�F�	�Z���؀��~��TѼ��!��~p�����ݽe�bw'��-A���V�s�e��   �   �,+�3�-�ж+�&%����&����L�ὤ�Ľ�y���B��:��Cp�˕t����� ��G�὆��N�J�2�������Qi־�������+���;���E���I��uF��<�N8-�Z�����̪پ����R����G�k����K�r��
��틼�� �83�����jB����*/J�
q���e��2�ew��g�<#��   �   X���N���$����@�P���3ӽ½(B��� ��\v��`���� ��.5���Ѣ���˽Л��_2�`�m�x
��Y>Ⱦe�����<�0��G�z�Y���e�r�i��f��Z��yH��1����������Ǿ啙�NZc�Q!�^�׽x���	�DVr���Po;P�c;��Ẑ�4��h��-/��]�@n��ؗ��Dʽ�A��   �   7����Z�������鼽�����o���Ǭ�����P��$󑽲������8󜽗���p轲����I�!?������=��K����)���F��4`�R�t� ؀�](�����<�t���`���F���)�f�T�޾�����`|��)2���t���,����`����:�:)<|#U<h#2<�0�;�F��x�t�^�ݼ$�"�H�T�����2����   �   nQf���,d��o5��5���(J��;�������~���S���Ȕ�R��->��B���`3ʽ�,��&�:�\��^��׷�������\�8�*�W�!�s�_̈́�����X�������ℿG�s�g�W�L@8����:[�,举Z8��y�?��]���ϛ�V"��\�x��;�jr<�)�<���<�ւ<�S<@�:��fl��@y�l ���E��   �   D,�f�J�2�e�II}�y���5H��⦕�(������m���<��&��b.������qս<*��/�bh��!����ɾHB�
!�XiB�@�b����ǈ��5�}��y�M������>{b�qA�8a��?��-���⸎�/�H����N�����(�\�\��y�;^�<�s�<���<�W�<�x�<�a-<��;Xvۻ�2��μ}��   �   �Q��f8���T���n��g��ns��(��]M��/������x-���㚽6���̺��NQٽ���%92�kul��͜�7I;�y��#���E���f�`*���ٍ�>[���[���ύ����l0f�ϛD���!��� ���ľ�����L����V��z�*���]�pX�;є<��<���<b��<"�<DQ`<���;021�|b?�r��T���   �   �C,�ׁJ�~�e�oH}�􉈽�G��6���q���� ������;��$%��v-�������oս�)��/��`h�� ���ɾ�A�R	!��hB�H�b�d��1����풿6}���񒿸������Kzb�ApA��`��>��W���C���D�H���_���,�(�|�\��~�;H�<�t�<��<�W�<�x�<@b-<`�;uۻ,2���~μ#��   �   �Pf�{���c���4��>��I��򜠽�����|��<R���Ɣ�ZP��i<��P���41ʽ*��y&�3�\�9]��'���m�������8�R�W��s�Ā�ߋ��V����ᄿ=�s���W��>8�p��-Y�⸾(7����?�W[�� Λ�S"�l�[�x��;�nr<
+�<���<Pׂ<TU<�$�:����k��`x＊k �I�E��   �   ����+Z������缽*���:n�� Ƭ�j�������R��������𜽆������{����I�Q=��P���F��w����)��F��1`�:�t�`ր��&��~���+�t���`�u�F���)���~�޾k���7]|�/'2����苑������`�`��:�?)<'U<�%2<P4�;@C����t���ݼ��"���T�3�������   �   ��0��7��������>�r�⽿1ӽ�½�?��D���s���~�������1��΢�x�˽#���\2��m�����:Ⱦ�����3�0��G���Y��e���i��f�i�Z��vH���1����\���5�ǾE���XVc�a!��׽u����(Jr���
�P"o;`�c;`��H�4��g���.�:]�n�������ʽcA��   �   \,+���-�:�+�j%����!
���������Ľ�v���?����n<p���t��������f��Ո���J�0���ԣ���d־��������+���;�N�E�A�I��qF�&�<��4-� ��:��9�پ�����O����G��g�^�����r�T�
�&狼\� �0&��<���@��?���.J��p���e���1�:w��g��;#��   �   �/n���n�rWh�V|[���I�+�4����1���_��7#����}�O\��*R���c���3���=���Q&�: \���l����R׾LL������!�g�$��+(���%����j	�� ��jݾ�x̓���e��',�s����j��^%^�V�	�f
���Ӏ�`{���Ѽ��!�~p�f����ݽ�d�<w'��-A��V�.�e��   �   JV����������a���ӂ�ecf�!bE�[�$����Jս����|���2O�_�4�P�5�6FV��5���F��~f��'.�0�a�#�������(�ʾP��nd�����f��U�����"��tYҾ`����՗�d�u��A����ֽ���:/P�B��r�ۼ��Ӽ��U�8����D���c��, ��}E�H3j��ȅ�8o���᜾�   �   6yԾ�VҾfɾ�������đ��,v���I�� �f����������6�J�����p�RI�F0���y���J��O,��,Z��5��nꜾ�_���þ�wϾ�uԾHSҾ�bɾ���o�����e)v���I�� ��������Ҳ�� �J��������VI�h3���}��IM��R,��0Z��7��$휾	c��^�þ%{Ͼ�   �   h��N�R������v\Ҿ囵��ח��v�W
A�����ֽ:����/P������ۼ·Ӽ~���8�Z�����d^���( ��yE��.j��Ņ�dl���ޜ�ES���~��蛚��^���т��_f�)_E��$�F��Hսo����{��3O��4��5�(JV��8��J���h��*.���a�J���)���,�ʾ���(h������   �   �-(�ٴ%����?��� ��mݾ�4Γ�<�e��),�����Sl���&^�Q�	����8π�ft���
Ѽ��!�ovp����#�ݽ�a�is'�<)A���V�V�e��*n���n��Rh�Cx[��I�8�4�/��/�����
���"����}�&P\��,R���c�2��򭶽����ES&�#\�s��������U׾|O��V���#�~�$��   �   c�I��sF�(�<��6-�ĕ������پ����"Q����G�6i����7�r���
��勼P� �0�� ���6�����&J�6l��J`���+��s�d��7#��(+���-���+�@	%�������(��0�Ľ�u��L?��V���=p��t���������Ὅ����J����������f־��m����+���;�c�E��   �   }�i��f�H�Z�=xH��1�K�������Ǿ����=Xc��!���׽�u��@��Hr�P�
��Co;`d;�Q�Ԣ4��[���'��]�Pi��X���Nʽ�;������}������:���%/ӽ�
½�>������s���~��_���3���Ϣ�l�˽^��$^2��m����|<Ⱦ���;���0���G���Y��e��   �   �'��P�����t�1�`���F���)�����޾�����^|�Y(2�
��̌��b��X�`� ��:�E)<�/U<,12<hP�;� ��<�t���ݼ�"�9�T�4����{��x���&V��S�������伽����hl���Ĭ���������Ћ��b�����ջ��z �}���I�&>��b������P����)�8�F�
3`���t�/׀��   �   }W��T���nℿU�s���W��?8�'��PZ�w㸾�7����?��\���Λ�6T"���[����;$rr<�-�<P��<܂<�`<`��:ܧ��b���n�If �ϛE�Kf����a��b2��L}��vG������Α��|��R��%ǔ��P��=�����(2ʽH+��4&��\��]��䶿�^���I�~�8�-�W��s��̄�����   �   �}��0�
���T���zb��pA��`�n?������������H�I��ܫ����(�,�\�@��;(�<�u�<��<FZ�<�{�<hi-< �;�bۻ-��$yμP��@,��~J�Ξe��E}������F����������� ������;��l%���-��(���zpս�)�=/�bah�@!��i�ɾ�A��	!��hB���b����w����풿�   �   ��̿ZVɿ�]���ǯ���������T�\�
�/�r����ƾd�����=�D��=��~���X��� %<"��<�*�<�d�<XI<p�;�� �U��[��T�����k�/���@�� L��eQ��Q���M��G��>�M�6�uv2��7���J��t�����۽AY�{TY�p_��*�ξg�	��1� Y^�E+���V��M����l��Wɿ�   �   m�ɿ�'ƿqY��������t��`"Y���,��u�7kþ�]����:�����5��C����ƻ�v<��<M�<��t<ı<��Y:\^�И��"�^��8�2���I�PZ�	�c���f�"�d���]�h�S�:)H�f7=��t6���8���I�Ir��m��i�׽t���U�ɔ�P˾�d�2�.�	�Z�c���Q̙��!��q\��O"ƿ�   �   !��9漿ᐳ��O��҄z���N�ߔ$��Q��4,��nރ�	2�W$�Fu����� ��ȡ�;��><�<<Ȫ�;@��P18�4���L��9��a��Ȁ�ȑ����������d��D���!���z�f�e�� R��C�g�=��]H��j������̽���j�J��G�����:� ��J&�*�O��!{�=j��+䤿�t��;м��   �   �G���b���ǥ�(A��S���g�J�>����S��ʫ���s��$�^~н��o���T��k�:8j�;@IV:ؿ�|�������?�~�{��-������_MŽ|ѽ�ֽ�@ս��ͽd���x��.�������w�C\Z�m�H��G��_��2��컽:��'�9������>���C�W��=4?�g��܆�����䂥�X7���   �   �b���՛�"&���	��23q�:UN��@*�z���Ͼ����'Z�ɧ����&\�~�h
O�h�ʻP��(o��ܼW�0�;J}��h��$�Ͻ@�����	�U]����-����9������~ҽ�8���җ��*���[�oK���S���|�Kߦ�{��$��he��!��եѾ���L�)�@�M��Kp�����N��������   �   �㈿�����H2k��xP�DS2�|/�q꾥$��6k����=�:�.���I���d-��BL��h�����a`[�'P����н:�̓�T8�z�L�r[��Cb�/�a�gQZ�qL���9���#������꽮꿽������z��V��K��2b��珽NƽZ���C��w��,���<����L�0��N�o�i����g���   �   H�d�6a�p*V���D��b.��C�v���d�ľǬ��Oka�) !�`�ܽ4����9����+ѼL7�jd*���z�����^��"8��B���g�ax��0��tA���g��"-��"ϗ�����}�FC]�>4;�C��!���8ܿ�NT��<�j�XJ�/K�
]r�<������D� �H�]�v�������$Y���Z9,�P�B�!�T��v`��   �   D�8��5��+-�*��J��P��Ⱦ#Ơ���x���9����fW��&�}� ^1�U�����"�;�JX��	9���w��y.��Q^�*;���Π�������Ⱦ��Ծ��پ�V׾��;����驾�����Pv���G�Lg�L�𽷢���Յ��Q���9��8I��逽(f���b��U�/�j�l�?��'"¾l��Hl
�����{+��5��   �   5.��9�|��ȟ���&޾�#��|��r����G��n���۽T휽�;b�E'1�&8'�.E��酽�Խ�����4�V3m��䕾���Y�־K�󾆅��1��0��;����̣��h*޾�&�����L����G��p�4�۽��<b��&1�6'�R*E�煽�н����4��.m�╾¯����־��:���/��   �   o�پ�R׾��;#���橾V����Lv�|�G��d�
�𽚠���ԅ��Q���9�&;I��뀽Vi���f��L�/�O�l��A��6%¾��gn
���G~+��5���8���5�.-�],��L��S�Z�Ⱦ;Ƞ���x���9�U��DY����}�3^1����p��>�;��T��d4��t��u.�.M^�e8���ˠ�������Ⱦ��Ծ�   �   �d���)��̗� ����}�H?]�1;����o����ٿ��R����j�WJ��K�`r�����!�余� �k�]���������i\����;,���B���T�{y`�&�d��8a�-V���D��d.��E�T�����ľs����ma��!!�w�ܽP��6�9���� &Ѽ./�^*�:�z�������Q4���B���g�xu�� ��,>���   �   c>b�5�a��LZ��lL��9���#�/�����翽ۓ��W�z��V���K��4b�8鏽�ƽ��w�C��y��B�����辏�D�0�J�N���i�d��h��d刿M�������4k��zP�U2��0�Ys�R&��ll��1�=�J�`��bI� �鼴)���E��$��v��UX[�,K����нu6����O8���L�[[��   �   L���)�+����;�^���zҽ�5���З�N(���[��nK�e�S�v�|��ঽ]}�b$�-ke�#��̧Ѿ����)��M��Mp�%�������B���7d���֛�R'���
��5q��VN��A*�{���Ͼ�����(Z�ƨ����'\� �`O�P�ʻ����n���ܼ��0�A}�\c����Ͻs����	��Y��   �   �vѽҲֽ�;սl�ͽT`���u���~��1���.w��ZZ���H�)�G��_�^3��]�3����9������?��FE�i���5?�� g��݆�����񃥿m8���H���c���ȥ�B����+g�\�>�x������ʫ�ʍs���$�Vн��o��������:X~�;@%W:؛�v�N��!�>���{��(�����HŽ�   �   z����������8b���������z�%�e�A�Q��C��=�^H�Dj�J����̽d��s�J�SH��� ��ޥ ��K&�%�O�(#{��j���䤿ku��Ѽ�����漿�����錄�O����z�~�N�r�$��R���,���ރ��2��$ὒu����Ｐ��p��;��><�#<<���;����l 8�T��������8�9a��ŀ��   �   ٿI�mZ�b�c�;�f��d�׻]��S�<(H��6=�Nt6�ޞ8��I��r�-n�� �׽���U��ɔ��P˾/e���.���Z������̙�"���\���"ƿԄɿ$(ƿ�Y��T��)����t���"Y��,��u�rkþ�]���:����6���B����ƻy<��<&O�<��t<��<�GZ:U�~���p�X��$�2��   �   ��/�>�@�BL�]fQ�r�Q��M�+G�<�>���6��v2��7�	�J��t����۽WY��TY��_��M�ξ~�	�9�1�Y^�S+���V��Y����l��Wɿ��̿SVɿ�]���ǯ�����v���6�\��/�X��s�ƾB���^�=����<�����(���@%<D��<�*�<�d�<4I<�o�;��T�U�:\������B���   �   ��I�Z��c���f�m�d��]�J�S�M'H��5=�)s6���8���I�'r�Dm����׽!���U��Ȕ��O˾�d���.���Z�(���̙�U!��\���!ƿ�ɿV'ƿY��������9t���!Y�U�,�3u��jþ&]���:����(5���@����ƻ({<n�<�O�<H�t<8�<@QZ:xT�6���(�*����2��   �   2���*���C���a��\�����n�z�U�e�L�Q�\C���=�n[H�Pj����R�̽�����J�G������� �J&�^�O�!{��i���㤿�s��yϼ�X��o弿���>fN����z���N��$��P��2+���݃��2��"��s��R�� ��ز�;�><�%<<���;����x8����������8��a�nŀ��   �   [vѽW�ֽ(;ս��ͽs_���t���}������c	w��WZ�U�H�p�G�|_��0��D껽6���9�Ґ���=��+B�m��3?��g��ۆ�����健�H6���F���a���ƥ�-@��o��Lg���>������辺ȫ���s���$�|н�o������ Ϗ:8��; QW:�廨����>�v�{��(��T���GŽ�   �   ���)�Ո������%��yҽe4���Η��$���[�IjK�[�S�n�|�ݦ��x�;$��fe�G ���Ѿ�����)���M��Ip�ኇ���������a��Aԛ��$�����1q�bSN�?*��x���Ͼ ����$Z�������!\�����N�p�ʻ����n���ܼ:�0��@}�/c����ϽH�����	�cY��   �   +>b���a�cLZ�glL���9�3�#�p��^��濽Ց����z��V���K�.b�叽gƽ�����C�}v��H������g�x�0���N��i��%f���∿����D���/k�HvP�FQ2��-�bn�{"���i����=�:���DI�x���#��B���������W[��J����н^6���vO8�w�L�1[��   �   fd���)���˗�����-�}��>]�D0;���������׿�|P����j��	J���J��Wr�&������� �J�]�����e���V��/7,���B�v�T��s`�e�d�@3a��'V��D�4`.��A������ľ�����ga��!�2�ܽ�����9�J���4 ѼB+�N]*�R�z�m������84�k�B���g�mu������>���   �   X�پoR׾Կ;����橾���9Lv���G�d���t���B҅�ZQ���9��2I��怽xb���]��n�/���l��<��<¾���:j
�V��-y+�25���8�R�5�)-��'��H��L�v�Ⱦ�à���x�H�9�0��:S��H�}�X1�������P�;�2T���3��Xt��u.�M^�\8���ˠ�������Ⱦ��Ծ�   �   -.��9�l�������&޾�#��+����+�G�n���۽뜽w6b�!1�p0'�<$E��ㅽv̽�5���4��*m�aߕ�������־�����-��+�*7�"��e����"޾� ��������G��k���۽J霽�4b�,!1�-2'��'E�7慽.н�����4��.m��ᕾ������־��6��z/��   �   ?�8��5��+-�	*��J�fP�e�Ⱦ�Š��x���9����uU����}��X1�k�������;��P���/��q�>r.��H^��5���Ƞ�j�����Ⱦ��Ծ3�پ[N׾��;a���㩾`����Gv�F�G��a�k������Ѕ�jQ���9�!5I��耽ge��b��,�/�O�l�
?��"¾e��Dl
�����{+��5��   �   F�d�6a�i*V���D�pb.��C�@���&�ľ~����ja�u!���ܽB	����9�����Ѽ�#��W*��z��������0��B���g��r�������:��a��{&���ȗ����!�}�W:]��,;�,��v����Կ��N���j�T	J���J�+Zr�H������ �'�]�k�������Y���W9,�N�B��T��v`��   �   �㈿뷆����@2k��xP�4S2�h/��p�m$���j����=�������I�4��� ��$<��������P[�F����н�2��{��J8���L�
	[��8b���a��GZ��gL���9���#���� ���⿽����c�z��V�2�K��/b�~揽�ƽ����C��w��#���5����J�0��N�o�i����g���   �   �b���՛�!&���	��*3q�0UN��@*��y���Ͼ^����&Z�E��\��#\�����N� �ʻ���,�n���ܼ��0��7}��]����Ͻq���R�	��U�.���%�/��[����(��quҽ@1���̗��!���[��iK���S��|�lަ��z轝$��he��!��ΥѾ���J�)�>�M��Kp�����O��������   �   �G���b���ǥ�'A��Q���g�B�>����6���ɫ�8�s���$�z}н��o�z����� �:���;�'X:8u��䕼y��$�>���{��#��z��VBŽ�pѽ�ֽ�5ս��ͽF[��5q���z������0w�UZ�H�H�[�G�%_��1��d뻽���9������>���C�T��<4?�g��܆�����傥�Y7���   �   #��;漿㐳��O��τz���N�ٔ$��Q��,��Tރ��2��#Ὂt��(��X�����;�><\.<<x��;�*��L8��������i�8�"�`�����������������^����������z�j�e�5�Q�C��=�s[H��j�
�� �̽���W�J��G�����8� ��J&�'�O��!{�<j��,䤿�t��=м��   �   n�ɿ�'ƿqY��������t��^"Y���,��u�-kþ�]����:�L�뽙5��\A����ƻ�|<��<�Q�<��t<8�<@�Z:�J�������ú�]�2��I�|Z�z�c��f���d���]�D�S��%H��4=�~r6�R�8���I�zr��m��6�׽c��t�U�ɔ�P˾�d�/�.��Z�b���Q̙��!��p\��Q"ƿ�   �   ���v��"������mL˿U����Ր��`g��1�I��V㺾jf~��=$���Ľ�yN��ȡ���U�0�<d�><P	<��.;�Ȼv7���Fؼ����g5���O�e�`��h�&kf��r\���K���6��]�P 	����0�߼�_�hO�ջY��%���E����:�����߭¾G��=�4���i�֑�	x����˿t��k���p���   �   ���z� ��������&ȿ����t���c�c���.��_��ݷ��Pz���!�����DL�룼�w�Hb�;��<8��;`o���r5�Щ�����T1��[U���p��������`ӂ��&y�FSe�e�L�.�1�"p��P����d������+X�^ɡ�����b7�45���^�����.�1���e��s��������ȿ�Dῗ����� ��   �   ����v��&�`�ֿ�������⇿��X��&�u\������qn�z��,��tZF�8B��(��`��:@]�:���LUd��Tּ�;"���Y��?��f���Nt���������Ʋ�����Qҙ��臽v@i��C�L�#��_��-
��o��!T��%���5��,.�Q�~�IƵ�A���U�(�=�Z�s����l��~"��<�ֿ�U鿫U���   �   ې���	�׿b�ƿ̌��������z��H�ƒ�U�]e����[�\n�ˇ���>�Ĥ��|B*����`=:��"��o��ePU��������6Jսl���+��P�����/��\��_�ݽ[½�����E����]��6�n�"�=(�.�O�1o���׽�����i��Ԧ�<(羐��	I��_{�#���;X��=ƿ�׿���   �   �lο�.˿^���ܱ�����~��|
`�{2����!�ʾ���:�D�����Ai��D�7�J/ּ�����W������H<�4���)����n��>-%��7��`D��fJ�XZI��A��3�z�!� ��n��\+���白A�s�eI���9�zM�qU��z�������RO�쓾�; �	��2�
�_�F!��w��e6�������ʿ�   �   ��,��N���_$���ֈ�mij�͘A�-�Ɍ�z���My���*�2�H⍽p-4�d,�(����7�p�b�I��D�ݽ���{�3��vV���u�}��b��϶���J�����Hw����g��1H�cv'�V��\5ս^u��A��:V��Q��w��������t�1�7W}��ȯ�.L�����@��h������E��������   �   =����������,&��ee��D�x�!�_� �V�ž���7`Q�-�����2��RX7�,�!��T:�db}�XZ������Y�%��FT�nn���;��e���R���x̾�Ѿc�ξ	ž����-ɡ�H���g�ۤ:�v�~�ܽ����u$��Y]�g��w��ƞ˽���*[Q�zw��K�þ.��� �B�C�b��������EE���   �   ��r�Fo�.�c��Q�Ug9������n�о_�����n�+��?�Q죽�+k��cC��M�|���H����ؿ1��j�aT��#���DվG4�V��[��Q�cS���c���<�۾f���B{��Y�z�RMB�@����ս���r�t�xv^���y��M����*�&��h����{̾�n ������6���N���a��[n��   �   ��=��;��2��#����}���w;���"3}�e�<��������*����_�o�Y��T���γ�����c�1�vq�{���F�ƾ�&��!��@0�(,:��=��;��2���#������5{;p���6}�2�<�ҋ�����+����_�b�Y�~R��6˳�������1��q�������ƾ��-$��!��=0� ):��   �   6O��P�i��ђ��>�۾����x���z�JB������ս0����t�w^���y�BP��k"��&��h������̾�p ����M�6���N�V�a�F_n�4�r��Io�t�c��Q��i9������L�о������n�I+�EB���3,k�+bC���M��|���D���� �1�j�YQ��`���@վ�/�ı�eX��   �   fѾ�ξ�
ž�����š�aE����g�V�:�es���ܽ���#��EX]�&g�Fy����˽��� ^Q��y�� �þ����: ��B�5�b�]!��I���G����q���r����'��&"e�D�c�!��� ���ž�����bQ��.�6�������W7�z�!�P:�X[}��U��m���V�%��AT�xk��48������(����s̾�   �   g���YG��]���mt����g�r-H��r'����;1սnr��W��8V��Q�,�w�l¨��"����1�7Z}��ʯ��N쾰��׎@���h�[���bG���eï������-�������%��8؈��kj���A�� ���"���lOy�/�*���㍽,-4�p*�����R2���b�>����ݽ�����3�~qV���u��y�����   �   �aJ�nUI�n�A���3�Ř!����C��F'��p䙽��s��I���9�?zM�LV��,�������TO��퓾�;j�	���2��_�w"��qx���7������:�ʿ7nο%0˿�_��ޱ�,�����4`�z|2������ʾ�����D�����j��U�7��,ּJ�N������@<�b��$����p���(%��7��[D��   �   M�*��l,��V��6�ݽ�V½0����B��z�]� �6���"�t<(���O�p��׽���B�i�֦��)羭�+I��a{�&���_Y��]>ƿ��׿s��=��o��I�׿��ƿ͍��{���R�z��H������8f���[�o�t����>�ܢ���:*����H,:����{���GU��z��T���Dս¿�p(��   �   ��������²�J���ϙ� 懽 <i���C���#�^��,
��o�j"T�p&���6齮-.���~�;ǵ�����.�(�M�Z����Zm��W#��*�ֿ�V鿭V������w��
��+�ֿ����n��Aㇿ��X���&�F]��D���rn���0-���ZF�A��x�����: ��:����tCd�FJּT5"�hzY��;��6����o���   �   ��������т�5#y�\Pe��L�*�1��n��O� ������f,X��ɡ�z��Zc7��5��:_��a����1�$�e�Gt������-�ȿE� ���Ҫ ������ �����M�8'ȿ1���������c��.��_��ݷ��Pz���!�9����DL�L꣼ a�`j�;8�<���; )��(h5�����}�Q1��WU���p��   �   ��`� h�wkf��r\�8�K��6��]�� 	�L��߼`�O��Y�&&���E����:�Ԉ���¾b��^�4���i�#֑�x����˿���v���r�����p��������XL˿@����Ր��`g���1�-��)㺾&f~��=$�p�Ľ�yN��ȡ���U���<t�><l	<��.;�Ȼl7���Fؼ���h5��O��   �   ���}���_т��"y��Oe�h�L���1��m��N�X���\���*X��ȡ�4��zb7� 5��a^��̀��1�)�e��s��>���Z�ȿ3D�"���M� �h��4� ����i�m&ȿ�������Ĭc�J�.� _�*ݷ��Oz�ߡ!�%���.CL�X裼�M��m�;p�<X��;�$���g5�����j�Q1��WU���p��   �   o�������²������Ι��函�:i�U�C�G�#�c\�+
�Bm��T��$��f4�,.�R�~��ŵ�T�����(�o�Z�񅈿�k���!��i�ֿU鿱T������u��-~�t�ֿ9�����$⇿��X�+�&�*[�����vpn�m�+���WF�@=��������: ��:����tBd��Iּ"5"�=zY��;������o���   �   �L���>,�bV����ݽV½k���B��x�]���6��"�S9(�ɒO�~m���
׽���	�i��Ӧ��&羨��I�`^{�B���4W���;ƿ_~׿���v�濷�⿲�׿"�ƿ��������7�z�fH������d���[��l�����4�>�����T3*����L):�������GU��z��;����Cս���\(��   �   {aJ�FUI�:�A���3�o�!����[��:&��D㙽@�s��I���9��uM�>S��������PO�C듾�;�	���2�>�_�3 ���u���4��������ʿ�jο�,˿}\��>۱����~}��y`�yy2����%�ʾ
���D������f����7� &ּ(똼4L��" ��L@<�,���#����c���(%��7�x[D��   �   X���DG��B���Ht��2�g�-H�lr'����/ս�p������3V�\Q�szw������_�1�wT}�ǯ��I�^����@���h�����9D��b릿Ͽ���B*�������"��hՈ��fj���A�k���\����Iy�A�*�v�6ߍ��'4��&������0���b�������ݽ�����3�nqV���u��y������   �   YѾ �ξ�
žԟ���š�*E��'�g� :��r�2�ܽT���� ���R]�?g��t��B�˽i��RXQ��u����þ����	 ���A�v�b�'��Ϻ��uC��b��̵�������$��ke�D�J�!��� ���ž픒��\Q��*������ ��2R7�ڜ!��M:��Y}�U�����8�%��AT�qk��,8������#����s̾�   �   0O��P�]�������۾з��Cx��y�z�pIB�,��
�ս&�����t�Rp^���y�2J��4�e�&�5h�����q̾m �;����6���N���a�KXn��r��Bo�̛c��Q��d9�=�����о����yn��+��:�Y製�$k��\C� �M�l{���C����ٻ1��j�OQ��Z���@վ�/�±�bX��   �   ��=��;��2��#����}���w;����2}���<�$������>(��s�_�"�Y�O��ǳ�v�����1���p�ڝ��J�ƾ���!�-!��:0��%:���=��;��2�9�#��xy��>t;���T.}���<���
����&����_���Y��P��,ʳ�������1��q�������ƾ��-$��!��=0��(:��   �   ��r�Fo�(�c��Q�Eg9������<�о"����n�v+��=�:ꣽ�%k�(\C��M��x���?����=�1�Tj�lN������<վ�*�:���U�sL��M�˒�������۾9���Pu����z��EB����d�ս�򜽒�t�Np^���y�ZL�����&��h�����p̾�n ������6���N���a��[n��   �   =����������(&��Ze��D�g�!�J� �'�žؖ���_Q�_,��������
R7���!�rI:�RS}�uP�����d�%�$=T��h���4��é�����^o̾�Ѿ��ξ�ž ���_¡�DB��`�g���:��o��ܽj���.���Q]��g��u����˽<���ZQ�iw��A�þ'��� �B�C�b��������FE���   �   ��,��N���]$���ֈ�dij���A�����N����Ly� �*��
�^���I(4�i%�h����+�o�b� �����ݽ�|�O�3�:lV�˩u��v������篓��C�����Pq���zg��(H��n'���c+ս�m��j��~1V��Q�c{w�I������,�1�W}��ȯ�%L�����@��h������E��������   �   �lο�.˿^���ܱ�����~��s
`�{2������ʾ[��ϠD������g��;�7�V$ּX昼\D�������8<����<�����x��\$%�I�7�rVD�_\J�=PI�lA�"�3���!�0�����!���ߙ�V�s�[I�X�9�RuM��S��f���-��VRO�p쓾�;�	��2��_�G!��w��f6��	�����ʿ�   �   ې���	�׿a�ƿ̌��������z��H����;�>e����[��m������>�Ĝ���,*�h��@:���n���?U��u���󳽲=ս���$�dI����(�,P���ݽ8Q½n����>����]�l�6���"�I8(�ǒO�
n���׽h��a�i��Ԧ�6(美��	I��_{�#���;X��=ƿ�׿���   �   ����v��'�_�ֿ�������⇿��X���&�f\������qn�9�
,���XF��<�������:��: ݉�1d�L?ּ�."�'sY��7��Ԟ��Tk��ާ����d�������"˙��⇽�5i�5�C��#�,Z��)
��l��T� %��&5齜,.�;�~�CƵ�<���T�(�<�Z�s����l��"��<�ֿ�U鿫U���   �   ���z� ��������&ȿ����s���a�c���.��_��ݷ��Pz�_�!�ĕ���CL�|裼`@� t�;X <X��;`Ἲ�]5�t�����M1�JSU�2�p�~��B���5ς��y�JLe�D�L��1��k�M���������*X�ɡ�~���b7�/5���^�����.�1���e��s��������ȿ�DῘ����� ��   �    �'���$��u�N������eܿ����ޒ���b��+(������KgV�N����r����K��/9���$;@{�ȑ�L���*���N�*��W�߈{��̊�п���O��x���ִ���e�!qA��`�lc����������¼�$�y�d�������e��誾�(���E+�N�e�V��|k��Y$ݿ�. � ��҉� �$��   �   ��$�� "�����v�����Y�ؿ$?��2����_�mq%�b��&Z��D�R�&�ʊ����� �^���3����듻�	V��ȼ@���#L�U�{�u�����������u���4a��|ߓ�Jł���]�=4�WG�=޼�J���#м>-�q�c����������a����R��[b(���a�w葿6t���ٿ�L��Ɯ�x ��"��   �   ���t��������G���ο�����҉�T�T�����{ྫྷ����I����?��+#��;��<��b��Y���/��/�6�p��阽Fn���νA߽_b�8{�g�ܽE�˽4���	���d|��G����� ����3��%wb�V��7����V����e��{ �"�V�/ڊ�լ��kϿ&��<�����Z[��   �   �����x��6����j޿�h������ls~�X�C����ξU�����9�\8�F[����藿��ġ�h�̼���b^�Eޘ��gŽ�B�:s����j'�R,��*�wh#�G�����&1�~���1f���j�u9��!� ,��ab��r��`��i�E�����xӾ ���zE����U���r��%!޿MJ��pm��q��   �   ,��/���U��࿐ǿڈ��B���Ic�]�.�l[��`��K�|���&�V�ӽ�~��0�*������C�
����R��K���d���B:��U�A/l��{������}~�W�r��_�C�F��p*�b��l�)���f]����X�^KI���f�+˝��,�0�:��~S��v�(}/�@�c����=����ƿ�)߿�z�}���   �   �_���ݿ�pӿѵ¿�8��l���C=v��ZD�\��C'߾�-��[�S��퇾� �PZB�b�=�� j������ܽ���Ɯ=�Y�i�p���❾ロ�㷾���퐹��ΰ������g��w�w���L���#�D���ȸ������
u�"s��=���cϽEs���_�������߾���(�C��u��ړ����{���mҿ^aݿ�   �   |��������ұ�_����h��nIy�J�M��$�����^X���2���v8�����~۪�]~��Af������J�����G�#�s:X�zX��L��S
ƾᾝ������ H�Ed�B����徸�˾4{��^1��a f�=�1�\O�hXƽ���I`��Rڍ��µ�� �HA:�v@������ ����"�w'L�V�v����X���°�����   �   y��Mŗ�hy��dԄ��k�	�I�D�&�����j˾Ɩ�aX��j�<,ӽ�
������^0��O���U���*�`[f��䖾㫾�%Y������*|)��3�ڳ6��4��@+�G�Sf�xt�Z�ľ$ٜ���q�v84�	���c���	���M�������(Խe.�؃U�����nbȾ����,$��G��h�򄃿�r���4���   �   Z�q�@n�|b�lP��r8���<!��(Ͼ�1���l��*�����蠐�FΎ�󴬽����	%�Re�ᚾl9ʾ-��������5���M�1�`��m�a�q�0n��b��P��u8����X#�,Ͼ�4����l���*�<��d��,���*͎�h���r���%��Me�0ޚ��5ʾ���������5��M�b�`��m��   �   d�6�b�3��=+� D��c�p���ľP֜���q�W54���0a�����N��4����+Խ�0�I�U�����eȾ���l/$�G���h�冃��t���6�����vǗ�t{��Eք�b�k���I���&�����m˾Ȗ��cX�^l�H.ӽN��(���R.���K���P�� 
*��Vf��ᖾ����T�f������x)��3��   �   NE��a�	����徆�˾�w��t.���f���1��L��Tƽ����_���ڍ�Vĵ��� ��C:�PB��P���p��ȷ"�.*L���v����Z���İ�#��Ǝ��󸺿�Ա�Q���sj��dLy���M��$�z����Z��Y4���x8�����gܪ�n\~��>f�©��DF�����W�#�j5X�ZU�������ƾ&�M���ڃ��   �   D�������ʰ����|d���w�'�L�&�#�����δ��F���u�X!s�\>���eϽ�t�z�_�u�����߾���^�C�^u�(ܓ����|���8oҿ�cݿ�a� �ݿ�rӿ��¿s:��ݼ���?v��\D����h)߾f/��![���������XB���=��j� ����ܽ����=���i��l���ޝ�����޷��   �   �����w~�e�r���_�w�F��l*�����|��pZ����X�aII���f�̝��.꽱0�X;��HU��Zw��~/�S�c������A�ƿ�+߿�|���6��2����V���ǿ&���)C��{Kc���.�f\��a���|���&�c�ӽ�~����*�������C�M����L������	���=:���U�1)l�[{��   �   �M,���*�Zd#���O��j+���db���j�T9�n�!���+�bb��s��F��߆E�����Ӿ��|E�p��V���s���"޿�K��Hn��r�n����@������0l޿�i�������t~�j�C�����ξ�����9�J9�t[����L���\����̼�� Z^�٘��aŽ�;�Vo�k{�$f'��   �   �\��u�C�ܽ��˽�������^|�]�G�F�h� ��������wb������өV�ꤟ����M �4�V��ڊ��լ��lϿ5�����2�� \����u���d ��H��οz���!Ӊ��T����Z|�&���K I�����?��~"�r8�����U�Q���$�o}/�t�p�*嘽^i��Ȁν�;߽�   �   ,������^��Gݓ�VÂ�q�]�z�3�.E��9޼�H���"м-���c�G��������a�"�����b(���a��葿�t��u�ٿ9M����� �2"�"�$�� "�
���v������ؿe?��g���_��q%����RZ��v�R�&�Ċ��l����^���3� 2깐ړ���U��ȼ~��EL���{��傟��   �   ࿑��O������󴁽e�eqA��`�d��$���$����¼,%�ӎd�4����O�e��誾)���E+�x�e�%V���k��q$ݿ�. �(��ډ��$� �'���$��u�D��}���Mܿg���ޒ�W�b��+(�ֶ����gV� �������K� %9�p�$;�u�d��������:�*��W��{��̊��   �    ����񦽴^��)ݓ�4Â��]��3��D��8޼HG��� м�+�i�c�@���<����a�a�����b(���a�@葿�s����ٿ1L�����. ��"�p�$�@ "�j��Hv����Өؿ�>��Ў��,_��p%���뾛Y���R�p%�݉��0����^�P�3� �@ٓ���U��ȼh��0L���{�救�܂���   �   �\罫u��ܽV�˽Ŭ��.��*^|�r�G�<�� ���������tb�&�����ϧV�z������� �\�V��ي�nԬ�kϿA��������Z�@�Xt����R���F��ο���҉�G�T�,��hz�ʣ��lI���&>��? ��5���� S�>P��<$�@}/�I�p�嘽Pi����ν�;߽�   �   �M,���*�@d#�[��"���*�;��a��`j��9�&�!���+�^b��p��R���E�����<Ӿ&��xyE�2��T���q���޿�H���l��p����6����������i޿og�������q~���C����ξ+���A�9��5�Y����$�������l�̼E��Y^��ؘ�waŽ�;�Oo�b{�f'��   �   z����w~�I�r�o�_�?�F��l*����H��&{��\Y��?�X��EI�ܽf��ȝ�H*�`0��8���Q��u��{/�u�c�������	�ƿ:(߿�x�x��"�����S����}ǿc����@���Gc���.�.Z��^����|���&�"�ӽ�{��٪*�7��W���C������L��Փ�����=:�~�U�+)l�T{��   �   >�������ʰ�����^d����w�νL���#�������������u�s��:���`Ͻ[q�_�_�ᯠ���߾p��/�C�4u�ٓ���������jҿ-_ݿc]ῴ�ݿ�nӿγ¿�6��չ���:v��XD�����$߾�+��[���T�����~��SB�7�=�Aj�r��G�ܽ���ԗ=�y�i��l���ޝ�����޷��   �   KE�}a�������h�˾w��I.��]f�@�1�9L�qSƽ����\��׍����� ��>:��>��f��������"��$L�U�v�%��V���������1���p���]б�S����f��2Fy���M��$�����U���0���s8������ת��U~�9:f�_���fE����+�#�P5X�RU�������ƾ'�L���ڃ��   �   c�6�^�3��=+�D��c��o�ľ֜�/�q��44�.��L_������J��.����$Խ�+�x�U�g���x_Ⱦ���z*$�G���h�����p��q2��C��×�Lw��l҄���k���I���&��~��g˾�Ö�0]X��g��'ӽ������?,��-J���O���	*�gVf��ᖾ�����T�e������x)��3��   �   Z�q�?n�|b�dP��r8���*!��(Ͼ�1��p�l�l�*�I��^�������Ɏ�n�����꽱%��Ie��ۚ�Q2ʾT���;����5���M���`���l�R�q�>n�4xb��P��o8�I�����$Ͼ/��Z�l���*����@��윐�Lʎ�����<��p%��Me� ޚ��5ʾ���������5��M�e�`��m��   �   z��Lŗ�gy��`Ԅ��k���I�7�&�����j˾�Ŗ�t`X��i�(*ӽ��������*��G��K��l*��Qf��ޖ�Z���P�͇�����u)�*3��6���3�R:+�A��`�Sk���ľӜ��{q�R14����,\��T��5J��4���0'Խ�-���U�����bbȾ����,$��G��h�󄃿�r���4���   �   }��������ұ�]����h��dIy�>�M��$�^���4X���2���u8�����
٪�V~��7f�䥃��A�����{�#��0X�YR�������ƾ]
������uB��^�������
�˾�s��0+��of�q�1�hI�Oƽ<���[��$׍�p���l� ��@:�X@�����������"�w'L�U�v����X���°�����   �   �_���ݿ�pӿε¿�8��i���:=v��ZD�O��!'߾�-���[����ꅾ�G�~�QRB�i�=� j���j�ܽʚ�(�=�٧i�Xi��۝��{��fڷ�����G����ư�'����`���{w���L��#�����6������4 u��s�
;��"bϽ�r���_�{�����߾���&�C��u��ړ����{���mҿ`aݿ�   �   ,��0���U��࿏ǿ؈��B���Ic�S�.�`[�t`����|�(�&���ӽ�|���*�������3C�����G��Č��ˎ��8:���U�'#l��{�<���q~�.�r�΢_�:�F�9h*���z�ཧv��V����X�=CI��f�5ɝ��+꽥0��9��mS��v�&}/�@�c����=����ƿ�)߿�z����   �   �����x��5����j޿�h������gs~�Q�C��j�ξ1�����9�D7轮Y���������<����̼��{Q^��Ә��[Ž5�tk�2w��a'�I,�<�*� `#�p������$��]���j��9���!�-�+��]b�Gq����"�E�r���lӾ����zE����U���r��%!޿MJ��pm��q��   �   ���t��������G���ο�����҉�O�T�����{ྕ���sI�T���>��B ��3������F�H�����v/���p�����pd��p{ν�5߽W�p潿�ܽ`�˽H���F���W|��G�
�� �����Z���tb�k�������V����`��z �"�V�/ڊ�լ��kϿ%��<�����Z[��   �   ��$�� "�����v�����Y�ؿ!?��1����_�kq%�Z��Z��$�R��%�N���m�� �^�`�3� K�(ɓ��U��ȼ���	L���{�T���*���\���尿\���ړ�����2�]���3��A�l4޼ D���мW+�&�c�L���^����a����N��Zb(���a�v葿6t���ٿ�L��Ȝ�z ��"��   �    nO��K��o@���/�������v3߿໳��W����O�/]���˾���-(��qŽ��S�T)ɼH�/��m��,�<؝�������6���m�B������౽�<��Y���\w������������a���0����Ƽ<����`ȼ}������ݽ��3�շ��,kѾ�`��R�3��ܓ�� �2��U��,0���@�L�K��   �   R�K��G�l/=�
�,��S����!�ۿ����#���.L�R��QeȾ��z�%� ný�T���Ӽ�xV�T�*�4�x��μ.�`Y�����ߥ�@滽��ʽ0�ѽ��ϽYŽ��������R��6�M����L���fż��ټ�C����4۽#�0�@h����;����CO��Ȋ�����kݿ �����(9-�T9=�
�G��   �   �>A���=�J�3���$��R�������ѿ�ڨ�뷂��qB��
�uȾ��{�Õ��ӽ�,�W�����������FQ𼆥0�$w�W桽:�ǽL��������
�,t��~������tٽE涽L9��7�c��d-�n��h�� -�TŃ�;Խ��(�r����þ�i�E�	��� ���ӿo����}���$��3���=��   �   &z1�P�.���%�0?�rk�L鿣N¿]��6>q�h/3�����ӯ���h�B��M���@R_��������� �#$\�2뗽>�ɽK}��^?�I�0�;uC�B�O��"U�uR�EEH���7�"�0�	�FmོO��/����R�dz7�hF�A����ɽ�	��p�ҳ����5���r��ʜ���¿�Z鿆8� ��bT%��>.��   �   �B�6��A��w���lѿ�3������`W���D�&�����P���Rۭ�9n���D�9�R��-���e��;����u�&D�i��&���z���L���Ǟ�n���� �����6�q�FZN�r�)��K���ν�����B~��bm�ỉ�������hkW��埾ӥ�Z� �)X�4ˋ������п�����ʤ�Vj��   �   04	��(�(� ��]�g}ӿx��&���q�H�9���	�o�ľ�䇾��6����ϧ�4��^'���M����ѽ0��e�:���m��������H�þƧ־J$㾳�羵��6lپ�Ǿ&����ᖾ�x�C�E��������XT��)f����4I���E;�Ҵ���ƾ�
���9��p��i���鴿�ҿ�뿔 ����   �   <翦���ٿ��ǿ���𘿌O}�FJ��1���徶r��~�d�`q�i�ٽ>�� Y��9��������'N�����檾*�о�Q��C3�m��!�,a$���!��\Z�~U��X�վ�5��z%����W�ٓ!���)���P棽�o����@���f�ڇ��t.�wj��H�@{������a��kLƿӜ׿���   �   [g��Ц���᰿T֢������x���L��0#��u�������Q���u;�5�.Ž:M�����H�㽪����T��u��/d��[�?����(��$?�q�P���\� �`��]���R��A���+�������J"�������
\�� �;��x���<���
=Ƚ�}�ߩ:�I��Oҷ�����yV!��J��'u�����>��8����︿�   �   sO����������2�b��$B�! ������wþ�'��=�Q��j��A޽XѶ������ڽb����M��q�������a��k���:?�b�_�g�|���������Q��� ����������b��'B��# �޴���zþ�)��k�Q��l��C޽�Ѷ�����!�ڽ����M�o������(]�����c7?���_��|�5 ��3����   �   ��`��]��R���A�e�+�ȓ�k���������\�`� ���ߨ��F����>Ƚ����:�5K��@շ�����Y!��J��+u����EA������r�j��k���o䰿�آ�����^!x�M�B3#�my������`S��Jx;���.Ž|L������㽆��Z�T��r��a`��YV�g��G�(�.!?�q�P���\��   �   �]$���!����iW�KP����վ2���"����W���!���𽎝��C壽Dp����5���
f�����1従l���H�UC{�����!d���Nƿs�׿�����Z��jٿ�ǿ+���򘿉R}��J��3���徙t����d��r���ٽ���5W�������S���"N�����⪾�~оoL��?0��i�A!��   �   M��l��6gپ[�Ǿ���sޖ�H�x�ȉE�L�ò彴��kR���e�����yK���G;�j���ƾF
���9��q�Ek���봿�	ҿx��� �t���5	�R*�j� �`�kӿ3�����V�q��9���	�M�ľ懾��6���ϧ�����$���I��׉ѽp����:���m�,��������þ��־���   �   �Þ�����L�������F�q�/UN�?�)�>H���ν�����=~�`m�2̉�|������cmW�D矾���� �+X�ű�g��G�п��������k�D�x��.B��x���nѿD5�����abW�A����H�����P�J��ۭ�M7n�ՉD�&�R��)���_�����rq�� D��i�t#��w���H���   �   mU��oR�4@H�Q�7��"���	�dg�	K��r+����R�w7��F�&A����ɽ�
���p�pӳ����[5�r�r�̜�6�¿&\�f9����tU%��?.�H{1�f�.���%�@�2l�FM鿰O¿5���?q�`03�����ӯ���h��������Q_���=���� �\�旽��ɽ�u��;���0�pC���O��   �   \��p��{�����joٽ�ᶽ�5��Q�c�,`-�0��h�& -��Ń�Խ��(�%���*�þOj�E��	��]!���ӿ����x~�T�$��3���=��?A���=��3�6�$�S�����H�ѿ)ۨ�\���jrB���
�ɾ�ӓ{�%���ӽ�o�W������y������F���0�w��᡽��ǽW�齭��*��   �   ��ѽ��Ͻ"VŽײ��*���:��ǒM�C��8�� dż,�ټdC�N����4۽��0��h��p�;���DDO�Ɋ������kݿt��(���9-��9=���G�ʼK�t�G��/=�X�,�(T����r�ۿ_����#��/L�~���eȾ􃾔�%�nýz�T�йӼprV�D�*���x�μ*��[Y�𫊽,ܥ�)㻽��ʽ�   �   �<��j���tw�����ض��Оa��0��TƼ�����aȼ���W���n�ݽ8�3�����akѾ�`�;�R�M������2 �B��U��,0��@�P�K� nO��K��o@���/�z�����Y3߿�����W��r�O�]�t�˾����(��qŽs�S��(ɼL�/�Xl�l�,��ם�������6���m�>������౽�   �   �ѽ|�ϽVŽ�����������M���8���bż��ټKB������3۽��0�h����;T��`CO�qȊ�?����jݿ������8-��8=���G�ܻK���G��.=���,��S�\����ۿ����d#��*.L�����dȾ��ɛ%�mý�T��ӼpV�Є*���x�� μ*�m[Y�쫊�&ܥ�&㻽��ʽ�   �   X��p��{�����<oٽ�ᶽT5����c�N_-������,�ă��Խ��(�򾂾l�þi�^E��������ӿ����D}���$�\�3��=�>A���=���3���$��Q�������ѿ�٨�I����pB�X�
�dǾ���{�����ѽ���W� ����w������F𼵞0��w��᡽��ǽS�齭��(��   �   fU��oR�&@H�8�7��"�~�	�gཋJ���*���R��t7��F�
?����ɽ����p�ѳ����5�Z�r�ʜ���¿QY��7���`S%��=.�y1�2�.�x�%�:>��j��J�aM¿P���<q�.3������ѯ���h������fM_�{������� ��\��嗽�ɽ�u��;���0�pC���O��   �   �Þ�����E�������!�q�UN��)��G�Кν����r;~��\m��ɉ�̣����siW�j䟾���� �e'X�ʋ������п�������i��A�����?��v����jѿy2��ӡ���^W����侅���)�P���$ح��2n���D�_�R�+)���_��Ѕ��dq�� D��i�t#��w���H���   �   J��f��.gپM�Ǿ���Zޖ�	�x�z�E������R��xP���b������E��JC;�V����
ƾE
���9���p�&h���紿�ҿ���R �½��2	��'��� �][�:{ӿ������R�q�*�9��	�
�ľㇾ�6���-̧�z��6#���H��>�ѽD��|�:���m�'��������þ��־���   �   �]$���!����bW�6P����վ�1��t"��3�W�&�!��𽒛��n⣽*l��������f����+徒h���H�={�ߌ���_��JƿG�׿d��z	���9ٿJ�ǿ����>L}��J��/����Op���d��n���ٽ ���T��H�������"N�����⪾�~оnL��A0��i�C!��   �   ��`��]��R�z�A�[�+����L����Ә��]\��� ����*���T����8Ƚj{�צ:�G���Ϸ�����%T!��J�n$u�����<��ė��9��d��-���m߰��Ӣ�q���&x�v�L�g.#��q��蒹�NO���r;���})Ž�H��3��������T��r��V`��SV�f��H�(�1!?�u�P���\��   �   uO����������(�b�x$B�! �����vwþv'����Q�j�G?޽�Ͷ�������ڽ��6�M��l��?����X�� ��94?���_���|�����р��M�����D��9��H�b�!B�G �!���tþ�$���Q��g��<޽�̶�^�����ڽ3����M��n��r���!]�����d7?���_�"�|�7 ��4����   �   ]g��Ц���᰿R֢������x���L��0#��u��ȕ��XQ��?u;���*Ž�H��V�����=���T�/p���\���Q쾮���(��?���P�i�\���`���]���R���A�	�+�ߐ�������镓�\��� ������՞��:Ƚ�|�J�:��H��8ҷ�����wV!��J��'u�����>��:����︿�   �   =翨���ٿ��ǿ���𘿂O}�9J��1���徂r���d�xp���ٽP��dS��`���ό��XN��
��6ߪ�zо>G��P-��f��!�4Z$��!����YT��J��/�վ.��c��y�W���!�3��r����ࣽl���v��hf�����d.�sj��H�	@{������a��nLƿ՜׿���   �   04	��(�(� ��]�c}ӿu��#����q�>�9���	�G�ľ�䇾ƪ6���̧����	!��E���ѽ�}��:��m����������þ��־�������bپ��Ǿݤ���ږ��x���E�4�@�彀��N���a����7G���D;������ƾ�
���9��p��i���鴿�ҿ�뿕 ����   �   �B�8��A��w���lѿ�3������`W���%������P����ح��1n���D���R�7%��<Z���~��#m��D��i� ��is���D��������������4�����q��ON��})�aD�8�ν�𝽴5~�Ym�ɉ�.���̅��jW��埾ĥ�W� �)X�4ˋ������п�����̤�Xj��   �   (z1�P�.���%�0?�rk�L鿡N¿[��.>q�_/3������ү�2�h��������"M_�z������ ��\�ᗽ�{ɽ�n���6�ٝ0��jC�|�O��U�?jR��:H�m�7��"�ǅ	��`�|E���&��8�R��p7�bF��>��,�ɽJ	���p�ҳ����5���r��ʜ���¿�Z鿈8� ��bT%��>.��   �   �>A���=�L�3���$��R�������ѿ�ڨ�귂��qB��
�aȾ�Ԓ{�e��yҽ���W����s���﫼�<𼇘0�[w�ݡ���ǽq��{������lm�Kx������iٽ�ܶ�V1���c�!Z-�<��*�a�,��Ã�(Խl�(�Y����þ�i�E�	��� ���ӿp����}���$��3���=��   �   T�K��G�l/=�
�,��S����!�ۿ ����#���.L�N��GeȾ��K�%��mýd�T�@�Ӽ8lV�,~*���x��ͼd&�WY�n���T٥�໽��ʽ��ѽ/�Ͻ�RŽү��`������x�M�������^ż��ټWA�L����3۽��0�4h����;����CO��Ȋ�����kݿ �����(9-�V9=��G��   �   ��|��ww���h�t�R��9�j*�����XԿ�A���w�;1����1>��L��Y������P��d$���p��L祿|k����2�	8q�����̿��Oʽ�cٽֲ߽=�ܽ��нT輽Y9��B��!�P�;[�����Ǽ���
6�!�����zT�ť����B14�x�z��B����ֿ.���3��9��$S�$�h��~w��   �   ,�w���r�V8d��N�` 6����j���ѿ�����)s��X.����C����I�V��"��'����������м��+�T��̌�#⮽:�ͽ�I潒���҉����"��V�ֽ���DY����r��7��	� �d����w;�c6���o�MQ����4���6*1�Gov������!ӿ\�������6�
OO��Gd�b�r��   �   L�i�4e�d�W�2�D��T-���E���i�ǿ(��̥g���%�ju��A���@�O��b����1-��N ����N3+�Kl�������ʽWR��v��Ha���(���,�x�*���!�����,�ؽ�̭�v����K�wU$��q ��L��㛽E���72H��6����辷a(��\j�8����,ɿ����H!�h�-��qD�ԺW���d��   �   0�T���P��E���4�� ���	�}[忏���yN����U����ɁҾwҋ�E�3�g;�0���SN�;�E�Y�k��	����������9��U�6�j��y��~��{��pn��,Z��)@�+�"��{�<�Ͻ�C����x��VY�Zk�2e�����-c:�)(���վ^����W�~D��������忎�	����~.4��!E�|�P��   �   p0<�V9��/�DS!��k�`���Ϳ��������z>��6��Ỿ$#{��D$�$ؽ����,����+���8��Ϥ�g����@��l�E��}���h=��H����m��,����X��솢�ϓ���nt�-rH����Z���亽���"���֥��Z\�L�)��'���f���m	��?�󂀿������ͿQ������y ��.�ԙ8��   �   �,"��������k����׿>��|���e]�K$��꾅�����[����4н ֦����)ŽWS�;�,�0�a� "���鮾�
ξ��3 �)��<K
�5��v��p�; ҾM���K����i��3�f ���ѽz@���창Vٽq��6W_��(���*�<�$�S]�"��Y#����տ����4 ��&��-��   �   �<�>D�^  �~�%_ҿv���P���Up���8�/	�-Oľ�͈�EY<�����ͽ����Hֽ��	��9�b�x��E���̾�������3&�j�5��@�V�C���@�mc7��H(�����O��P[ѾBS��Ǿ�n�?��<�`t߽YŽ2�ӽ4>�D>�{a���fľb���"8���n��*��gz���hп��S@������   �   mp޿�>ۿ�ѿա��-v���?���s�rNB�J6��3ݾ���>U`��/�6�ѽZD޽��
� ];����>��a�IU���+�7QI�V�c�*�x�"$��l���K�����z� Ff��L��v.�H����r��&̂�Ÿ?�pQ��|��Խ�?��;�_�]7����۾a���q@�y,q���������ľ�~ϿSaڿ�   �   Z���;���㤿S����Ɔ���f���>������wѬ��Sz�Q4�����7޽�mݽ���O�1��.w�m�����微��	<���c�O"���*��5���^g��3�����q椿ſ��Ɇ���f��>������6Ԭ��Wz��4�� �S8޽�lݽ���a�1�d*w�W���ѣ����<���c� ��o(�������d���   �   �٭���z��Af��L��s.�����{��n���ɂ���?�lO�{� �Խ�A򽚁���_��9��%�۾����t@�&0q�%���#����ƾ�	�Ͽddڿ�s޿�Aۿ�ѿ~����x���A��j�s�.QB�`8��6ݾ�� X`�@1�E��ѽ�A޽@�
�sY;�������\�xR�]�+�MMI���c�u�x��!���   �   7�C���@��_7�E(����@J���VѾ�O�������?��9�;q߽�WŽ��ӽb?�MF>�Pc��_iľD��[%8���n��,���|���kп���iC�� ��|>��E�� �<쿓aҿ���yR��SXp���8��	�oQľψ��Z<�H��tͽ����Dֽ��	�ʔ9���x��A����̾8���r���/&���5���?��   �   H
��1��s�~k�j�Ѿ0���H��t�i���3�p���ѽ%>���밽4ٽ����Y_�~*���-�&�$��U]��#��D%����տ0����� (��/��."�N����Ɉ���	׿��[~���g]��L$�H�����Q�[�V��Fн�Ԧ����h$ŽP�ӏ,���a�x��U宾�ξ4�0 �����   �   �h������_T��邢�E����ht�+mH����:��Zຽ�����������u]㽣�)��(���h��/o	���?�!������ïͿ*S��$���z ���.�r�8�2<��9�t�/��T!��l�3����Ϳ��������{>��7�㻾�${��E$�oؽ��������(���3��2��*����@���l����i����8���|���   �   w�~�& {��jn�X'Z��$@���"�xx���Ͻ�?��V�x��RY��Wk�4e�����ld:�4)����վ���6�W��E���������r�	�����/4��"E��P���T�Z�P�H�E���4��	 �~�	��\忌¸�?O���U�����Ҿ&Ӌ���3��;⽐���PN�;�>�Y�Vf����h���+���9���T��j�jy��   �   ��,���*���!������ؽ*ȭ����x�K��Q$�Ao �߁L�䛽K���;3H��7���辘b(��]j������-ɿ�����!�6�-��rD��W���d�p�i�Fe�V�W� �D�2U-��������ǿ�(����g�9�%�!v�iB����@���������/-��K �n��?-+�oCl�ඞ�+�ʽ
L�����]� �(��   �    ���T������ֽ'~���V����r�J7�J}	���h���8w;��6���o��MQ�'�������*1�pv�7����"ӿ������ �6��OO�dHd��r���w�0�r��8d�j�N�� 6�:�����GѿЭ��*s�Y.�5 �k����I�P��W"��
��0��� �м����T��Ɍ�߮�ޙͽDF�ȹ���   �   ޲߽K�ܽôнh輽x9��]��k�P��[���缀 ǼГ�V6�^!��I��{T�<ť���l14���z� C����ֿ@���3��9��$S�0�h��~w���|��ww���h�d�R��9�V*����kXԿ�A���w��:1����>���L�fY��f�������#��\p���(k����2��7q�����Ŀ��Oʽ�cٽ�   �   ����T������ֽ~���V����r��7��|	���Ⱦ��v;��5��Po��LQ�l�������)1��nv������!ӿ*��P��T�6��NO�FGd�ʛr���w���r��7d�|�N���5������vѿ)���)s�PX.�*�ﾷ����I���!��������L򣼔�м����T��Ɍ�߮�ܙͽGF�˹���   �   ��,���*���!�����Ƒؽ�ǭ������K��P$��m ��L�n⛽����[1H�?6����#a(��[j������+ɿ����� ���-��pD�ܹW���d�&�i�e�Z�W�J�D��S-�d��.�����ǿH'����g���%�&t�A��¥@�7��t����--�tJ �����,+�3Cl�ж��"�ʽL������]��(��   �   v�~�! {��jn�K'Z��$@�ھ"�Rx�>�Ͻ$?����x��PY��Tk��b��n���a:�F'����վ}��p�W��C���������Ɲ	����`-4�L E��P���T�~�P���E�P�4�� ���	�Z�X���}M��m�U����#�ҾHы�{�3�~8�t���TMN�X;�0�Y�
f�����N���$���9� �T�!�j�ky��   �   �h������\T��₢�8����ht��lH�R�����xߺ��������Ƣ��TY㽌�)��&��Je���l	�j�?�����K���m�Ϳ4O�����<x ���.�B�8��.<��9���/��Q!��j�R��_�Ϳ�������x>�W5��߻�[ {��B$���׽~��Z���'��63��ם�����@���l����m����8���|���   �   H
��1��s�vk�]�Ѿ��}H��4�i���3����ѽ<���谽�ٽi���T_��&���(쾘�$��P]�� ���!����տ<�����
�%�F,�:+"��� �B�݃���׿Xk{��?c]�+I$�9��w�����[����н�Ѧ���N#Ž�O���,�h�a�p��R宾�ξ8�0 �����   �   8�C���@��_7�E(����.J���VѾ�O��4��%�?�J9�*o߽�TŽ}ӽ�;�KA>��_��8dľ���� 8���n� )��Nx���fпG��W=�����:;��B������쿌\ҿ/���N��RRp�>�8�G
	�YLľ~ˈ� V<����ͽ2����BֽV�	�x�9���x��A����̾8���s���/&���5���?��   �   鉶�٭���z��Af��L��s.�����{侨n���ɂ��?�qN�x㽝�Խ^;��|���_� 5��p�۾?���n@�)q�𚑿N���v���;{ϿN^ڿTm޿�;ۿ�ѿ����s��q=��M�s�nKB��3�0ݾA
��;Q`��,���ѽ�>޽d�
��X;�������}\�vR�]�+�PMI���c�y�x��!���   �   [���=���㤿Q����Ɔ���f��>�������CѬ�KSz�o4�3���3޽hݽ@���1�&w�n�����待���<�F�c����&�������a������i��᤿ɺ���Ć���f���>�ۜ����9ά�Oz��4�����2޽�hݽ�����1��)w�7����������<��c� ��r(�������d���   �   np޿�>ۿ�ѿӡ��)v���?����s�gNB�:6��3ݾ���zT`��.��	�Xѽ�<޽N�
��U;�|��p	��EX��O�%�+��II���c�ܙx�=��q���a���D�z�q=f��L�Ip.����8w�,k��ǂ�F�?�L��u���Խ�<�{~���_�.7����۾\���q@�z,q���������ľ�~ϿUaڿ�   �   �<�@D�^  �|�!_ҿq���P��vUp���8�	��NľC͈�MX<���`ͽ�����?ֽ��	���9�J�x�f>��5�̾����_��,&���5���?��C���@��[7�lA(�R���D��GRѾL�������?�\6�mk߽�RŽ�|ӽ�<� C>�8a���fľZ���"8���n��*��iz���hп��V@������   �   �,"��������h����׿:��|���e]�K$����G�����[�S���н Ѧ����*Ž�L���,��a���<ᮾ� ξ���- �ځ��D
��.��p��e�_�Ѿ����D����i�=�3�����ѽA9���簽�ٽP���V_�h(���*�8�$�S]�"��[#��³տ����6 ��&��-��   �   p0<�V9��/�DS!��k�^���Ϳ��������z>��6��Ỿ�"{��C$�n�׽�}�������#���.���������@���l���l����4��x��d��ܔ���O���~������Ubt��gH��� ��ں�=������졤��Y�q�)�a'���f���m	��?�􂀿������ͿQ������y ��.�֙8��   �   0�T���P��E���4�� ���	�}[忏���vN���U������ҾEҋ���3�z9�S���KN� ;�íY��a��N���Z������3�9�{�T��j�y���~���z��dn��!Z��@�v�"��t�D�Ͻp:����x��KY��Qk�`b��֗ｔb:��'����վX����W�D��������忎�	����~.4��!E�|�P��   �   L�i�4e�d�W�2�D��T-���D���i�ǿ(��ȥg���%�Vu��A����@��뽈���z,-��G ����K'+�
<l�l�����ʽ�E������Y��(���,��*��!�|���8�ؽ>í������K� L$�~j ��}L�⛽����1H��6����辶a(��\j�9����,ɿ����H!�h�-��qD�ԺW���d��   �   ,�w���r�X8d��N�^ 6����j���ѿ�����)s��X.����5���[I����!���������T�м=�Y�T�Tǌ�,ܮ���ͽ�B�������~���콘�ֽ�z�� T����r�7��y	����L����t;�|5��Jo��LQ����.���4*1�Gov����� "ӿ\�������6�OO��Gd�b�r��   �   �ז��c������fw�|�V��5��y���P��e	��ZL�������e�m�!������r!@�D���qż�����"���`�j*������x�Խ>������j1�%& ���۽Qk��D����s���6�`�	�0���v�@	U��n�� ~�ot��~���;��+O��Ǐ��k����������6��W�ıw��͉��h���   �   �����@��O߆��`r�n�R�l�2��)�s�b���ǋ�%I���
�fŷ��0j��M�����5�F����������'B�T�������н(򽺶�ί��1�����	�X����׽��YJ���9V��W"�Xn	�Z��Q[�b�������ip�b��f����K�[k���W��b1�P���3�n�S���r�����:���   �   �a���j��J�}��e�&H��b*��u�
<促ر��3��a?���s+���^`�fA�~���[�ǯ(���,�' Y��&���ľ�]����&�&�}8�ɆC�%�G���D���:��*�n�����m�Ƚ�b����m�.�@�/�<�o�2���؃��f��k������A������d�����*=�H�*��mH��d���}�FJ���   �   ��y�v�t�6�f��3Q�b�7�g���$Qӿ�b���u�}G0��+�顾�vQ����z������pj�褆�ſ�������5�-X�T�v�o����Ώ�9ڒ������6����z���\�S;�*Z� c�& ������t�}��L�������4
�alV�����p;��L2��w��a��9Կ0M��r�$�7���P���e��jt��   �   ��Z�8�V��K���9��:$��!��@�ӊ�����I[���o�ؾ*g���j?������	��I��T,��νd�#�0�bE`��k��h4���z��Gʾ2�վFھ��־�̾�㺾�����^���'f�j.6��g���׽�V��z⤽�;��sj�qC�|��-۾"8�^]\�ف������T�2��xv#���8��J�XV��   �   ��:� �7��m.��; �h��ɚ��`�̿僤��}~��9=��|��ɻ�Z�~�q,�/��~�ƽ$�Ľý���8dI�:��hإ��Sʾ�	�N� ���/�5H��������nw��;�/��H����N�.��BC�d�̽��ͽ܌���m/���������k�=��j~�3%����˿�$��b����]-�J�6��   �   ������bA�h��H��Ͽ7������T����\S��흾�,Z������:�߽P���W!���W�#(���ϻ���쾩��&)���?��ZQ���\�Q;a���]�Y�R�=�A�%O+�<9�����&������2�\��1%��^�4F彋���ؗ��[�j��j�'��s�S�7A�����ZYͿ�#���C�P���   �   /���a��m��"ܿ�$Ŀ״��i㋿�d_���+�:����J��{��z}8�B��Q��� 0��"�b�Y��L����ƾ����#��F�a�g��邿%̎�8����^�����LϏ��1����j��H�lW%�h���ɾ�x����\��$���������g�8��B�������d����*��]�����=���+¿�ڿ���l���   �   ,�ȿƿ����#˭�?��������[��l.�)����ƾ 0����O��j��{��4�����UN������ž���,���X�	��dޘ�>*���d���Hſc�ȿEƿ�����ͭ�����ۋ��s[��o.�U����ƾ12��h�O�Gl�'|��3����MRN�[�
ž���ى,���X�����ۘ�f'���a��gEſ�   �   �[������̏��/��Rj�1�H�\T%��e�"�ɾ>v���\�H}$��	���������8��D������ i��@�*�[�]���������.¿#ڿ1�Sp�����+e����� %ܿa'Ŀ'���Z勿�g_���+�����-M���|��F8����m���u.�;�!�3�Y��I����ƾ���#���E���g�炿xɎ�m����   �   �6a�	�]���R�5�A��K+�06�����"����Ҝ\��.%�]��D����0����[�7l��6m�P��O T�C������[Ϳ�&�X��pE�0��x�����C�����J�PϿ9��������T�����U�|�.Z�k��q���߽�K��CT!���W��$���˻�D�쾀�	#)�j�?�bVQ���\��   �   �D�t��p����q���;,��E���N�����>򽸕̽ԗͽҍ��xo/����=��)	���=��m~��&����˿9'��܃���l_-�D�6���:��7�xo.� = �ƈ����M�̿t���,�~��;=�~�5˻�h�~�r,�;/���ƽ��Ľ���T��/_I��6��Xԥ��Nʾ��	�����+��   �   �@ھ��־�̾^ߺ�����i[���!f��)6�bd���׽2S���ऽ*;��k��rC�r}��*/۾�9�o_\�1���;���Y�f���w#�\�8��J�ZV��Z�.�V�RK�(�9��;$��"��B�7�������J[��� پ h���k?��������F��h(��v	ν��O�0�d?`��g��90��v���Aʾ��վ�   �   �֒�P���3����z�	�\��;�-V��\�@�������}�OK������(5
��mV�����F=���2��w��b��~:ԿN��s�h�7�4�P���e��lt���y�B�t�Јf�B5Q�z�7��g����CRӿ�c��a�u�pH0��,�z꡾_wQ���z��&��kj�꠆�q���T��� ���5�Q'X���v�𽇾�ʏ��   �   ��G�?�D���:���)�������v�Ƚ�^��k�m���@�c�<��o�n���l���f��l�������A�E����e������=��*��nH�4�d� �}�K��Eb���k����}��e��&H�`c*�jv��<�ٱ�]4���a?�����+��_`��A��}��j[��(��,�QY�g"�������V�d��&�&�)8�?�C��   �   �/�����	�������׽��H���5V��T"�Rl	�4���P[�������Vjp��b�����?�K��k��X��2� Q�Z�3��S�z�r�8��,;��쓓�#A���߆�ar���R���2�0*�����b���ǋ�bI�ڧ
��ŷ�!1j��M�K�����F������s��0#B����������ϽF$򽦴�����   �   k1�*& �$�۽nk��]���j�s��6���	�ԕ�Vw��	U�;o��_~��t��~��<��+O�ȏ��k���������6� �W�رw��͉��h���ז��c������Rw�f�V���5��y����O��G	���YL���������m���j���!@����xqż��꼰�"�h�`�M*������j�Խ8�������   �   �/�����	�������׽���G���5V�rT"��k	�^���O[�����a��:ip��a��<��]�K�+k��OW��	1�bP���3��S�>�r���`:�����Z@���ކ��_r���R���2��)����1b��&ǋ��I�A�
��ķ�0j�*M�h���¡F�*����/��#B����������ϽJ$򽨴�����   �   ��G�@�D���:���)��������F�Ƚ�^����m���@���<�uo�����	���f�3k������A�!���d����忪<���*��lH���d���}��I���`��3j����}��e�%H��a*�Nu�;俯ױ�D3��`?�a��k*��]`�6@��{��@
[���(���,��Y�B"�������V�i��(�&�+8�E�C��   �   �֒�P���3����z���\�n;�V�D\����I�����}��I�����:3
��jV�����:��L2���w��`���7ԿvL��q��7�T�P�Z�e�
it��y���t���f�p2Q�&�7�f�6���Oӿ�a��Q�u�0F0��)�W衾�tQ��}��w��#��#ij�Z������!��� ���5�S'X���v�򽇾�ʏ��   �   �@ھ��־�̾Zߺ�����][���!f��)6�d���׽�Q���ޤ�+8���h�,oC��z��Q+۾�6��[\�����"�������,u#�(�8�0J�bV�ԇZ�8�V��K���9�29$�` ��>�1���P���F[��>�ؾ�e��gh?���������D��L'���νn�3�0�Y?`��g��=0��v���Aʾ��վ�   �   �D�u��p������q��;�+���D����N�O��8=򽐓̽��ͽ׈���k/�D�����4���=�th~��#����˿W"�������[-�Z�6���:��7��k.��9 ����A���;�̿����z~��7=�3{�&ǻ��~�cn,�j*��¬ƽ��ĽI������^I��6��Rԥ��Nʾ��	�����+��   �   �6a��]���R�2�A��K+�(6����"����[�\��-%��[�VA����c����[�h��Ng�;����S��?������VͿ!�&���A�z�����ȁ��?����+E�\Ͽ�4��E���5�T����"P�f띾 )Z��������߽�I���S!�o�W��$���˻�?�쾀�#)�m�?�fVQ���\��   �   �[������̏��/��Jj�)�H�RT%��e���ɾv��c�\�>|$�h�����`��Z�8��@�����Na�� �*�˒]��������)¿�ڿ��ei�����4^�����ܿ�!ĿZ���NዿOa_�ٻ+�����G���x���y8�R�������,�I�!���Y�lI����ƾ����#���E���g� 炿zɎ�o����   �   .�ȿƿ����#˭�=��������[��l.�����ƾ�/����O�\i��y�n1�����NN��뎾�žL���,�.�X����_٘��$���^��DBſ��ȿ� ƿ����Dȭ�����r���[��i.�����ƾ:-��l�O�{g��x��1�8��uQN��
žy��؉,���X�����ۘ�i'���a��kEſ�   �   2���a��k��"ܿ�$ĿҴ��e㋿�d_���+����vJ���z��:|8�V�������+���!��Y��F����ƾ����#��E���g��䂿�Ǝ��~���X��$���ɏ�-���zj�C�H�Q%��b���ɾs��;�\��y$���������9�8��B�������d����*��]�����>���+¿�ڿ���l���   �   ������bA�h��H��Ͽ7������T����+S�s흾�+Z������*�߽�E���P!��W��!���ǻ�G��|��)�n�?�RQ�L�\��1a�_�]�z�R�}A��G+��2������p��\��*%��Y�,?�ȣ��L���[��i���i���r�S�8A�����[YͿ�#���C�R���   �   ��:��7��m.��; �f��ǚ��]�̿ფ��}~��9=��|�Aɻ���~��o,�@+��Ϋƽ�Ľ��齉��LZI��3��wХ�Jʾi�� �@��\(��@����������l���;�'���A����N����8�J�̽�ͽ����l/�T��������g�=��j~�3%����˿�$��b����]-�J�6��   �   ��Z�:�V��K���9��:$��!��@�Ҋ������H[���B�ؾ�f���i?�����Z���B���#���ν���0��9`�{d��0,���q���<ʾ��վ&;ھE�־o̾�ں�i����W���f��$6�T`�U�׽�M��Bܤ�17���h�-pC��{���,۾8�]]\�ہ������W�2��zv#���8��J�XV��   �   ��y�v�t�6�f��3Q�b�7�g���#Qӿ�b��
�u�tG0�z+�|顾�uQ�r~��w�����idj�Ɯ��*�����������5��!X���v�����SǏ��Ғ������/���z�+�\�j;��Q�vU�h��L����}��G��n���u3
��kV�[���X;��G2��w��a��9Կ0M��r�$�7���P���e��jt��   �   �a���j��L�}��e�&H��b*��u�
<俄ر��3��a?���R+��+^`��@�
|���[�ӧ(�9�,��Y�<�������P���@&���7��}C���G���D�I�:���)�H�������ȽbZ��ҕm���@��<�?�n�,���+��Cf��k��
����A������d�����*=�H�*��mH��d�}�FJ���   �   �����@��P߆��`r�n�R�l�2��)�s�b���ǋ�"I���
�Wŷ��0j��M�����i�F������J��OB�V��������Ͻ� 򽠲����Z-�����������B�׽��HE��A1V��P"�*i	�r��DN[�d���Z��_ip�b��d����K�Zk���W��b1�P���3�p�S���r�����:���   �   �
��Q��.�����zZr��&K���&�fL��ѿ�����c�3��о����7#�zG���:c�N��0���z?���B����l먽�mν��0m��)�yt�6������N���ӽ����t���O����s	����FVp��TȽ3'��b���zӾc��e�M��	�ӿ�s��A(�|cL�V]s��@��OO��,���   �   � ��" ��R����	����m��G��Y$��>�AοU?��y�_����B3;z��o�!����Hj�[H �.��,,��e��9���½�g��?����� ��>$��{!�̚�lr
�:��W�ǽ�[��c�q���8��X�*�,�FDw���Ƚ�z%��f���	о�k�b�����Lп�K�(z%���H���n��@��4˚�����   �   3���d���
���݁��`���=� ��/���%ſ�����U�D'�p�þ6{���vý�2���NI��M��g~�XA��7ٽ�����"�}:�)�M��Z��^�)�Z��dO�]�<��o%���
���߽�ѭ�.����RZ���U�����*�ɽc� ��l�ƾ���
W�-��A}ƿ�����Zb>�%a�qԁ�]���A���   �   ���c���M�����k��M���.����g�鿕9�������FD�W��@���:�j�ׅ�Z4ǽA#��0���丛�d�ƽ���!�%��L���q�/Ӊ��T���"���a��4����p��)Q���:u�4�O�\:)�d*�dyͽ.��ͤ���#���Nͽ?���&n�9ٶ�*����E��a��~!��ũ��B���.��MM��k��`��vF���   �    �v��:r��;d�4YO�t�6��C�����ѿ�!��s�s�K�.�P���C���LV�^��xAн������g��r��:F�P{������ ���;�Rᾘ!�������⾿�Ͼ�)���ě�\�m7J���ʜ��Ľ����S�ս1]�Q:Y� ޣ����/���t�������ѿ������D�5�VN��;c��q��   �   ��P��M��QB���1��������R��9���>���mR�{��}9Ѿ(���C	A��	
�%ὰg߽j��*� �a�[���.0����� ��t���$���-��"1��O.�%�%�Ͷ���-��Ļ�� ��{�e�C.���G|�%��8<�1C�`��XCҾoK�µR� 6��_㵿Q�ῒ�j��R�0��AA� oL��   �   ��,�x@*�t�!�T���s������ ���Pl��/�g���P᯾�[s��!-�!��N�����5���q�!����ѾN�}� �e<�T)U�^�h��u��&z��>v��j���V��8>�]a"����9Ծ'���u���7�U2�L����	��~.�|t��C�������\/�8�k��X������!I�l�����D!�֮)��   �   �y��h
����/@���ؿձ��{����w���>�����˾l#����M�Ƙ��o	�X��a5�s�X~����ݾ�y�4�5��i\��ހ��g��5t��-妿����f���\��n���3����^���7���-"�F(��߆u��%7��X�DZ
�|,�f�M�����Z˾��}�=��`v�/ᙿ�)��y׿X^�!���	��   �   �B޿��ڿ��п�G��w��8蒿�s���A����Wݾ�O���fg��\-�K�����8�,�MAf��\����۾[��r$@���p�+���훩�̾��}ϿNڿF޿L�ڿնп�J��1���꒿�s��A�0���ݾR���ig�z^-����ݛ��,��=f��Y����۾���
!@���p���������Ⱦ�'zϿ�Jڿ�   �   �����c���Y�����������^�.�7�e���G%����u� #7�zW�9Z
��-���M����?]˾��v�=�pdv�|㙿V,���׿�a�`#���	��{��j
�����C���ؿc����
����w�P�>����|�˾3%����M�y��ao	����^5�es�{��`�ݾw���5�|e\�8܀�7e��Bq��⦿�   �   �!z��9v��j�7�V��4>��]"�L��*5Ծ�#��u�6�7�V0�����+	�A�.��~t��E�� ���._/�a�k��Z������K������F!���)���,��B*�h�!�������񜾿���{Sl��/�Q���:㯾^s��"-�����K��u��U�4�,�q�����Ѿa��� ��`<��$U�r�h��~u��   �   �1��K.�U�%�N�����|侯�������D�e�Y?.����Py�.�彾<��2C�����EҾ0M�-�R��7��V嵿�������>�0��CA�TqL��P�<M��SB���1�,�����U⿉;���?���oR����h;ѾO���[
A��	
�h
�
d߽����*���a������+���������p���$�s�-��   �   ������6�⾜�Ͼ%�������U�W2J��(��Ľ�����ս�]� <Y�}ߣ�@��J�/�ȹt�9�����ѿ��������5�XN��=c�P�q���v�=r��=d� [O��6��D���*�ѿ�"��G�s���.����D���MV����R@н= �����:꽴n��5F��	{�����2���ޣ;FMᾡ��   �   �]��&����l���M��Y4u�ߪO��5)��&��sͽD��?����"���Nͽ���n(n��ڶ�-��<�E��b���"��W���C���.�0OM�zk��a���G��A���~���H���V�k�^�M���.�d����鿌:��y����GD���"���#�j����3ǽd!�����������ƽĖ���%��K�j�q��ω��P��x���   �   �^�(�Z�"`O��<�l%�m�
�2�߽ͭ�Ρ���MZ���U����g�ɽ� �n�ƾ̻��W��-��6~ƿ����Jc>�J&a�*Ձ�3���B�����e�����jށ���`�J�=��������ſM���QU��'��þ�6{����ýM1���JI�W�M��`~��<��@1ٽN���"��x:�[�M��Z��   �   ,<$�Gy!����^p
����5�ǽY��B�q���8�\V���,��Cw��Ƚ8{%�Lg��=
оvl��b�%����LпL��z%�$�H�p�n�GA���˚�|��?!��� ������/
���m�Z�G�Z$��>��ο�?����_�"��t3;���m�!������Fj�>F �J��w,��e��6��@½&d��=�7��V� ��   �   zt�:������N��/�ӽ��������O�r��t	�����Vp�'UȽC3'��b���zӾ��R�e�:M��/�ӿ�s��A(��cL�r]s��@��XO��2���
��K��.��}��`Zr��&K���&�PL�κѿk���ׁc��2�ډо���7#�)G��S:c��������4?���B����O먽�mν��(m��)��   �   /<$�Ky!����Zp
����'�ǽY���q�,�8��U��,��Bw��Ƚrz%��f��N	о�k��b�����Kп�K��y%�:�H�>�n��@���ʚ����C �����ھ��u	����m�z�G�\Y$�X>��~ο�>����_�x���2;�����!�����gEj��E ����6,��e��6��;½'d��=�<��Z� ��   �   �^�,�Z�&`O��<�l%�b�
�
�߽�̭�x����LZ�@�U��~��v�ɽ�� ��k�Zƾ����	W��,���|ƿ���t��a>�$a��Ӂ����A��K���c��!
��݁���`���=�h�����;ſ����U�x&�L�þj4{�~�ý!0��YII�l�M��_~�r<��01ٽJ���"��x:�a�M��Z��   �   �]��(����l���M��Q4u�ЪO��5)��&��sͽ������� ��5Lͽ���8%n� ض�b����E�a��� �����B���.�`LM� k��_��ZE��틎�@���C����k���M���.�������[8��ȇ��5ED�K��º���j���1ǽ������곛�.�ƽ���x�%��K�n�q��ω��P��~���   �   ������9�⾚�Ͼ%�������U�,2J���L�� Ľj�����ս_[�38Y��ܣ����A�/���t�����+�ѿ���b����5�NTN�l9c���q���v�L8r��9d�HWO�؇6�<B�����ѿ ��6�s���.����+B���IV�)��8=нF���N��꽂n��5F��	{�����7����;NMᾪ��   �   �1��K.�V�%�N�����|侠���y�����e��>.����w佪��
:��.C����-AҾ�I���R��4���ᵿ/��H������0��?A��lL�N�P��M��OB���1����0���P��7��=��kR�����6ѾC���PA�
���a߽����*�R�a������+���������p�Ó$�w�-��   �   �!z��9v��j�6�V��4>��]"�D��5Ծ�#���u�{�7�//����p	�|.��xt�SA��v����Z/�h�k�	W�������F�����R!���)�h�,�V>*�n�!�~�|�����Y�������Ml���/������ޯ��Ws��-�M��H��b����4�͠q�n���Ѿ^��� ��`<��$U�x�h��~u��   �   �����c���Y�����������^�'�7�Y����%���u�"7��U��W
��)��M�����W˾z���=�2]v�ߙ�'����ֿ[����	��w��f
�����<���ؿ���+����w���>����[�˾� ����M�����l	���]5��s��z��J�ݾ w���5�~e\�:܀�:e��Eq��⦿�   �   �B޿��ڿ��п�G��v��5蒿�s���A����'ݾMO���eg�K[-�������,��9f�=W���۾C���@���p�\���h����ž��vϿGڿ?޿O�ڿ'�п�D������咿�s�L�A���@ݾ�L���ag�6Y-�#�������,��<f��Y��n�۾���!@���p���������Ⱦ�+zϿ�Jڿ�   �   �y��h
����.@���ؿұ��x��v�w���>���|�˾#��{�M�����l	��
�[5��s��w��,�ݾNt�:�5�la\��ـ��b��bn��ߦ��󩿴`���V������R
��@�^���7�s��q��!��r}u�7�#T�.W
�w*��M������Y˾v�x�=��`v�0ᙿ�)��{׿[^�!���	��   �   ��,�x@*�t�!�T���r�俾���
 ���Pl���/�5����௾�Zs��-����VF��Z��[�4��q������Ѿ���� �]<�` U���h��yu��z��4v��j���V��0>�kZ"�S��^0Ծ���Qu���7��,�����N	�}.�{t�DC��i����\/�5�k��X������#I�l�����F!�خ)��   �   ��P��M��QB���1��������R��9���>��vmR�i��<9Ѿ�����A��
����^߽M���*�"�a�J���Z'��Q����m���$�v�-��1��G.�v�%������bw��������^�e��:.����ks����%:��/C����CҾbK���R� 6��`㵿S�῔�j��T�0��AA�oL��   �    �v��:r��;d�4YO�v�6��C�����ѿ�!��n�s�>�.�"��C���KV�Ș��<н1�������꽦j�u0F�H{�Ѓ������ʞ;�G᾽������X�Ͼj ��Ƽ���N��,J�����`�ýƔ����ս�[�N9Y��ݣ�ʞ��/���t�����ѿ������D�5�VN��;c��q��   �   ���c���M�����k��M���.����g�鿓9�������FD�H��
�����j�����0ǽf���~������Ǫƽ*���%���K�?�q�̉�M��o��cY������h��	J���-u�D�O�71)��"��mͽ&��������Kͽ��)&n�ٶ�����E��a���!��ȩ��B���.��MM��k��`��wF���   �   2���d���
���݁� �`���=� ��-���&ſ�����U�<'�O�þ�5{��Dýl/��6FI�|�M�,Y~�
8���+ٽ����{"�Xt:���M���Y��^�!�Z�R[O���<�h%���
�2�߽ȭ������FZ�>�U�z}����ɽ�� �Tl��ƾ����
W�-��D}ƿ�����Zb>�%a�qԁ�]���A���   �   � ��# ��R����	����m��G��Y$��>�AοU?��w�_����23;`���!�ؗ��Ej�)D ����
,��e�(4��$½�`��;������ ��9$��v!�B��6n
������ǽ&V��C�q�\�8��R���,�(Aw���Ƚcz%��f���	о�k�b�����Lп�K�(z%���H���n��@��3˚�����   �   �
�������{�����eU���\���3�d����]����t��;)�����h��0� �ҽVA{��%�hj�
�#�_OX� b����߽Ρ�ַ����(�AV���������A�� R���+_��*�4F��,�DV����ֽY�2�1퐾�⾍�*��`v�_|��}K�,����4���\������5��Ֆ�������   �   a���|S��.����������bX�&�0�*��;dݿ���ׯp�>s&�ݾ�V��*�.��ҽ�Z���3��#�dn@���|��u����ҽ�������>�"���,��F0�%-�y�#��L��� ��8ֽ���������dG��i*���:����I�ֽm1�~ώ�;�޾��'�_Pr�������޿��� �1���X���6˗�,����N���   �   b���K�������3���t���L�~R(�zQ��Dӿ%���� e�mc�ޛҾ/e��s�)�*YԽ/	���v_��0d�H�������뽔���R/�U�H��]�[*j���n�D�j�r1^�xXJ�.1�L��3�� n������Ak��pf�
���$7ؽ�+�����LԾzx��f�����ANԿ,��<�(��VM��t��,��n���/���   �   R���:���$��T����^�.<��h��k���Xÿ���*S�:����¾��|���"���ؽ@!��zѕ��Y��h?ؽ�m�Z�2�d�[��-��F��ڪ��  ���[��rd��d��;<���F��HG^�5�����1ܽz��hK��⎥�E ܽ%�$�����þI���T�G5��mĿ;������<��G^�����َ�����   �   +܆�����x�bY`�څD�0�'�r>�R��N宿�Ⴟp<�;�[����f�E!����p�½��ν������$�Y�U��J��>[����¾A:ݾ/>�����_�2 �o6��޾&<ľ2̦�e����cX��'�$� ��8ҽ�ƽ�%�����h�|������ڵ<��7���-������(��F'��C���_��Qw�Y؃��   �   r�a���]���Q�|H?��%)�8D�� ÿ�w����a��"���྄�����O����,���������8��Qs����ekǾi �+��G�!��0�l�:��3>��;���1�@�"� �������ɾ=�����u��:�Z��P���O�� Q�/Q�b���Ᾰm"��*b��q��;�¿��־�Be(�@d>�d�P��S]��   �   ��9���6�ҽ-�������
���	�˿�棿~}�͉<�oK��򼾒Â��G:�$��*�8�v!C�f&��oc�����m+�<�,�C�J��e��z� Ń��.�����#�z��Pf���K��.�";��i��Ů��9���D����rF	�	�{!;�� ���4��%R�Ta<��}�tn���!˿��V:����H-�
y6��   �   x��(�2�H�n��Ƭǿ�����ℿ��L�����ھḚ���\��\(�����G�.=C�n˂�$�����2z�܄C�-�l��t�����6����岿����C�������霿�M��X�n���D�Q~�tJ�w*��Đ��4UD�@������(�]�n���}�ھ��.L��R��&��3�ƿq�FR�2������   �   ���/B��0߿�Ϳ����E��8=����O����U0��𫾤2x�J:����Zp�;�9�Hzw�mS��V2�+��w�N�<|���R�������̿�N޿B��Y���E꿃4߿M�Ϳe��
H��R?���O����#4���5x�:����xo��9�Xvw�pP��.�T��КN��y��P��������̿�J޿����   �   ]���@��ߜ���朿K���n���D�i{�F�>'������qRD�������(��]������ھS��\L��T���(���ƿYt�T�2����$z��*�&�����}�ǿ����x䄿��L�	���ھͺ����\��](�L���E��9C��Ȃ�������w� �C���l�Vr���������ⲿ�   �   �+�������z��Kf�T�K��.�$8��d�a®��6����D�����E	�S�#;�4"��7���S��c<�
}��p��+$˿��<����~-�h{6�X�9���6���-����`��ٷ��a�˿�裿�}��<�M������Ă��H:���N)�v5�xC��#���_�����H(�u�,��J��e��z�@��   �   !/>�K;���1���"�Ҹ�A����ɾ����=�u��:����*���N���Q��0Q��c����ᾘo"�`-b��s��U�¿���^��g(�df>���P�fV]�$�a�&�]��Q��J?��')��E�a ��!ÿ^y����a�"���ð����O����\���������8��Ks�����fǾ������t�!���0��:��   �   \\��. �f0�z޾I7ľ
Ȧ������^X��'�"� ��4ҽpƽC%彆���h���������<�!9��i/�����*�XH'���C��_�Tw��ك��݆����.x�l[`���D�~�'�z?���࿙殿�₿�<�,�����@�f��!���὚�½4�νL���"�$���U�RG���V����¾�4ݾ8�B����   �   NW��`���_��t8��lC���A^�G5�1��,ܽJ ���H��|���C ܽ�$��
�g�þ`��ET�Q6���Ŀ�������<��I^����ێ�"������V;���%��U��f�^�L<��i�Dm���Yÿؚ��MS������¾��|��"�ōؽF��6Ε�HU��+9ؽ�i�g�2�y�[�p*��-B�����������   �   &�n���j�[,^��SJ�1�Ŀ�T��qi��x����<k�Cmf�O���b7ؽ��+������MԾSy��f�M���EOԿ����(��WM�>�t�m-��o���0��c���L������y4���t�t�L�S(��Q�3Eӿ�����!e��c�~�Ҿ�e����)��XԽ���}r_��*d�J��� ���j������N/���H��]��$j��   �   OD0��"-��#��J��� �v5ֽ�򩽀󁽪aG�lg*�C�:�c����ֽ�1��ώ���޾�'�Qr����O�޿@��|�1���X�{���˗�����CO�������S���������J����X�j�0�\���dݿH��� �p�ms&�Lݾ�V��&�.���ҽ�Y����3��}#�Yj@���|��r��/�ҽt������Ƈ"���,��   �   (�CV����������A��CR���+_�J�*��F���,��V���ֽ��2�c퐾b�⾽�*��`v��|���K�B��ڡ4���\������5��▮������
������u{�����UU���\�~�3�L�����\��[�t��;)���ྮh���~0���ҽ�@{���%�j���#�	OX��@��|�߽ġ�ʷ�����   �   QD0��"-��#��J��� �m5ֽ��d�SaG��f*�g�:������ֽ1�Lώ���޾\�'�Pr�m���j�޿�����1�|�X�����ʗ�����3N��տ���R������2��������X���0�����cݿ�����p��r&�TݾJV��R�.���ҽY����3��}#�j@���|��r��,�ҽt������ˇ"���,��   �   -�n���j�a,^��SJ�	1����0��:i��$���;k��kf����X5ؽ2�+�v����KԾ�w�$�f������MԿ�����(��UM�Ȼt��+��1m���.��a���J�������2����t���L��Q(��P��Cӿ_ߞ��e��b���ҾJd���)��VԽ����p_��)d����Ӡ��T������N/���H��]��$j��   �   SW��`���_��u8��iC���A^�05����+ܽ�����G������pܽ��$�!���þu���T�z4��a Ŀ�������<�ZF^�����؎���������8��a#��S��H�^��	<��g�Mj��1Wÿ����	S�����¾E�|���"� �ؽ���͕��T���8ؽ�i�X�2�v�[�r*��2B�����������   �   a\��. �l0�z޾F7ľȦ��g^X�l'��� �43ҽDƽ�!����կh��������d�<��6���,������'��E'�x�C�Ԍ_�Ow��փ��چ�)��6x�2W`��D���'�D=�e���㮿�����
<���|���B�f���6�ὂ�½�ν������$���U�KG���V����¾�4ݾ8�L����   �   &/>�N;���1���"�ϸ�:����ɾz�����u���:�ޒ�����ZJ���N�,Q�d`�����l"��(b�ep��c�¿ӄ�t���c(�>b>��P�2Q]���a���]�H�Q�ZF?�
$)��B����ÿBv��,�a��"�4��~�����O�%�������:����8��Ks�����fǾ������w�!���0��:��   �   �+�������z��Kf�Q�K��.�8��d�>®��6����D�b���C	�s��;����(2��{P�_<��}��l��C˿C��8���&�,��v6���9�B�6���-����������z�˿�䣿�z}�8�<��I�𼾁���CD:�%�|'�S4��C�U#��s_�����F(�u�,��J��e��z�C��   �   _���@��ᜪ��朿K����n���D�_{��E�'��6���TQD�$��}���(��]����Lھ���HL�Q���#���ƿ�m濂P�D������u��&�2�n����ǿ
���������L�x	��ھ8�����\��Y(�����C��8C��Ȃ�h�����w� �C���l�Xr���������ⲿ�   �   ���2B��0߿�Ϳ~���E��6=����O���'0�𫾥1x��:����l���9�rw��M��&*쾳��p�N��w���M����[�̿nG޿ӻ����q>�b-߿��Ϳx
���B���:����O����+���-x�u
:�9��m�a�9�buw�*P���-�K��ΚN��y��P��������̿�J޿����   �   x��(�2�H�m��ìǿ����ℿ��L���u�ھw���A�\��Z(�����B�6C�fƂ�/��:��+t�^}C�8�l��o�������x߲���Z=�������㜿oH��S�n���D�Bx�A�#������ND�`�Y}���(��]����E�ھ��(L��R��&��4�ƿq�GR�4������   �   ��9���6�ҽ-�������	����˿�棿~}���<�WK���Â��E:�g��&�)2�9C�� ���[��̟�M%���,���J�9e�^z������(������z��Ff���K�%.��4��_�]����3����D�ׇ�bB	�M��;� ��>4��R�Ma<��}�tn���!˿��X:����J-�y6��   �   t�a���]���Q�|H?��%)�8D�� ÿ�w����a�z"�������e�O�������j�����~8�0Fs�(	���aǾ���z����!���0�ͫ:��*>��	;�`�1���"�d��Y���ɾ�����u�,�:�ˏ������H���N��-Q��a����ᾩm"��*b��q��=�¿��ؾ�Be(�Bd>�d�P��S]��   �   +܆�����x�bY`�څD�2�'�r>�Q��M宿�Ⴟc<�$�	����f������K�½�ν������$��U��C���R����¾*/ݾ2�����"Y��+ �K*��t޾@2ľ�æ�X����XX��'�g� ��.ҽpƽ� �'���h�,������ҵ<��7���-������(��F'� �C��_��Qw�Z؃��   �   R���:���$��T���^�0<��h��k��Xÿ���#S�+��Z�¾�|�r�"��ؽ ��eʕ�rP��3ؽ�e���2���[�"'��p>������H����R���[���[���4���?���;^�<5���O%ܽ����FD�������ܽ��$� ���þ<���T�G5��pĿ>������<��G^�����َ�����   �   b���K�������3���t���L�|R(�zQ��Dӿ%���� e�dc���Ҿ�d����)��VԽ����m_��$d�f���%���|��^���J/���H��]��j���n���j�8'^�
OJ��1������&d�� ���{5k�Igf������4ؽY�+�Ǽ���LԾtx��f�����DNԿ.��>�(��VM��t��,��n���/���   �   `���|S��-����������`X�&�0�*��;dݿ���կp�<s&�ݾ�V��˹.���ҽ�X����3�*{#��f@�f�|�p����ҽ����q��f�"�x�,��A0� -��#�?H��� ��1ֽ�墳����F]G��c*��:����)�ֽ1�`ώ�,�޾��'�^Pr�������޿����1���X���5˗�,����N���   �   ���Z���ȷ����M��`�e�
�:����a�\ܯ��7~��/�`l�����O7���ڽ�����-��V��t+���a�v���������}6��� ���,!�`�#��Ī��������ؖ���c���-�����/�DC���jܽ�78�͊��J1꾏j0��~�wR����鿮���d;��Uf����r:��rԷ��\���   �   ��������������������a���7��2�3��A���z���,�e��*̒�Zt5��4۽�Ɇ�3<�^+���H����������ڽ���p3��*(�Wn2�H	6��2�4�(�Ԯ����<�۽�8��ꄽ�_K�b|-��>����l�ܽ�V6�\���d�|-�`�z�����K�J��>88�Bb�`,���������������   �   ����/Z������\����� �U�P�.��d�<-ۿ/�n��$���ھ����0B0���ܽ�̒��i��m�tǑ��޽�I����\���5��P�R�d�FMr��w���r��Re��P��n6�,��E���6��X���dp��ok����D޽^1�d��yp۾F%�.�n�I��^�ۿ���%/���U�+���Y��=ا�AN���   �   ��}��H���_��F/h�ڋC��=!����B�ʿ)&��J*[���ʾ�$��z�(�x��d���5қ�� ��*�ཥ����9�Jd�J��
ř�����.1��K����W���娾�"��Iw���$e��x:�٘�J�~l��0��]�����ҍ)�Y�����ʾ����[��e��I�ʿ���fV!�.�C��h��D��(��z���   �   �x��$k��-�����i��VL�T�-�@D�A���O���ʇ��3C���+��Xho�.� ��a꽮=ʽ<�ֽ���%+�0^��w��8����@ʾ�徫U��̩������5���&澫�ʾw=�����_���+�~�(�׽rd˽k��rx!��p�>����B�@xC�;5n����迈;�ض-�JL���i�掁��O���   �   ��k��Xg��6Z�ګF��V/�g����� ʿk����[j��/(�,N��H��}VW��V��c������./��x?���|��#���$Ͼ8q���Q�	(�}�7�m�A��2E�A�A��7�2d(�b���+���Ͼ�����}�T9@���������`��p��M�W�ύ����P(��pj�J�����ɿ`^���/��/�PKF���Y�"g��   �   �KA�&�=�6,4��H%���������ҿ�����S���qC��@��þ�h����@��/�*��i���NJ��	��y���i����O�3�Y�R�:�m�Z���,���_��@ǈ��pgn��S��4��#���܌���p��>�J�J7��^�H��A�u���:�þ�C��aC��;������Z�ҿN���Ԗ��$���3��=��   �   x���w�
�y��￑~ο=���G����T�i����� ����d�O.�}��&�"��.J�z����ɸ�������!�%K�2v�ɏ�����Q���u������U���9���5[��� ���v�ΩK�&�!�"����3��4ᇾ|�J���"�B%�p*.��d�����⾎[���S�BZ���e��*	ο�￶.�����R��   �   >`���x������Կ�N��௢��Ɔ�{W�<>%�X{��Nױ��?��"@�� �� �?@����Z���f��&�$���V��y���N���޼�C8Կq�濓F�/d���|�o��P�Կ�Q��z����Ȇ��
W��@%�L��ڱ��A���#@�_� �"� ���?����@�����3�$�ԔV��w���K���ۼ��4Կ��濰B��   �   �����������BX��K����v�	�K�"�!�����`0���އ���J�b�"�3%��+.��d���x��
^�>�S�Y\��-h��(οN￠0����"U�����y���z�3��a�ο����1����T�������"�� �d�	.����L�"�|+J�唇��Ÿ�����d�!�!K�S-v�NƏ����@N��[r���   �   ~��mĈ�^~bn���R��4�� ������&n����J�5��]�����A������þ�E��dC��=��䄩��ҿq������0�$�*�3���=�hNA���=�x.4��J%�������;ӿ����tU���sC�:B�&�þ�i����@��/�������mJJ����t���d꾴��a�3��{R�*�m�����S����   �   �-E���A���7�P`(����%��B�Ͼѯ���y}�$5@���������_����!�W�~�������Q(��sj������ɿa��01��/��MF�l�Y��$g���k��[g�(9Z� �F��X/��h�����ʿ�����]j�1(�SP�9J���WW��V��a�������+�t?���|�����Ͼ k��N�(�.�7��A��   �   ��7�����l澟�ʾ)9��x���z�^���+��z� �׽*b˽���.y!�bp�䔵�6D�zC�{�o������<�d�-�6L��i�D���Q��z���l��|���&�i�HXL���-�TE����QQ���ˇ�35C���7,���io�o� �W`꽼:ʽo�ֽ���{ +�6^��s�������;ʾE��PO��v���   �   ����gS��ᨾ����s���e�t:����O�,h��\��췩��⽘�)�6����ʾ@��L�[��f����ʿh��|W!���C��h�F��R)�����o�����UI���`���0h�
�C��>!�z��W�ʿ�&��x+[����ʾ$%����(����V����Λ�������~��n�9��Cd��	�����S����,���   �   �v�!�r��Me��P�Wj6��
��?��2�����8_p�Flk�'��~޽1����q۾&%�j�n��I��k�ۿģ��&/��U�����Z��?٧�SO��ȱ��3[�����d]�������U���.�^e��-ۿ��n�{�$�^�ھ󕌾\B0�s�ܽ*˒�U�h���m�VÑ��ٽ������X��5��P���d��Gr��   �   �6�?�2���(���������۽�5���焽T\K��y-���>�Z��ǫܽ:W6��\���e�}-�#�z�z���ML濮���88��b��,��|������}������f�����������;	���a���7��2���w���z��,����?̒�Tt5�T4۽;Ɇ��<�*+�e�H�謃�����L�ڽ���1��'(��k2��   �   �,!�b�,��˪���� ���ؖ���c��-�z��6�/��C��Xkܽ488�����1꾿j0�V�~��R��������d;��Uf�����:��~Է�]�����Z���ȷ����=��B�e���:�����`�8ܯ��7~���/�l�����ZO7�h�ڽ������-�@V��t+�j�a�P����������p6�������   �   �6�D�2���(���������۽�5���焽�[K�fy-�Ն>������ܽ]V6��[���d�L|-��z����`K����78�� b�,������
���b�������K��������������a�.�7�`2��������z�S�,���得˒�ys5�B3۽�Ȇ��<��+�&�H�Ѭ������L�ڽ���1��'(��k2��   �   �v�)�r��Me��P�Vj6�z
��?���1��P��*^p��jk����h޽n1�����o۾� %�c�n�vH����ۿ���,%/��U�����X��Pק�<M������Y������[��J���U�z�.�>d�5,ۿa��n��$�q�ھ�����@0�^�ܽ�ɒ���h���m�Ñ��ٽ������X��5��P� �d��Gr��   �   ����lS���ᨾ����s���e�t:�Ҕ���ng��2�������T�)�t���U�ʾD��}�[�e��3�ʿ���~U!���C�^h��C���&�� ��������F���^���-h�x�C��<!�����ʿ%���([��}��ʾf#����(���ང���͛���J��_��^�9��Cd��	�����X����,���   �   ��;������p澟�ʾ%9��n���W�^�D�+��z���׽�_˽���zv!�3p������A��vC�4퇿�l�����t:�x�-��L���i�����#N��w���i��ϸ����i��TL���-�C�E��aN���ɇ��1C���)��meo��� ��\꽒8ʽ�ֽ"��> +�^��s�������;ʾL��XO��|���   �   �-E���A���7�R`(����%��9�Ͼ����|y}��4@� ��:���$\������W�������VN(��nj�������ɿ\��&.�/�.IF�X�Y�Dg���k�Vg�4Z���F��T/�~e�����ʿ�����Xj��-(�JK��F��=SW��S�,^��&���;+��s?�z�|����zϾk��N�(�3�7��A��   �   ���oĈ�`�bn���R��4�� ��������m����J��3��[����)A�������þ�A��_C�f:�������ҿg������$���3���=�TIA���=��)4��F%������(�ҿi���)R���nC��>��þwf��]�@��,��������IJ����U���d꾰��`�3��{R�.�m�����V����   �   �����������DX��L����v��K��!�j���,0���އ�|�J���"�c"�m'.�i�d�E�����KY���S�XX��Gc��]ο���,�����P�@��~u���.w���ￓ{ο����/���{T���Ϧ�Y����d��.�,����"�]*J������Ÿ�����^�!�!K�R-v�PƏ����BN��^r���   �   C`���x������Կ�N��௢��Ɔ�uW�.>%�*{��ױ�T?��u @�a� �"� �e�?����:������y�$�T�V�|u��0I���ؼ�w1Կ���>�V\���t��濁�ԿyK��#���4Ć��W�<;%��v���ӱ�N=��@�{� ��� �A�?�o���������(�$�ДV��w���K���ۼ��4Կ��濳B��   �   z���w�
�y��ￒ~ο<���E����T�W��P�⾰��|�d�.����"�'J�C���Y¸�*���]!�NK��(v��Ï�����K��o�� �������ŏ��;U�������v��K���!�o���,���ۇ�&�J���"��!�>(.���d�C�����[���S�AZ���e��+	ο�￸.�����R��   �   �KA�(�=�4,4��H%���������ҿ�����S���qC��@���þh����@��,����V��FJ���������_꾚����3�swR�D�m�����������������쁿r]n��R��4����������j����J�61�SZ�w��AA�䋇���þ�C��aC��;������\�ҿQ���Ԗ��$���3��=��   �   ��k��Xg��6Z�ܫF��V/�g������ʿj����[j�o/(��M�|H��	UW�yT�]������m(�go?���|�����ϾHe���J�6(���7�z�A�n)E�M�A���7�Y\(�h�����*�Ͼ����@s}�0@����<���KZ��/����W�_���ؔ��O(��pj�J�����ɿb^���/��/�RKF���Y�"g��   �   �x��%k��.�����i��VL�V�-�@D�A���O���ʇ��3C����*��Bgo�v� �r\�N6ʽ��ֽ	���+�|^�;p��p����6ʾ���I��.��;���������j�ʾ�4����b�^���+�w���׽
]˽N�뽼v!�op�쒵��B�8xC�:6n����迊;�ض-�JL���i�玁��O���   �   ��}��H���_��F/h�؋C��=!����A�ʿ(&��D*[��~�aʾ?$��?�(����~���ʛ����R��~����9�>d�G��%������(������N��.ݨ����@p���e��n:����f⽞b�����
���⽖�)�����Q�ʾ����[��e��J�ʿ���hV!�0�C��h��D��(��{���   �   ����/Z������\����� �U�N�.��d�=-ۿ0�n��$���ھb���gA0���ܽ!ɒ�;�h�y�m�L����Խ�����)U�ֽ5�	P���d�"Br�p�v��}r�9He�$�P��e6���9���,��&���Wp�!fk�x���޽�1�(��Vp۾?%�-�n�I��a�ۿ���%/���U�,���Y��<ا�BN���   �   ��������������������a���7��2�3��@��z���,�U��̒��s5��3۽TȆ��<�4+���H���������޿ڽ����.��%(�i2��6���2�/�(�/��x���۽|2��儽�WK�Bv-�x�>����@�ܽQV6��[���d�{|-�^�z�����K�J��@88�Bb�a,���������������   �   r����7��8����������0g���;��;�-g꿎���`2�!y0����
����6��Uٽ��x)����&�2]�ߖ��@�������8����������$���Y����&��!�������b[�'%�����A'�����>ؽ<6����-l�o0�ͺ~��I���꿠��j�;�L�f��{���ף�U���76���   �   �r��E����z��xF��ů��j�b�2�8�>��ʸ�ŭ��{�v�-�b$��ڒ���4�1�ٽǄ��7���&��D��������>�ؽ���J�`2'��Y1���4�P61�u�&�������dؽU��������B���$�0�5��΃�^�ؽ(^4��v������3-�r�z�%{��*[�����r8�${b�1����9��x�������   �   =������>�������b}���nV���/����ܿҊ����n��	%��)۾Ǔ��5�/���ڽ�ʐ���d�i�i��ʏ�v���F�[���5�lO��/d��wq�J�u��Mq���c��O�Ƥ4�$��@���
ӎ���g���b�ُ���ٽ�$/��8���ھ�$��tn�cN����ۿ���<o/�MV�u������|���$���   �   ����ڼ���͖�Xφ���h��&D�j�!�p9��=˿ӡ��0�[����m?ʾF
��i1(�߽�����Ι��>�� ߽�)��'9���c�����ۀ�������<���䱾�N���k������Xc�v�8�L��� ޽AE��^㘽�����"޽�'�<���F�ɾ����[��w���˿d#���!��$D���h��������ˡ��   �   �
���������&j�<�L��7.�r���F�JƵ��!����C�9��4����n�� �����KȽ��Խ����*�5�]��w��@ҫ��|ʾ���������X�;��S������ʾ\n������]�� *�ׂ�6�ӽ�pǽV��K��_|n���3�|sC��
������>����N.���L�ܹj�N1������   �   ��l�0�g�̣Z�r�F��/� �������hʿ\C��1�j�g(��h龋 ����V�or��r��\��Zf�[�>��c|�DB��}ϾC ��/���r(��
8�HB�^gE�V�A���7��5(��k��}��,Ͼ�ۣ���{�5c>�l��h8��5������MV���:�GR(���j��E��C{ʿX(�����/��7G���Z�\h��   �   &�A�TY>��l4��n%���J���,ӿ6ީ�u����C�G�͝þ����?��)���d����I��솾�*��2����U)4�Q/S�Z�n��������R��Gꈿb����Vn�+�R���3�#��6d��ɳ������<I���Ī�\���?�"�����þOF���C�[���� ���fӿM���9���%�V�4�,y>��   �   �c����2����￤�ο�ȫ�ѝ��+T�Xt��d�?���)~c���,�Z���!��`I�ma��<ڸ�Hb���!�:�K��w��R��뛢��䰿�����	��7ܹ�µ���a�����%�v��sK��!�9���\���2+��(I��t!�y��1�,�wc������⾉��VOT�7Ɖ������ο�𿒿��\�Z���   �   u���>��B��ԿkQ�����O���n�V��%�K��Q���H���>��A��J�$�>�R��ڀ���[���O%�>W����q�آ���տ�\���i�������@�ԿjT������}�����V�l%�A���S��gL���>�B��I���>�=}��}��QW���L%�L:W��򆿰����6տ�X�����   �   E���ع������^������v�pK��!����� ����(��FI�is!�h��z�,��yc����������RT�Pȉ�����οb �~��_����f����4�ގ�c��t�ο9˫�����* T��v�h�B���n�c���,����*�!�"]I��^���ָ�D]����!�3�K��w�8P��ޘ��Y᰿%��   �   +O��q爿�����Qn���R���3���J_�Ƴ�����9I��}�Щ������?�����<�þ9H���C�������4iӿt����:���%���4��{>���A��[>��n4��p%����L��E/ӿ/੿�v��ޙC��H���þH����?��)�������x�I��醾�&����꾲�b%4��*S�D�n���������   �   �bE���A��7�2(�3h��w��WϾ�ף���{�_>����5�����~��OV�b��<�9T(�J�j��G��m}ʿ�*�������/�B:G�H�Z�2 h���l���g�P�Z���F���/�v��S����jʿ�D��y�j��h(�k��!��ԩV��r��p��R ��#c���>�Y]|�4>��xϾ#�������n(��8���A��   �   �����L��B���ʾj��S��']�{�)����ӽ�nǽ��	��9~n�=﴾z�TuC���������@�T��jP.�z�L�:�j��2�����0��\��@��^�j��L��8.�����H鿥ǵ��"��*�C�:�%6��,�n�> �a���HȽ��Խo��*�6�]��s���ͫ�vwʾ��征���Z���   �   J8��C౾�J���g��J���%Rc���8�h����ݽ�@������@����"޽ج'������ɾ��,�[��x��
˿@$�̰!�6&D�x�h������.͡�����7���$ϖ�]І�|�h�&(D�T�!�$:��>˿����b�[�t��m@ʾ�
���1(�P߽샦�g˙��9��~߽�%�}"9���c��톾���z|��T����   �   ��u�Hq���c���N���4�] ��:�
��Rώ�m�g���b�K؏���ٽ�%/�69��<�ھͿ$��un�2O����ۿ���p/�4NV��u���������+%��P�����-���I����}��|oV�(�/����vܿ^���r�n�
%�D*۾���a�/��ڽ.ɐ�M�d�3�i��Ə�*��&@�~���5�gO�a*d�rq��   �   J�4��31���&�;������ؽy��b����B�N�$���5��΃���ؽ�^4�w��n��S4-�6�z��{���[�^��zs8��{b�����(:���x��;���:s������c{���F�����ַb�~�8�t����Dŭ�{���-��$�ے���4�ĖٽDƄ���7�`�&��D�阁����z�ؽ��@H��/'�W1��   �   ���%���Y����2&��!������c[�l'%�$���A'�{���>ؽJ<6�R���ul龟0�	�~��I��꿸����;�l�f�|��أ�a���=6��r����7��,����������g���;��;�g�j���&2��x0���龷
����6�{Uٽ��)������&��1]������������8�������   �   N�4��31���&�;������ؽn��K���þB���$���5��̓���ؽ�]4�bv��i�徒3-�(�z��z���Z�Ɵ��r8��zb�嗈�A9���w�����r������Wz���E��X�����b���8����*�濍ĭ�� {��-��#�fڒ��4���ٽ�ń���7���&���D�Ԙ��w��x�ؽ��CH��/'�W1��   �   ��u�
Hq���c���N���4�X �g:�
��ώ�g�g���b��֏���ٽ$/��7��L�ھ^�$��sn��M��պۿ`���n/�8LV�|t����������#��+������<��������|��~mV���/�j���ܿ���j�n��%�T(۾ג����/�
�ڽ�ǐ���d�%�i�>Ə��
��@�w���5�"gO�g*d�rq��   �   P8��H౾�J���g��J���Rc���8�G��<�ݽ<@��bߘ�q����޽��'�W����ɾ��^�[��v���˿�"�̮!��#D��h��������jʡ����t����̖�;Ά��h��%D�T�!��8�i<˿������[�x���=ʾ
	��j/(�h߽���:ʙ��8��߽�%�h"9���c��톾����|��Z����   �   �����L��G���ʾ
j��K��]�>�)�P���ӽylǽp��W��zn�촾 ��qC��	������=� ��|M.���L���j��/����	��cߊ�����|j�N�L�6.�4���D鿯ĵ�^ ��ОC��7��2���n�� ����FȽ��Խ���*��]��s���ͫ�wwʾ��徉���`���   �   �bE���A���7�2(�4h��w��PϾ�ף���{��^>�����2��b�����KV���7龘P(�T�j�{D��Zyʿ�%�����8�/��5G�,�Z��h�Ƚl�^�g�4�Z�.�F���/�j��S���yfʿ�A����j�e(�f�m��Q�V��o�m������cb�J�>�]|�!>���wϾ�������n(��8���A��   �   .O��t爿�����Qn���R���3���:_��ų�����F8I�X|��������?�M���(�þ�D���C�̄������dӿd���N7���%��4��v>���A��V>�Dj4��l%� ��F��/*ӿܩ�Gs��۔C�E��þ���<�?��&���������I�]醾�&����꾮�`%4��*S�F�n���������   �   H���ع������^������v�pK��!�����͉���(��*I��q!����*�,�esc�<����|�D��RLT�Kĉ�'��'�ο�𿺽��Z�0���a�P���/�����￥�οQƫ������T��q�&a�z����yc�L�,���\�!� \I�|^��Uָ�']����!�-�K��w�8P������[᰿)��   �   z���A��D��ԿlQ�����O���k�V��%�!���P���G�A�>�?��F�J�>��x��z��0S��J%��6W�����좿�����տ2U�%�����\���o�ԿKN��a���������V��%��
���M���C���>�.>�7G�%�>�7|�s}��&W���L%�H:W��򆿯����8տ�X�����   �   �c����2����￥�ο�ȫ�Н��%T�It��d�յ���|c���,������!�"YI�1\���Ҹ��X����!�g�K�Aw��M��핢�)ް��ﹿ���tչ�M����[��K��ӟv�lK���!����� ����%���I��o!�����,��uc�;�����x��NOT�5Ɖ������ο�𿔿��\�\���   �   *�A�VY>��l4��n%���J���,ӿ4ީ�u����C�G�y�þs����?�'����J���I��憾�"����꾔��!4�^&S�U�n�L�����KL���䈿�����Ln�>�R���3�����Y�����ɛ�� 4I��y��������?�����N�þ9F��C�X���� ���fӿO���9���%�X�4�.y>��   �   ��l�2�g�̣Z�r�F��/��������hʿ[C��+�j��f(��h� ��"�V�+p��k�������_��>�GW|�S:��'sϾA���0��k(�n8�M�A�>^E�\�A�5�7�.(��d��q��B�ξ�ӣ�H�{��Y>�����.��|�����PLV�A��9�7R(���j��E��C{ʿZ(�����/��7G���Z�^h��   �   �
���������(j�>�L��7.�r���F�IƵ��!����C�9��4����n�C �x��~DȽp�Խ���b�*�s�]�Cp��mɫ�hrʾ,��E����������vF��k�從ʾ�e�����]���)��{���ӽ�iǽ7�罓��B{n�F��rsC��
��	����>����N.���L�޹j�O1������   �   ����ۼ���͖�Xφ���h��&D�l�!�p9��=˿ӡ��,�[����4?ʾ�	��,0(�b߽����nǙ��4��߽�!��9���c�ꆾ���8x�������3���۱�6F���c�������Kc�\�8�"����ݽj;��ܘ�_����޽ڪ'�ػ���ɾԛ���[��w���˿d#���!��$D���h��������ˡ��   �   >������?�������c}���nV���/����ܿҊ����n�z	%�z)۾����l�/�F�ڽǐ�<�d�ƪi��� ���9�Ν�?5�ObO�$%d��lq���u�nBq�2�c���N��4����3�G���ʎ�6�g�s�b��Տ�&�ٽ,$/�E8���ھ�$��tn�aN����ۿ���<o/�MV�u������}���$���   �   �r��E����z��wF��ů��j�b�2�8�>��ʸ�ŭ��{�r�-�T$��ڒ���4��ٽYń�P�7�p�&�'�D������ ��
�ؽ���E�T-'��T1���4�11�n�&�������0ؽH��������B���$���5�(̓�8�ؽ�]4�uv������3-�p�z�%{��)[�����r8�&{b�1����9��x�������   �   ���/������.��YC�� ,_��!6�r��+��?l��cdw���*�⾑���)/��ͽ=o���� � ��xjK�y���	����ٽ�?�����=O�B.�������T����(׽���ޱ���7E��W��e���O��h��ʽ��,�H2��"F�%�)���u�;k���t�2&�`A5��K^����U���̰������   �   �;��4���i�����~��[�>3���� �����8Ks��'�}P޾�j��9E-�N�ͽ�v�0�&��9��r3��{p������>ͽb<���2�~���O)�%�,���(������Gq��5ʽ<o���!j�8&-�*��̒ ��p�UʽK#+�@����ܾu�&���q�ᵧ���޿r��jG2�&EZ��3��Ɍ��h۬������   �   ﴱ��s�����i���hw�>CO�A*����P�տl����cg������ӾPJ���(��DϽ�����R���W�i��$6��t����RF-�$�F���Z�ُg�
�k��g���Y�0cE���+�P���}�C̭��ł�R<Q�|vL�T΃���˽^ &�"��8ҾU���'f��џ���Կ�U�j�)�\�N��3w����Ȝ��8����   �   ����g������������`���=� �������3ſ����(�T�K���þ�{��� ��8ӽ�)���ʏ�����9Iӽ>e
��K1���Z��Ɓ�
쓾�;���W��;\��Z���ה������ʀ���X�!F/�mz�׸Ͻ�b��e���x���нg���y���������S��j��@�Ŀ7��Ƣ�Զ=���`�IƁ����*���   �   �r��+c��z���a���E�,�(��/�>�-4��{ԃ�&7=��������le�6���Uܽ�����;ɽD2��	#���T��4�������bþG�ݾ��& �6Q���������ܾ�¾�Y��������R��%!�<���Fƽ����wٽ�K�y�c�ȭ��v���<�D���=����!��C�p�(��JF���b���z�����   �   �Dd�X�_���R�$@�P�)�r���8�6ĿD��c��"����!��}�M�A����S��v���6���r�TP���OȾ���r����"�R�1���;���>�>;��c1�$"�������i�ƾ�����fp�L 5���
����3뽭�`}L�/�����ྺi"�?�b��J��WĿ!��ZT��~*���@���S�*`��   �   $�;��8�,|.�� ��O��F���x̿_c���8~�2�<��Q��X��t���r7�[������<1A�����ݶ����\A��c.���L��2g��|�����oֆ��j��P<{�`f��`K��K-�JL��Kᾣv���À�ʭ?�U�M�����6�DX�� ��M�S=��~��Ф��0Ϳ�V������� ��&/��w8��   �   ������`��|F�9���ǿ$������k�L���X�پHl����Y���$��s����@�Z��+�����D��$_E��|o��������╫�R���2��x�������� ��T3���n��2D�����.��e��T�?��c�2�� �$��Y�ㅙ��Sھx3��mM������㦿�ȿG�
����C��   �   :�\���߿��Ϳ����:���!��vbO�� ���R��
xt�8
6��|����e6�)(u�d窾���{��TiP�Ԃ��������ο�࿝�����_�x�߿�Ϳ�!��Q=���#���eO�D#�����T��q{t�6�)}���\c6�4$u�a䪾��쾜���eP��т�&�������ο:������   �   4/��2������������0��n�/D�*��2��l+���b����?�Db���`�$���Y�*����Vھ�5��pM�����e榿k�ȿsJ����� �:E������X��FH�c�{�ǿW&��� ��R�L�.��\ ھ=n���Y�m�$�vs�����@�����'�� ����:[E�xo�����������N���   �   �ӆ��g��7{��f�]\K�/H-�HI�G�s��Z���1�?��R�[��J�6��Y���"���N��=�S�~��Ҥ�a3Ϳ�Y��z�� ��(/�Bz8���;�@8�X~.�� ��Q��I��{̿Le���;~�u�<�/S�
[������#s7�4����"��4-A�ʹ��񲭾��+>��_.�*�L��-g�J|�ӣ���   �   d�>��9;��_1�F "�e�������ƾ:����`p�8�4��
���� 2�7�"L�̈́���ྚk"���b�qL��'YĿ����U���*��@��S��`��Gd���_�N�R�&@��)����&;�Ŀ�E��Fc���"�"�D#����M�,A�'��O��s�K�6���r�bL���JȾ�y�������"��1�Z�;��   �   �M����z���ܾ�¾yU��{����R�b!!�*���:ƽ���xwٽ�L�B�c�^�������<�z�������t#�E���(��LF�ʚb�l�z�랅�Ct���d���z���a�r�E���(��0��?�5��}Ճ��8=���ܞ���me�t��ZTܽ ���07ɽ�+���#���T��0��,����]þ��ݾ���� ��   �   �W�����������
��<ǀ��X�_A/��v�
�Ͻ�^���������н#����y������S��k����Ŀ�8��У�&�=���`�Uǁ����Z+�����������������f�`�̿=�������4ſ����R�T���zþ�{�� ��7ӽ�'��:Ǐ�ĭ���Bӽ-a
��F1���Z�xÁ� 蓾D7��DS���   �   |�k�\�f���Y�{^E���+�����w㽈ǭ�����7Q�$sL��̓���˽!&����XҾ-���(f��ҟ���ԿVV�4�)�d�N�5w���������>��������t��Հ��(���iw�DO��A*�b��	�տ�����dg�5��9�Ӿ�J���(�fDϽ0��1�R�z�W�\���0��#�����A-�O�F���Z�^�g��   �   �},��(�=��� �^m���1ʽml��Bj��"-����h� ��p�rUʽ�#+������ܾ��&���q�[���}�޿����G2��EZ�64��G����۬� ¹�!<���������|���Q~��x[��3����] �/����Ks�1�'��P޾	k��4E-���ͽ`�v���&�`6��n3��vp�l����:ͽ08���0����M)��   �   ?.�������f���)׽��� ����7E�,X�@f��dP���h�;	ʽ��,�z2��hF�U�)��u�`k���t�J&�|A5�L^����e���̰��������)������.��IC�� ,_��!6�Z����l��*dw�u�*���b����/���ͽ�<o������ ����jK�M��������ٽ�?��v��6O��   �   �},�"�(�B��� �]m���1ʽcl��j��"-�H���� �3p�jTʽ�"+�����ܾF�&���q�������޿B��$G2��DZ��3��k����ڬ����	;��������������}��n[��3�&��u�|���zJs�t�'��O޾bj��\D-���ͽ��v���&��5�Jn3��vp�d����:ͽ,8���0����M)��   �   ��k�f�f���Y��^E���+�����w�]ǭ�����6Q��qL�R̃���˽s&����wҾ˰�	'f�1џ��Կ@U�λ)���N��2w�_��盡�>���糱��r���~�����Tgw�0BO�>@*�D��M�տ�����bg�Χ�W�ӾdI��@(�XBϽ�����R�v�W����0�������A-�P�F���Z�g�g��   �   �W�����������
��>ǀ��X�TA/��v���Ͻ^������N���н���a�y�x����V�S��i��5�Ŀ�5������=�~�`�UŁ�g����(��Q������E�������*�`�L�=������u2ſ�󓿔�T�&���þ��{��� �5ӽ�%��Ə����nBӽa
�hF1���Z�vÁ�!蓾I7��JS���   �   �M�!�������ܾ�¾xU��v����R�*!!�d����ƽ���#tٽJ�8�c�L���j�J�<�G��������B��(�4IF�z�b�Z�z����]q���a��|z�P�a���E���(�n.�<⿚2��CӃ�R5=����ě���ie�����Pܽ�����5ɽ�*��C#���T��0��&����]þ��ݾ���� ��   �   i�>��9;��_1�K "�g������ƾ*����`p���4�f�
�8��_.�f��zL�~���6�h"��b�LI��3UĿӿ��R�}*���@�2�S��`�Bd���_�x�R��!@�|�)����G6�ĿgB��qc�'�"�����L�M�N>�u��]M�s���6�;�r�LL���JȾ�y�������"� �1�^�;��   �   �ӆ��g��7{��f�a\K�0H-�GI�G��r��'����?��Q���)��6�{V�����TK�=��~��Τ�o.ͿT����� ��$/��u8���;��8��y.�� �6N��C��v̿=a��.5~���<��O�V��\����n7�P������t,A�����Ͳ�����$>��_.�)�L��-g�O|�գ���   �   7/��4������������0��n�/D�%����<+���b��r�?��`�f��.�$�]�Y�����TPھC1��jM��~���ᦿ��ȿ�C�@���� A�қ����^���D�����ǿ�!������.�L������پ�i����Y�:�$��p�4�z�@�}��R'�������3[E�xo�����������N���   �   =�\���߿��Ϳ����:���!��tbO�� �����Q��wt��6�<z����_6��u�n᪾������5bP��ς������^�ο�����l{�QX�Q�߿q�Ϳ���#8��Q���^O�������N��st�]6�Xy�����a6�/#u�䪾[�쾎���eP��т�%�������ο=������   �   ������b��~F�;���ǿ$������d�L�����پ�k��y�Y��$��p�����@�B��$�����&���WE��so�^�7�������xK���+��������������.��tn�0+D���B'��`��.�?��^�����$���Y�v���NSھf3��mM������㦿~�ȿG�
����C��   �   &�;��8�,|.�� ��O��F���x̿^c���8~�(�<��Q��X��詁�Jp7������Ƀ��(A�ﶁ�-���&��!;�\.��}L��(g�
|�����І�8e���1{��f��WK�bD-�F��A��n��H���w�?�2O�7����6��W������L�E=��~��Ф��0Ϳ�V������� ��&/��w8��   �   �Dd�Z�_���R�$@�R�)�r���8�5ĿD��
c��"��ᾒ!���M��>�j��.J�Zp���6���r��H���EȾ�s�����8�"��1��;���>�O5;��[1�o"������ҽƾA����Zp�V�4�I�
�M�齈,�x��{L�����J�ྩi"�7�b��J��WĿ��ZT��~*���@���S�,`��   �   �r��,c��z���a���E�,�(��/�>�-4��zԃ�7=����[����ke�����Pܽ�����1ɽ�$��#�H�T�|-�������Xþ�ݾ��� ��J�����\��ݼܾ�¾#Q����'�R��!�����Mƽ����rٽEJ�c�c�t���^���<�C���>����!��C�p�(��JF���b���z������   �   ����h������������`���=� �������3ſ����"�T�>��JþU�{�m� �5ӽv$��VÏ�֨���<ӽ?]
��A1���Z����T䓾3���N��DS������{������À��X�Y</��r�T�ϽdY��A���L��:н2��]�y�i�����z�S��j��@�Ŀ7��Ƣ�Զ=���`�JƁ����*���   �   ��s�����j���hw�@CO�A*����Q�տk����cg����w�ӾJ���(��BϽ"��8�R�@�W�f
��,���潆���=-���F��Z���g��k���f�x�Y��YE�:�+����q�D­�����0Q�?mL��ʃ�N�˽�&����ҾL���'f��џ���Կ�U�j�)�\�N��3w����ǜ��8����   �   �;��4���i�����~��[�<3���� �����8Ks���'�kP޾�j���D-�(�ͽ��v���&�z3��j3�/rp������7ͽK4��u.�����J)��z,���(�Ǭ�}��>i��.ʽWi��j�~-�6��J� ��p��Sʽ�"+�$���ܾs�&���q�൧���޿t��jG2�&EZ��3��Ɍ��i۬������   �   '������޷�����R�w�J�O�Ȇ*��	�&�տ����tg�"n�)]Ҿ����� ��*���O�Q��Paμ`c�� �-���q������Ľv��:�������
��T�����F��ƿ�����6�f�fV"�L^ༀA��x���mC�t�����������Ͼ���#e��C���Կ����K)�jbN���v��͏����*����   �   �ޭ�����������r���K�J�'������ҿ	 ��u�c������ξ�������`����V��$�l���~�^�P�􈎽����F�1v����������D��\�i��6ݽ�C���׈�V3E��m��߼�����J�`첽�J�À��/̾��aa������п����&�d�J�fr�ό����©��   �   ]p��퓞�~��LR����d�7A�R�� � �!�ȿ{���SX������ľ|\z�<
�����|�l�R�4�V?9���j�j=��N�н������E�6���I��^U��Y��tT���G�Jz4��%�J��ʽ1"��,�^�2�-�0)���`��h��ܤ�hv��a¾�j��tV�zT���0ǿ���������@���d��[��z��(����   �   Tv��������2o���P�`E1�X�8O��������P�F����NC����h����;��G��7}��`���c���/��~�"���I�-�o����rW��yʞ������9���J������o�l�k_F�ZH����L��0n��K�q�M���`�����Tge�NE�����\E�����1���~���J:1���P��o��@���T���   �   �{�*�u�`-g���Q�Pk8�������;ԿB����v�<�0�e�����ˍS������ƽn8��yδ���-]��AD�cGz��������`fξ����Q�?S����ྀ�̾-���n���P;v���@�[����۽`@�����ִ�������P��u���m񾔡/���u�+����Կ6��`K��(9�:�R�H(h�̜v��   �   $�S�­O��3D��C3�,�����?������l����S����r/Ѿ�ό�<+=�@O��׽��ս����Q�'�]`��Ӓ��>��p���-���	&���.�@�1�|r.��%�j��M����Nͷ�����k\�o�$�}��rѽ �ҽ�B��&;�΋�75о� ���S��u��/�����ra	�P��ld4�=E��NP��   �   �Q/��,�L-#�n���Y���������kZm�%0�p�������Ro��&(��$�����V	��1���o�(:���!Ӿ�`�"�
?�E$X�9�k��x�0|��]w�tj�n�V��X=��!����о�5���l�@�.�E�R�˪ �b�&�%En��B������FF0�w�m�ja��p����h��T����v$�"�,��   �   �3���(���/��hٿ����Q���Ex���>�f4��4ʾ�ʍ�u.H����n�8��0�0�>Zp�VQ��C߾Y�a_8�(`�!��:Γ�Ԡ�� ��y�����������U���끿��]���6�?���ݾ����Xn��F/��Z�ܒ�#��H�_�d�ʾW���?���y��m������*ۿ[���z�d��   �   ɸ�Y�ܿq�ѿo����I���Ⓙ��r��#A�����ھv���`��q&�e�	��
�y	'��	b��b��5:ܾR���B���t�.��_���S@¿��ҿ�cݿd���ܿ��ѿ�����L���䒿��r�'A����|�ھ�x��9�`��s&���	��
�S'�b�`��56ܾ� �A�B���t��+��z���=¿x�ҿS`ݿ�   �   O���ဨ��񟿠����聿��]�N�6�����ݾ����!
n�D/�?Y�ƒ�L	�@H�������ʾ����?���y�Np��R���:-ۿ����|�`� 6��� ��!3��kٿ[��T��@Ix���>�k6��7ʾ�̍��0H����(n�����0��Up��M��{>߾c��[8���_����l˓�Ѡ������   �   �|�VXw�2oj��V��T=��!�)���о�2���l���.�
C�QP�� ���&�Hn�E��)����H0�� n�lc�������k翢V�r���$�T�,��S/��,�L/#�8��[����U�������F]m�F0�r���
����To��'(��$�,��zT	�Q}1�H�o�y6���Ӿ���"��?��X�2�k��x��   �   �1�fn.��%���.��~��ȷ�����bf\���$��w��bѽ��ҽ C��(;��ϋ��7о�"��S�Gw��(�����b	� ��bf4�<?E�8QP���S��O��5D��E3������m�þ���m���S�z��n1Ѿ�Ќ�a,=�ZO�׽/�ս�����'��`��ϒ��9��ک�������&���.��   �   M���^��K�̾���������4v�`~@�o����۽�<��o��\���F��>�P�nw���o�>�/�$�u������ԿR���L�r*9�6�R��*h�L�v���{�� v��/g�ڧQ��l8�F��~���=Կ�����v���0�6�����S�����ƽ�5��ʴ�J��X�{<D��@z�ﯙ�񌵾aξ�ᾶK��   �   c}���5��G����� �l�ZF��C�������0j���q�����R���H��he��F����H^E�����p��N�����|;1�0�P���o�B���U���w���������3o��P�pF1�,��P����h���k�F����7D����h�.��:��%E���0}�b\���]���'��µ"���I���o�g���vS��Lƞ��   �   wY�koT���G��u4��!��� �v�ʽ���Y�^�:�-�)�%�`��h��{��]iv��b¾~k��uV�7U���1ǿȏ�������@���d�D\��S	�����Lq��ϔ��H���R����d��7A����� �эȿ�{���TX�$��%�ľ]z�c
������l�:�4��99�/�j��8��R�нd�������6���I��YU��   �   6����KZ��f��2ݽ�@��Ո�*/E��j�p�߼<�����J��첽K��̀�Z0̾��Rba�o�����п\�� �&���J�r��ό����+é�Y߭����9��r����r�T�K���'�����ҿ> ����c�ֺ���ξ�������V`��(�V��"�t�����~�P�����4���N��s�Q��4���   �   ��
��T�����T��ƿ�����t�f��V"��^�B��D��vnC�ӛ��������F�ϾD���#e��C���Կ����K)��bN���v�Ώ�#���0���'����ӷ�����8�w�0�O���*��	���տ����ftg��m��\Ҿ������ �x*����O�P���`μ�b����-�}�q������ĽY��#������   �   :����PZ��f��2ݽ|@��Ո��.E�zj�x�߼����f�J��벽TJ�̀�p/̾��]aa�ʹ����п���r�&�
�J��r��Ό����1©�Wޭ����P�����^�r�f�K�֯'�6��	�ҿ�����c�%����ξ^���0��J_����V��!�<���L�F�P��(���F� t�T��5���   �   �Y�uoT���G��u4��!��� �b�ʽ�����^�P�-��)���`�	g����gv��`¾3j�%tV��S��?0ǿč��6���@���d��Z�����G���oo�����������Q��~�d�"6A������ �-�ȿCz���RX����\�ľ�Zz������X�l���4��89�{�j�L8��*�нS�������6���I��YU��   �   g}���5��G�����$�l�ZF��C�����n���i����q�M�������:��ee�5D��"���[E���5���}�8��B91�Z�P�X�o��?��bS��!u��{�����<0o�8�P�&D1�^��M����������F�����A����h�
�88��`C��x.}��[��]���'����"���I���o�f���wS��Qƞ��   �   M���h��S�̾���������4v�G~@�;��H�۽X;��u��:������w�P��t���k�4�/��u�񱤿/Կ<��,J�H'9�`�R�&h�Z�v��{���u�+g���Q��i8����^�$:Կ���c�v���0���(����S�f��b�ƽ�3���ȴ�j⽨X�L<D�s@z�毙�쌵�aξ�᾽K��   �   �1�ln.��%���1�����ȷ�����*f\�1�$�~v��<
ѽ��ҽV@�w$;��̋�3оX���S�Rt��o�����$`	�����b4��:E�zLP���S�b�O�p1D��A3�|��P���������j����S�'���,Ѿ�͌�6(=��L�t�ֽ��ս`�����'�Z`��ϒ��9��Ω�������	&���.��   �   �|�[Xw�8oj��V��T=��!�'���оl2����l�5�.��A��L�U� ���&��An��@������D0���m��_��4���f�jS����x$���,��O/�V,�B+#�����W�(�快}�����5Wm��
0�̡��f����No��#(� "����QS	��|1���o�S6���Ӿ�����"��?��X�5�k��x��   �   Q���倨��񟿣����聿��]�M�6�|���ݾn����	n�C/��W�2��Y�R�G�&�Z�ʾD��V�?�Q�y��k������'ۿ�����x�p��1���J��Q,���dٿ���O���Ax���>�2�I1ʾ"ȍ��*H�����k�Ό��0��Tp��M��X>߾W��[8���_����l˓�Ѡ������   �   ͸�_�ܿu�ѿs����I���Ⓙ��r��#A�����ھ�u���`�wp&��	� 
�'��b�E]��p2ܾ���B���t�)������	:¿ �ҿ�\ݿ3��бܿ�ѿF���G�������r�f A�f����ھ�r��_�`�In&�1�	�z 
��'�b��_��6ܾ� �8�B���t��+��z��� =¿{�ҿW`ݿ�   �    4���*���/��hٿ����Q���Ex���>�X4��4ʾIʍ�1-H���xk����l�0��Pp��J��):߾��8X8���_�,
���ȓ� Π�l���+����}���ܰ��"恿v�]���6����ݾ����n�@/��U�����W H���"�ʾC���?���y��m������*ۿ\���z�f��   �   �Q/��,�N-#�p���Y���������gZm�0�I��������Qo�%(�E"�۽�JQ	�9y1���o��2��4Ӿ��P�"��?�X�H�k�ix��|�%Sw�;jj�T{V��P=�!�0�șо�.��M�l�j�.��?�XJ�(� ���&�	Dn�qB������8F0�n�m�ga��n����h��T����x$�$�,��   �   $�S�ƭO��3D��C3�,�����A������l����S���8/Ѿ;ό��)=�&M�|�ֽ��ս;�����'�`�U̒��5��y�㾪�����+&�y�.���1�Pj.��%�J������ �Sķ�뤐�`\��$��p���ѽȬҽf@��%;��͋��4о� ���S��u��,�����ra	�N��ld4�=E��NP��   �   �{�,�u�b-g���Q�Rk8�
������;ԿC����v�3�0�<����ɌS�����ƽ�1���Ĵ��⽻T�)7D��9z�����S����[ξf�ᾷE��F������̾�|��v���.v��x@����۽�6�������������P��u��jm񾇡/�ڝu�)����Կ4��bK��(9�:�R�J(h�Μv��   �   Tv��������2o���P�`E1�Z�;O��������L�F����C��2�h��
�68��B��O)}��W���W��~ ��6�"���I�F�o��􈾑O��1�4y���1�� C��t�����l�nTF�+?� y���
��$e����q�d�������r��fe�E��ؙ��\E�����0���~���H:1���P��o��@���T���   �   ]p��쓞�}��MR����d�7A�T�� � �#�ȿ{���SX����j�ľ\z��	�@����l�~�4��39���j��3����н������N�6��I�TU�TY�[jT���G�hq4���o� ���ʽ���2�^���-�x)�+�`��f��!���gv�la¾�j��tV�yT���0ǿ���������@���d��[��z��(����   �   �ޭ�����������r���K�J�'������ҿ
 ��t�c������ξ��������_��f�V�� ������P�\���������q������ŷ�t��W��d�/ݽ=��.҈�@*E��f���߼\�����J�J벽FJ�%̀��/̾��aa������п����&�d�J�fr�ό����©��   �   L��'���{����~���\�t�:�^}�j���/¿������P�K`��r��˝l����Q���*&&�����ь� ����1�b�E�/���7ʧ��ƽ��ݽ�L콲��+�wٽ�5�����/�z�@�3�c�|Ȍ�ؒM�����������4��Մf�\׸�s)�pN�ʏ�|��g���/��v9���[�b�}�;���ﰗ��   �   ���@c��2���d�x��vX�|7����}���
�� ���HM�C���C����h�
O�������,���μ�ܱ����U'�j&m�
����½�P��_��rG�/�	��!�8��P@޽�s������5[��� 徼0鋼����]�֓���?c�Tȵ�&�
��J��z��v��{����|k6���W�R�x�J���ci���   �   �D��9	���%����j���L��I.�R�� 鿑絿'��"C�����b^����S���δ@�~b�Ъ��B?������V���v彜6�B� �`�1��o<�Ӥ?��+;��v/�ܛ��;���ܽ������v�B1,��������X(.��T�������X�����@����@������]�������.�-���L�Лj�uL���*���   �   *����z�dqk��LU��m;�W �~~��s׿x����?z���2�D���/����^N�a ���Re���O�	t��Y����ڽ��ZY2�(�T���s�j腾�x���я�ɹ�������o�wP��t-���	�"�н����la���=���S��Z������ΥI�y]�����6M1��[x�ӛ��X�ֿ</�xK ���;�"�U��)l�~.{��   �   Z�_���Z��N�vM<�\�&�(#�����z���V��2Z^�����پSo��h�:����l���s���Aj����½���S-�Hl^�o���U���Ÿ��aʾ�zվ�ؾ��Ծ��Ⱦ�o��ͤ���G����X���'�;������Lې�J���H��f`뽟#7��o����׾8���J]�?锿7K��� �Α�HQ'��R=���O�,�[��   �   �b>�"�:���0��"����/��j�οAY�����h�>���^��l^z���&��l��k��0`��U�ݽx^���F�����螦��&̾���Q���G�M�������"'�}�tR�9�ȾZf�����fA����Z�ս�;�����k�S�#���w��й���h�>�!���^����Ͽ����F���1#���1��P;��   �   n��r����� ������sп�a��������U�n%�PV�����S�DE��s�٬н���a�T�l���� �����no��,���B���T��_��Vc�c�^��S���@�� *��\���幾�-���JP��\���� �˽+"ݽ�v��iR�I5��B��i�*�V�������)ҿ:���
	���xH��   �   ��7���i��сݿM	ſiM���A��<�_�jr+����Tz���{�� 0�l�1��TS���X�FU��~��Ⱦ�D��&�mJ���l�����#�������tT��l�������f���j� �G���#���@Fžie����Q�������	�Y��/��|�'��IY��*�,�4pa����;����ǿބ߿Ɍ�v���   �   F�˿Z/ȿ�������՚�"���k�Z��w-� ���Mþ_ދ�GF��D�����2�5���G�s��'ž����U/�4]����	���0���m��c�ȿ��˿�2ȿ���⍮�Tؚ�N���
�Z�wz-�[��%Qþ�����IF�yF�|��P1�F�O�G����v#žV���R/�N]�H��c���--���j���ȿ�   �   �Q��Gi�����d��Vj�Z�G���#��}�uBž�b����Q�>�����	�Z�d�/�}|��)��^]���,��sa�?��������ǿ�߿9��&z��_����������ݿſ�O���C��t�_��t+�Q���|��C�{��"0��f��FP���U� U��{���Ⱦ*B�? &�nJ��l�l���b��������   �   �Qc���^��S���@���)��Y���Ṿ�*��FP�lY�2��Z�˽�"ݽ�w�lR�d7�� E�l��V�\���)���z,ҿ="���	����hJ�b��X��������u��/vпd��-⊿I�U�\'�
Y�ѭ����S�1F�Ysὔ�нF��?�p�T�ݏ����I��(l�,���B��T�Q�_��   �   ���ά��#�J��L�h�Ⱦdb��T��PaA�����ս�8���ﱽ�l�Ȯ#�F�w��ҹ������>�����-����ϿL���� �t3#���1��R;��d>�&�:�^�0�*"�2�����j�ο�Z��L���R�>��	�+���`z���&��l�<j���\����ݽ�Z���F�O݂������!̾�����bD�QI��   �   �ؾ0�ԾZ�Ⱦ�j������bD����X�=�'��3��v����א�T�������a�!%7��p����׾����L]��ꔿ�L�������R'��T=���O�B�[�~�_��[�܎N�O<���&�D$����u|��X���[^�!����پVp��q�:�`��d�������<f���½���N-�f^�����Q�������\ʾ7uվ�   �   Ώ����8~����o�]qP��o-���	���н�����da��=�
�S��Z��
���1�I��^�����N1�j]x�����Íֿ0��L ���;���U��+l�n0{�+����z�sk�NU�o;��W �>��t׿g���3Az�� 3��������g_N�Va �r���e���O��t�XT����ڽ���5T2�2�T���s��䅾�t���   �   �?�';�Dr/�ח�m8���ܽ������v��*,�`���D{��'.��T��6����X����������@�g����^��-��h����-���L��j�)M���+���E���	��W&����j�l�L�PJ.�ش���2赿����C�w������b^����῞�t�@��^�x���;?�}���PQ��vp��2�� ���1�Qk<��   �   �	�j����<޽rp������E0[���߾��䋼�����]�L֓�h�c��ȵ���
���J�f{����������k6�N�W��x������i�����c��������x�dwX�V|7������.��0��IM�l��D����h�O�T���\�,�ȼμ`ױ����hQ'� !m����Z�½�L�x[��5E��   �   ���(�wٽ6�����`�z�z�3��c�,Ɍ��M�����
��r���t��(�f��׸��)��N�.ʏ��������,/��v9���[�x�}�D�������L��"���s����~���\�^�:�H}�B���/¿������P�$`��r��{�l�w�������%&����0ь�H����1��E����ʧ��ƽ��ݽ~L��   �   �	�o����<޽vp������50[����޾�䋼8���X\�fՓ����c�ȵ���
���J��z��7��(��h��0k6�P�W�ʏx�����i��2���b��ɣ����x�\vX��{7�f�����d
�����+HM����*C����h�HN�a����,��μ4ֱ���(Q'�� m����P�½�L�v[��8E��   �   �?�';�Nr/�ߗ�n8���ܽ����^�v�n*,�����px���$.�S�������X�U������8�@�G���.]��X��D����-���L�j��K��*��$D��t���$��L�j���L��H.�����}鿮浿w��C�D�����}`^�J������@�]�l��>;?�>���(Q��Sp��2�� ���1�Tk<��   �   Ώ����>~����o�`qP��o-���	�r�нC����ca��=��S�?X��B���M�I�{\��Q��7L1�GZx�횦�3�ֿ�.��J ���;���U�J(l��,{�)����z��ok�
KU��l;��U ��}�4r׿N����=z�y�2�M�������k\N�b_ �� ���e���O�[t��S��|�ڽ���T2�$�T���s��䅾�t���   �   ��ؾ8�Ծc�Ⱦk������cD����X�%�'��3��ƛ���֐��������]뽬!7�Kn���׾���I]� 蔿�I�������O'�BQ=�ƊO�$�[�:�_���Z��N��K<��&��!�ۿ�Ly���U��X^�T����پ�m����:����R��������d��2�½ĕ��N-��e^�����Q�������\ʾ=uվ�   �   ���Ҭ��#�N��L�h�Ⱦ_b��8��aA����U�ս�6��~챽�g��#���w��ι������>�ࡀ�ƶ���ϿX������0#���1��N;��`>��:���0���!�H�����7�οnW������*�>�������Zz���&��g��f���Z����ݽ&Z�=�F�3݂������!̾��� ��cD�TI��   �   �Qc���^��S���@���)��Y����๾�*���EP��X�.��(�˽�ݽ,t�ofR�63��#?��g���V�ޘ��㐮�j'ҿf��V		�L���F�|�������v�����"qп�_���ފ���U�2#��Rᾗ�����S�RB�8n�2�н� ���T��܏�|��5�� l�,���B��T�S�_��   �   �Q��Ji�����!d��Zj�\�G���#��}�aBžyb��l�Q�J�������|V���/��|�N$���U����,��la����������ƿˁ߿p��s�����|����~ݿqſ�J���?����_��o+�v���6w��J�{�?0�l�x��M���T�QU�Z{���ȾB�6 &�fJ��l�k���a��� ����   �   I�˿^/ȿ�������՚�#���m�Z��w-����Mþ ދ�(FF��C�Y��%,�J���G�]�� ž���O/���\����}��X*���g����ȿ��˿,ȿg��.���5Ӛ�ك����Z�kt-��~�Jþ�ۋ��BF��A�£��,���Y�G����D#žG���R/�D]�E��a���,-���j���ȿ�   �   ��:���n��ՁݿO	ſjM���A��<�_�fr+����!z��4�{��0���h���J���R���T��x����Ǿ�?��%��
J���l�𦅿����*����N��pf��U����a���j�e�G�M�#��z�B>žo_���Q�{�������W���/��|��&��!Y���,�,pa����8����ǿ݄߿ʌ�v���   �   p��t�����"������sп�a��������U�f%�(VΆ�����S��C��nὨ�н`��}����T��ُ�n����i�m,���B�u�T���_��Lc���^��S���@�<�)��V�%쾭ܹ�a'���@P�[U����֊˽Dݽu�whR��4���A��i� �V�����뒮��)ҿ:���
	���xH��   �   �b>�$�:���0��"����1��l�οBY�����e�>���&���]z�G�&��h�f���W����ݽ�V�r�F�ڂ������̾��ʇ��@��E����� �	�G�j�Ⱦ;^������[A������ս\3���걽�g��#���w�|й���]�>����[����Ͽ����D���1#���1��P;��   �   \�_���Z��N�xM<�\�&�(#����{���V��0Z^�ݾ���پo��u�:�����������wa���½4���I-�`^���kM��
���mWʾ�oվ��ؾ��Ծ*�Ⱦ4f��c����@����X�8�'��+��
����Ґ� ������l]뽤"7�Co����׾,���J]�=锿6K��� �Α�FQ'��R=���O�.�[��   �   *����z�fqk��LU��m;�W �~~��s׿y����?z���2�,��������]N�
` �� ��*
e��O�t��N����ڽ���6O2�j�T�|�s�DᅾBq��6ʏ�Q����z���o�~kP��j-�p�	���нϜ��x[a�h�=�n�S��W�������I�D]�����-M1��[x�ћ��W�ֿ</�xK ���;�"�U��)l�|.{��   �   �D��:	���%����j���L��I.�T��鿑絿'�� C��������a^����>���̮@�FZ����4?�,�L��Dj�K/�� ���1��f<�m�?�m";��m/�Ǔ��4�0�ܽp�����v��#,�4����p���".��R�����:�X�����6����@������]�������.�-���L�Лj�uL���*���   �   ���?c��3���d�x��vX�|7����}���
�� ���HM�@���C��k�h��N�����̎,�̸μ,ұ�(��VM'�m��
����½�H�YW��C���	�;������8޽�l�������*[�����׾��ދ�P���[�Փ���	c�Dȵ�"�
��J��z��u��z����|k6���W�R�x�J���di���   �   ����l���p��SY�"�>���"�"����ڿ,��d~�>�5�
I���V��<�I����J�{�|�＠�T������N�ԝ���m�2�P�:[��I㠽�^��R���<ŽD����Y���P��=w�J�7���� 5{� ����}�*��Pe��JX]�6:ܽ��A�?���F�ϓ2�Άz��!��y�ؿBn���!���=���X�:�o�����   �   ���<�z��ik��IU�h;�K �$l�UD׿�`����y��h2�]��l���K�F������{� �������<M��ѓ���|6��Az��M��Ę��i>ҽ1�p��k�ܽ�!̽鲽Jv���a�t��h���h.�p�����lw��F^�N�ٽJ�>��M���)�n�/��tv�2{���0տ&`��]���:�R�T�FYk��z��   �   �q��l��(^���I���1�|��M6��WͿ�@���Tm�l\)�t{羬w���C=����Z^}�����4ü�˼~�HAP�$��W+���#������V��Lj!��.����t����ܽrT��*��:�2�$=༬1��,�� >�x$a�0�ҽz6�Ť���>㾸�&�=�j�n���zz˿R����*�1�"�I��i^�V?l��   �   4[�ܣV���J�J�8���#�$����k��#���A�Y��D��Ծ���E/���Խ�W����.�7���<�����	�����̪���4�"�O���d��q���u���o��;a���J�� /�������gZ����f����vS ��F�h��jȽ��(�Շ�`�о�n���W�؏���(����0����#��]9�$1K��W��   �   F5A��s=�RY3��M$�`���t���ѿ����U���JA�w	��λ��4w�����sȽ,߇�"T`�v�s������Pٽ�U�y=�n�j��u��)���S��i귾�׺�rӶ�|E��4�������c�`�5���
�L�ʽ��>�Y��/H�_!y��ʽ�n��<:r�MY��RC��/@�6灿Ok��T�ѿ�>��>��1%�V44���=��   �   �&���"�R��<�������ٿ�Z���_����_�R�%���à��DU�f����������ۓ�)��0����k(�(�_�)G��]����Ͼ�J��<�4�^
�^��������辻̾&��gC��NUX�Sh!�,���w��c��x-������[��y�Q��G��-��%1%��`�����,��tEۿ����  �<���#��   �   $6�4��
��"��<vԿ����8���r�6�9�^���¾�-��>3����LY��O�����Ľ���-�4�.�v�o뢾3NϾ�����S�,A)�H�8���B�o�E�Y�A��?7�
-'���������ʾ����.�o���.��;���绽5m��dE���4�#i1�򞄾����Z	�al:��|s�����q_���zֿ���D���-	��   �   ����޿�ӿmT¿�����ct�7B��^��ھ��� �U����(ؽlŹ���Ƚ���e�4�c�|��Z���㾅��"�/�N,N��i��~�0���ԥ��
��B|��f�g]K�~�,�4���߾���aw�F~0�����ýfH��ֽ�P�CeV�����?�۾����D���v�X���1|��>Ŀտ.�߿�   �   w˲�(r��r��?�������f���=���'j�R~��_n��&�kZ���½"�ý��򽡸(�zq�A����s羲��C@�
�i�mƈ��8�������+��gβ�u���t����������f���=��n�0���bn���&�8]��½ܙý&�򽰵(�q�����o����@@��i�Ĉ��5��躧��(���   �   D�������|�!~f��YK�+�,�w��U ߾����\w��z0����]�ý8H���ֽS��hV����О۾���D�zw������~���@ĿտZ�߿���$�޿�ӿ$W¿����𓿙ft��9B�#a��ھ\����U�e��L)ؽ�Ĺ� �ȽW����4��|�W��B㾘����/�>(N�9i��~������   �   .�E�0�A��;7�q)'�X��T���>�ʾ\�����o���.�H6��>份�k���E��'7�ik1�Ǡ������C	��n:��s����a��N}ֿ���޹��/	��7�֨������xԿн��
����r���9���c¾b/���?3����Y��U���҃Ľ|��ע4�W�v��碾tIϾԧ���P�r=)�?�8�d�B��   �   �Z
� ������Z���̾�����?���OX�d!���齨s���`���,��`��������Q��I�����3%�`������.���Gۿ8���x!�ؕ���#��&���"�����������ٿ_\��_a����_� �%�d�vŠ��FU�T������6���ؓ�h
��l���jg(�A�_�|C�����]�Ͼ7E쾤9��0��   �   �Һ��ζ��@���/��H��~�c�7�5�t�
���ʽB��Y�f,H�� y��˽�����<r�[���D�e1@�e聿�l���ѿ�@��z���2%��54�X�=��6A�@u=��Z3��N$�����v����ѿ����V��RLA�"x	�Fл��6w����<tȽCއ��O`�^�s�g���JٽSQ��s=���j�r��� ���N���巾�   �   �u�Y�o�q5a�;�J���.�t��ǒཤT����f���O �� �"�h��kȽ�(�&և���о�o�)�W�ِ���)�������#��^9��2K�:W��[�Z�V�P�J�t�8���#���E��y������~�Y��E�. Ծ���/�(�ԽW��t�.�2�P�<�������$��B����4�G�O���d�t�q��   �   %f!��*�ˋ��~�f�ܽO�������2��1�h)���&���;似$a�*�ҽw6������?㾙�&�m�j�1���i{˿s�������1��I��j^��@l��q�
	l��)^���I���1���77��Ϳ8A��oUm�])�;|�&x��D=�ʍང]}���� .ü4˼B�^9P�K���%����B	����8���   �   r�㽈�ܽ�̽�岽Ls��\a�*�������.�p餻h��v���^�
�ٽ��>� N���*���/�ouv��{��21տz`�^�(�:���T��Yk���z�J��ړz�@jk�ZJU�ph;�JK �Xl��D׿�`����y�i2���󾕉��l�F����6�{�ȵ�����2M�H˓����w6��;z��J��8����:ҽ;��   �   2ŽB����Y���P��==w�n�7����5{� ����#}��,��0f���X]��:ܽ��A�q���`F���2��z��!����ؿTn���!���=���X�H�o�������d��~p��SY��>�p�"�����ڿ�+��/~��5��H��uV����I�Z�뽦�{����8�T�0��`�N�0���fm��P�[��,㠽�^��B����   �   p�㽍�ܽ�̽�岽Js��Va� ��H����.�椻���t��$^�̬ٽ��>�gM��u)�8�/�ftv��z��Y0տ�_�r]�\�:���T��Xk�h�z������z�ik�XIU��g;��J ��k��C׿`��ſy�Ch2����Ԉ��i�F�6��x�{�\���H���0M�|ʓ�|��w6��;z��J��.����:ҽ;��   �   (f!��*�ы��~�i�ܽ O�������2��0��'��<$���7伞!a�ҽ�6�2����=�$�&�q�j�羝��y˿u���~�|�1�L�I��h^�4>l�\q��l��'^���I���1�Ȋ� 5��^Ϳ�?��_Sm��[)�z羶v��2B=�A��0Z}�����*ü˼���8P���t%����:	����7���   �   �u�`�o�y5a�B�J���.�p�����pT���f���^M �����h�nhȽr�(�9ԇ�"�о�m�e�W�����'��I �l����#��\9��/K�:
W��[�T�V���J��8���#�8��g��"�������Y�}C�BԾ���^/���Խ�T��N�.��/�Ԙ<�T��V�����%����4�<�O�|�d�r�q��   �   �Һ��ζ��@���/��J��~�c�/�5�\�
���ʽ�퐽��Y�)H�Uy��ǽ�����7r��W��9B�.@�8恿j����ѿ�<�� ���/%��24��=��3A��q=��W3�L$�"���r�� �ѿ'����S���HA��u	��̻��1w����pȽrۇ��K`�րs�����~IٽQ�ps=���j�
r��� ���N���巾�   �   �Z
�"������`���̾�����?���OX��c!�L�齇r���^���)���}��M����Q�F�����v/%�P `�����%+��]Cۿ'��������@�#�4&�8�"������������ٿ�X��O^��	�_�W�%�
뾽����AU���^�������Փ� 	��z���g(��_�dC�����P�Ͼ.E쾢9��0��   �   /�E�3�A��;7�s)'�Z��U���:�ʾQ�����o�6�.�*5��d⻽�h��BA��f0�af1����Y����	�j:��ys�Ծ��G]��$xֿ��𿺶�4,	�v4����v��6�sԿS���>����r���9�g��¾�+���:3����nT��4�����Ľɧ�_�4� �v��碾[IϾ�����P�n=)�?�8�e�B��   �   E�������|�&~f��YK�-�,�u��K ߾���_\w�]z0������ý�C��Uֽ8N��aV� ����۾S��D�&�v�;����y��e;Ŀտ�߿����޿�ӿ�Q¿����쓿P_t�4B��\��ھ]����U�����"ؽ9�����ȽV����4���|��V��"㾌����/�8(N�6i��~������   �   {˲�*r��r��B�������f���=���j�0~���n�(�&��W� �½/�ýƟ�L�(��q�����k�X�E=@��i�����u3��.���&���Ȳ�Go��So����������f��=����e�{��in�*�&�ZT��½��ýg��ȴ(�pq�嬩�go���v@@��i�Ĉ��5��麧��(���   �   ���	�޿�ӿpT¿�����ct�7B��^�~ھ��u�U�����$ؽ6����ȽH����4�͚|��S�������@�/�S$N��i�/
~�"������� ���|��yf��UK���,������޾��
Ww��v0������ýC��jֽ�O�zdV�P����۾y���D���v�T���/|��>Ŀտ1�߿�   �   $6�4����'��>vԿ����9���r�4�9�U���¾�-��*=3�
���T��س��~~Ľ��t�4���v��㢾�DϾO���VM��9)�L�8�;�B��E��A��77��%'���������ʾ������o��.�/��j޻��f���@���1�%h1���������I	�Vl:��|s�����m_���zֿ���F���-	��   �   �&���"�R��>�������ٿ�Z���_����_�M�%��뾮à�1DU�B��@���]����ӓ����\}���b(���_��?�����Y�Ͼ�?쾐6�}-�gW
�ށ�������辶̾����G<���IX�^_!�����m���[��>(��~��'����Q��G����1%��`������,��qEۿ������<���#��   �   H5A��s=�TY3��M$�b���t����ѿ����U���JA�w	��λ�34w���"qȽ$ۇ��H`��zs�􎞽5Cٽ�L�Jn=���j�cn������bJ���෾�ͺ��ɶ�m<���+������c���5��
���ʽ�落��Y��$H�[y��ǽ�����9r�Y��DC��/@�3灿Mk��R�ѿ�>��>��1%�X44���=��   �   6[�ޣV���J�J�8���#�$�����k��$���@�Y��D��Ծ����/���Խ�T��@�.��+�t�<�����������ס���4���O�K�d���q�\�u���o�0/a�x�J�h�.����0��NN��X�f����>H ����v�h��hȽ%�(��ԇ�A�о�n���W�Տ���(����0����#��]9�"1K��W��   �   �q��l��(^���I���1�|��M6��WͿ�@���Tm�j\)�f{羑w��:C=�L�མZ}�����%ü0˼�	��1P���� ���轴���,��b!��&���S{���ܽYI���
����2��$�|��x��X3伴 a��ҽ6������>㾳�&�:�j�m���xz˿Q����(�1�"�I��i^�X?l��   �   ���<�z��ik��IU�h;�K �$l�UD׿�`����y��h2�X��_����F�����{����L���)M�lœ�ě�ns6��6z��G��ܑ���6ҽj
཈�㽫�ܽ$̽Dⲽ(p���a�n��x���X�-�@Ӥ��	�<r��t^���ٽ�>��M���)�k�/��tv�2{���0տ&`��]���:�T�T�FYk��z��   �   ��V�8�R�n�F�t�5�H� �<G
���H���Ə�ɑU�����ξ\g���%�{��<������� `Q� 3����O� �ļJ���G�as��`���,��~��궏�ƚ����Y�J�&��oܼ�GW��Oe�X�<�EA<�E<�}л8�������B�*��Fɾ���kAR����F�����Nq	�R4 ��I5���F���R��   �   d�R���N�\lC���2�&-�h�S��5����^����Q�nC�v0˾���kB"��ḽ�<��H���{߻�����-�p���^a ��59�d�p�6���������]��.���R��!�شO�2��O���u㻠�Y;X�<8�;`������i㢽���R�}�h�ž�e���N������״��#�^T�
��.L2��aC���N��   �   ��G���C��_9�̨)�v��ҙ�lؿ�ʭ��b��:LG�G������;z�`$�����&�<��-�� �`��o��m��&�y\�8c��4k���׽e������ �|���?��P5ʽ���'��N1�<�мؾ8� Y/�@s� nA�4��b���d���p��ӻ�'�i�D�<���w����ֿ�/�t^�ֶ)���9��D��   �   b7�.�3�X=*�h&�^�
�^+ￃ?ǿ ����v���6�"��>&��� e�=��^%��@����!Ӽ���TZC�DR��BJ��|��R���v)�l�:� �E��oH�|3C��M6� �"���
���߽2���k��U� ����s�𜼖Z��Ȕ�vO���\�@D���b��H�4��'u�B��S�ƿq￬�v����*�(�3��   �   ��"�`��X��4n�C/����տNα�j���&[���!����}����J�����4Λ���I��"��B3�\�r��׫�d�����@��e�tb��\*������h���֖�����u���~]��E7��C�f�ֽ�d��tI�F:�H%���x'�@��K��TED����~s⾂� ��ZZ�'A�� ��OjֿI����\d�B ��   �   l��PQ
��e���׿Z��e����t�h�;��(
�q.þ�}���s-��޽ ��L:^���]�|���6Ľړ�<�7���l�O���լ�6�ľ�<׾���Jc�q᾿�Ծ���5T��|�� wb���-��m��fV���rv�&>�R B��҅�)�ӽ�)��������	���;��u�l��.���ؿ�W�$���
��   �   U�쿱s�n�ܿQ�ʿ>������N���K�~"����g��_�Y�l/�i�������r��Dח�:�Ͻ���~�J�݆��T���oӾ&`��؂������"�hs%��"����]�ok��4:ξH1��� ����A�,s
�01��^<��^~k�5˃��V�����Q�X�S��F2������L��Ѐ�3��������̿�E޿�L��   �   Z�������o��՘��	ґ��4y�M�V"�s���.~��A�}��-�ξ齤��������T��.ͽ�
�IQO�2���{輾2S�
����,���C���U���`�,Gd���_��S��?A�S*��&�=!�AJ������ĎH��h���ý/G����������x�-�����7��H���>3$��O��>|����M@���Ŵ�cս��   �   �8���S�����ޠ��J)c��UA�[i��������ʏ��OA�������ې�������[���S��
E�:1��\o������!�$PD��Kf������������2;��PV��b������-c��XA�l��������:����"A���2 ������죔��X��XQ��E��.���k��W����!��LD��Gf��������D����   �   �Bd�B�_���S�<A�*��#��뾑F��������H��e���ýJE���������H	�P�-�����:��Q����5$�*�O��B|�<����B��Wȴ�ؽ�������2r��.��� ԑ�B8y��M�}X"�(���ꀴ��}�W-���齺���'���~R��
�̽���LO�'����伾AN�����,��C���U�\�`��   �   �o%�O"�@��Z�f���5ξ~-������!�A��o
�p,��p9���{k�r˃�nX�����i�X�YU��}5���L�L�8Ҁ�3��������̿dH޿|O�2��zv��ܿ��ʿ+@��ٖ��q��d"K�r$�����i���Y�1���������p���ӗ��ϽN����J��ن��P���jӾ�Z����D����"��   �   �]澌kᾏ~ԾQ���P�����=qb��-��f��Q��~kv��!>���A��Ӆ�T�ӽ�)�����[�����	��;���u���%��N�ؿZ��%�b�
�����R
� g�Q���׿-︿yg��Q�t�U�;�
*
�t0þ.��tu-�[޽@ ��8^���]�x���{�ý���C�7�a�l�����bѬ�U�ľ�7׾����   �   �d���Җ�Ӷ��v��Zx]�v@7�&?�P�ֽs_��RI��4����w'��@��|��FGD������u�� ��\Z�mB�����lֿ'K�� ��e�hC ���"�������No�/1��b�տ�ϱ�8k��^([�>�!���;��E�J�I����Λ�n�I�."�t<3���r�ҫ���F���@���e��^��y&������   �   �iH��-C�nH6�I�"�^�
�P�߽����k�(N�����s�으dZ��ɔ�yP���\��E���d����4�<)u�C����ƿ�ￎ�v����*�V�3��7�V�3�f>*�X'�,�
��,￣@ǿ� ����v���6���A'���e�����%��$@�����ӼZ��RC��L���C���������q)��:�_�E��   �   b� ��������@/ʽ*�����n1���м��8��/� N��iA�n��2��je���p��Ի���n�D�����x����ֿn0�_���)���9��D�|�G���C��`9�z�)�
��L��1ؿ7˭�c���LG�ȓ������<z��$�1�����<��*��ȧ`���o�<c��X��p\�N^���e���
׽f^��
���   �   :Z��ؘ���N��<�����O���LH���]�`�Y;��< �;������ 䢽3��4�}��žf���N�򭋿Kش��$ῲT�j���L2�4bC��N���R�X�N��lC��2�n-������x����^����Q��C��0˾����B"��ḽ <��F��@p߻�����"�����:] �"19��p�.���������   �   u��㶏�ʚ����Y�d�&�,pܼ�HW��Ze�d�<�DA<|D<�л���Z����B�V��BFɾ����AR�:���c�����^q	�b4 ��I5��F���R���V�2�R�d�F�f�5�:� �,G
���*����ŏ���U������ξ1g���%��z���<����p���KQ� 1����O���ļ��G��`s��`���,���   �   7Z��ؘ���N��:�����O���(H���\�@Z;|�<��;`���|���⢽^����}�*�žse���N�]����״��#�*T�Ƭ��K2�XaC��N���R�b�N��kC�"�2��,����⿵���Q^����Q��B��/˾E���A"��฽d<�TD��`i߻���� �𵘼�\ ��09���p����|�����   �   _� ��������@/ʽ(��s��L1��м��8�@/�`<��bA�������c���p��һ�����D����=w����ֿh/��]�0�)��9�D���G��C�&_9��)�ȋ�<��jؿ�ɭ��a��.KG������/:z�$#�����p�<�0&����`�`�o��a����<p\�^��ne��b
׽R^��
���   �   �iH��-C�qH6�K�"�`�
�B�߽�����k��M���h�s�$眼�V��Ɣ�EN�t�\�1C��ha��@�4�"&u�"A��<�ƿ"������v�*��3�27��3�<<*�d%�x�
��)�+>ǿ������v��6����$��r�d�����"����?����Ӽ����PC��L��bC��t������q)���:�X�E��   �   �d���Җ�׶��}��\x]�q@7�?�&�ֽ_��6I��2�$��s'�b=��6��YCD������q�9� �&YZ�@�������hֿ0G����&c��@ �,�"�����m�)-����տ�̱��h���$[�[�!�X��H|��6�J������ʛ�@�I�� "��93���r�mѫ�e�����@�z�e��^��r&������   �   �]澏kᾒ~ԾT���P�����/qb�ԇ-�^f��jP��piv�z>���A��υ���ӽd)�����������	���;���u����a����ؿ+U�<#���
����O
�zd�q��e׿`븿Bd���t�2�;��&
��+þ |��q-�V޽'��V2^���]����z�ý�����7�$�l�z���QѬ�H�ľ�7׾����   �   �o%�Q"�C��Z�f���5ξx-��������A�uo
�h+���7���vk��ǃ��R��Z��%�X��P��V/�����L��΀�U���򵿌�̿C޿�I�}���p迻�ܿ��ʿ�;�������~�K�K ����We����Y��,����i����m���ї���ϽΉ�.�J��ن��P���jӾuZ����A����"��   �   �Bd�D�_���S�<A�*��#��뾇F������Q�H�te�5�ý�B������򲣽� �V�-�O���4�������0$��O�;|�퀓��=��*ô��ҽ�����;��m��j����ϑ��0y�BM�tS"�R���{����}�C-�>��ێ������O��!�̽��RLO�����d伾$N���|�,��C���U�[�`��   �   �8���S�����ࠀ�N)c��UA�\i�������������A������f���ş��T��bN��E��+��[h�������� �WID��Cf�v��:�����(6��]Q����������Q%c�3RA�vf�����������A�o��n�����2���9V��xP�+E�\.���k��9����!��LD��Gf��������E����   �   \�������o��ؘ��ґ��4y�M�V"�g���~����}�7-�߼齙���$���N����̽�CHO�3����༾�I�3��-�,�-�C�l�U��`�f>d��_�׭S�G8A��	*�	!��뾕B������ŅH�1b���ý_@�����ճ���齸�-����Y7��$���23$��O��>|����K@���Ŵ�eս��   �   W�쿳s�p�ܿT�ʿ>������P���K�z"��㾲g����Y��.����ރ���l��@ϗ�+�Ͻ����J��ֆ�M��fӾU���|���i�"�/l%��"����W�`���0ξ)��O�����A��k
�&��N4���rk�/ǃ��S�������X��R��"2������L��Ѐ�/��������̿�E޿�L��   �   n��RQ
��e���׿[��e����t�f�;��(
�W.þ�}��/s-��޽���$1^���]�����J�ý��O�7�H�l�����"ͬ���ľx2׾t��X�	f�NyԾ{����K��5	��kb�ق-��^���J��$av� >��A��υ���ӽ�)�н��������	���;��u�i��+���ؿ�W�$���
��   �   ��"�b��Z��6n�D/����տOα�j���&[���!����}��D�J�&����˛���I���!��43��r�̫�g콳����@�L�e�T[���"�����r`���Ζ�����\��r]��:7�:���ֽ8Y��^�H��,�(��Pq'��=������DD�꥘�^s�x� ��ZZ�%A������OjֿI����^d�B ��   �   d7�0�3�Z=*�j&�`�
�^+ￃ?ǿ	 ����v�}�6���*&��G e�����#����?�8��Ӽ`��ZIC��G��P=��$��~���l)���:�́E�TdH�V(C�C6�\�"��
���߽p��*�k�*E��䯼��s�|᜼\U��Ɣ��N���\� D���b��A�4�|'u� B��R�ƿq￬�v����*�*�3��   �   ��G���C� `9�̨)�v��ԙ�lؿ�ʭ��b��9LG�D�������;z�$�ڗ��ڏ<��$��0�`��so�$X�����h\��Y��`��^׽�W����� ��{��z�)ʽ����2�� 1�p�м �8���.�@� [A����:��2d�H�p�qӻ� �e�D�;���w����ֿ�/�t^�ֶ)���9��D��   �   d�R���N�\lC���2�&-�h�S��3����^����Q�mC�q0˾���AB"�pḽ�<�D���b߻@�������ZY ��,9���p�F���b������V�������K��@���B�O���@��pA��,Z;��<8$�;м��ئ��⢽v��3�}�_�ž�e���N������״��#�^T���.L2��aC���N��   �   
�-�t�*�z�!�Е� ����RS���ɗ���i��,������祾z>V����x���`��*��XV:`q|;@��:�з�@Em�T�ż�		���)���A���N���N���@� �&��\��E�� �`Sd;�$g<�(�<vB�<p�<��<��h�_Y�Tl��G��L���f�E�)�j�f�n@��-滿T���DX���!��*��   �   z�*�p�'��/�D+���~�߿&=��TB��?�e�@�)��^�5䢾@R������������8���s� H�:`�1�x�+����|S ���*��O���j�n�y��Bz��l��O�v�'��9�@ف���5�L�<��<�$�<ز�<T�	<�=l�8V��M��fD�����Q�q�&���b�ٓ�p�����޿�����)���'��   �   �j"�
��4��3�C���<տ{D��Y鍿�EZ��!���N(����F�r��Y������Jb�@�ϻ`:��i��JмN��ȢZ�g���^!���������{��Vk���\�������U`� E��`�� zݻ�c�;�3O<�X<0�;0�y���L�ьԽ�:��n���s޾��P�W�q֌�/a��,�Կ�p���=���(���   �   ��������Tj �a�俏�Ŀ�8���j��M/H�]f��о�����4���۽�My�:m��U�������L��26�XR�:���i߻�G�佗�2������P�b��)�\)��̽������`��
�d+�� �_��;@�ܺ�����b@���½�*��ه��˾����F��́��ڢ���ĿK��� ����=��   �   ���:g�X���t��.̿�i���K���g� <1�l)�PK��w�o������H�c���
��'׼|���%1�)f��1�����Y��'6��\P��d�\�p��(t���m�#T^�_3G�Jw*���
�TԽ�m���\A� ܼ�sj��_<��%��8�3�.\��R!�%�o�bq����b�0�TLg��t��o꯿ Ϳ��濒������   �   ��翯�㿹Vؿ��ƿ�~���E��
�y��mF�^�\�ݾ���E�P��8��k���P�ֵ��$���L�5ؔ���Խ���8<�ui��/��GU���>��:|�����nݳ����̘�"����\�(.�7V�����o���D�ϼ�^ؼ8�*��閽�+ �wL������ܾqs�HG��{�i2��P����ȿ�mٿ�a��   �   �¿a��U��IW���[����{��.O���#���� �����}���)�(�ڽ�%��z�D��R2�h�Z��d��>w������V�뉾�����fȾ ��n����!�."�zF�ͧ���߾��¾Ps��n����I�<�v˽nT��ڴ3�4��ȴ)�n ��MԽ,"(��}��[������B>%�\Q��7~�:���ʷ���u��W����   �   ׿��z�̯���E��	2m��I�:x%��Z��.žU���L�F�,V��~��� k�:FB��0Z�h�z����"���b�9�����\���r��(���,���5���8�F 5���*���������f ��0���4wX�N}��н���x�D�3��b� ���(y�n5I�y��ȾTD�M�'���L��p�G����Ó��Z���   �   GAv��lq� yd���P�#�7� ��J��v&Ǿݥ��t7W���?�ĽA�����H�)L�}�����̽���k^�ə���˾�����s�:�:S�uf���r�zEv��pq�}d�R�P�L�7�����"��*Ǿ����};W�r���Ľ]���H��'L�5�����̽���^�4ƙ���˾ ��Ӣ�#�:�k6S�qf�v|r��   �   �8���4�L�*����;��X�澗��)����rX��y��
нr��2}D��3�v�b�����x{��8I����N"ȾtF���'���L�tp�Q����œ� ]��%��Ě����G���5m��I��z%��\��1ž����x�F�JX�b����"k��EB�H-Z�헽Z��*�"���b��5���������o��%��,���5��   �   9��C�T����߾��¾�o���j����I��8�Rp˽mP��Я3�����)��!��2PԽ�$(���}�i^��R����@%�+Q�;~�#���蹧�;x������S�¿���DW��PY���]����{��1O���#��"�����3�}��)���ڽ�&��t�D�6P2��Z�\`��Hq����~�V��牾ɢ���aȾ����������   �   X���س�c���Ș������\�K.�PR�����o�R���ϼ�[ؼ�*�H떽z- ��yL�{��^�ܾ6u��G��{�4��2����ȿ�oٿd��������Xؿ��ƿW���*G����y��oF��_���ݾ������P� :�jm����P�$��� �h�L��Ӕ�[�Խ��v3<�bi�,��LQ��x:���w���   �   �!t�X�m��M^��-G�1r*�S�
�Խ�g��tSA�<�ۼ�`j�U<�$$��x�3��]���"���o�/s�����0�sNg��u���믿�Ϳ��濡���*�����Hh�U���D�忬/̿^k��M����g��=1�}*��L��w���������c���
�4"׼Ԫ��1�na���*��(��U��"6�WP���d���p��   �   L�y]�<%�S!���̽ѥ��&�`�lw
�4���>_� @;�]ܺ���Ld@���½	*��ڇ���˾'��	�F��΁�ܢ�ДĿ���Դ �����>�t���	�j��k ���俱�Ŀq9���k��z0H�:g�3о񗌾��4���۽�Ny��l��Q�������B��z/��R�惑�ٻ���~ �Ȏ����   �   ,u���e��W��v����L`�V=�TS��`Oݻ���;(@O<�	X<��;��y��L�+�Խ�:��o���t޾��g�W�׌� b���Կr��\>����֫�`k"����΀��3�1���J=տ E���鍿jFZ�n!�����(��l�F�2���Y��@��@Eb�nϻ� �8~i��?м�����Z�����6��������   �   �<z�@l���O���'�D1�с�`�5���<��<�'�<���<��	<�>l�8V��N�~gD�B����Q���&���b�jٓ������޿
��Z�**�<�'�ؾ*�ʼ'�(0��+�V����߿p=���B����e�|�)�_�h䢾@@R��������x��� 8���s��~�: �1�8�+���zO �L�*��O���j�­y��   �   t�N���@� �&��\�F��p��Qd;$g<�(�<B�<��<P�<��h��_Y��l�J�G��L��3g�l�)���f��@��I滿%T����NX���!�"�*�
�-�p�*�r�!�ƕ���v��:S��uɗ�S�i���,�J����祾2>V����mx���`���*� jV: u|;���:�η�pDm���ż�		�~�)���A���N��   �   �<z�0l���O���'�1�с���5�0�<t��<<(�<���<��	<�9l�fV�$M�xfD������P�9�&���b��ؓ�*���5�޿������)���'��*��'�|/��*������߿�<���A����e���)��]�㢾*?R�l�����������7� cs����: �1�`�+�P��$O ��*���O�f�j���y��   �   u���e��W��r����L`�8=�S�� Mݻ���;�BO<�X<@ �; |y���L���Խ�:�dn���r޾�����W��Ռ��`��m�Կp��>=�|�����j"�\����p2�(����;տ�C���荿�DZ��!����['��Y�F�Q���W��f���<b�0aϻ��0zi�>мȴ��Z���������������   �   �K�r]�9%�N!���̽������`�
w
��� 0_� V;�ܺ|���X_@���½Q*��؇���˾7��v�F��́�ڢ�r�Ŀ��J� �D���<���������i ���B�Ŀc7���i���-H�:e�Hоᕌ� �4���۽�Hy��h��K��<���\?��.��R�e����ػ���^ ����ښ��   �   �!t�S�m��M^��-G�-r*�K�
��Խ�g���RA�,�ۼhZj��J<�H����3��Y������o��o������0��Jg�ks��鯿��̿ו濜���
�����&f�G������Q,̿rh���J���g�h:1�(�_I��2w�K��0���Z�c���
�׼����1��`��J*������T�n"6��VP�l�d���p��   �   T���س�b���Ș������\�;.�4R�&���o���ܪϼPSؼ��*�j施�) ��tL��	��X�ܾ�q�AG�D	{��0�������ȿ_kٿq_�?��^��}Tؿw�ƿ�|���C��6�y�{kF�F\���ݾ�}��4�P�f6�1h��,�P�ܮ���v�L�jҔ�u�Խx�$3<�i��+��9Q��j:���w���   �   6��C�U����߾��¾�o���j����I�8��o˽�O���3�l��Z�)�����HԽ|(�J�}�^Y������.<%��Q��4~�k���µ���s�������¿	���R��+U���Y��L�{�$,O���#���`�����}���)�X�ڽ�!���D��J2�.�Z��^��*p�}���V��牾�����aȾ���������   �   �8���4�N�*����<��V�澒�����crX��y��	н���xD�"3�ؘb�䍫�}v��1I� ���ȾTB���'���L�Kp�P���e����X������5��������C��c.m���I��u%��X�,+ž��`�F�*S�z���k�0>B�(Z�/뗽��ར�"�N�b��5�����d���o��%��,���5��   �   HAv��lq�%yd�P�$�7� ��F��n&Ǿ̥��:7W�8� �ĽQ�����H�D L����޷̽h���^�aÙ�K�˾۾����:��2S�5mf�Yxr�=v��hq�,ud��P�ڨ7�G������"Ǿբ���2W����Ľ����N�H�� L�ϭ��7�̽���^�ƙ���˾��Ţ��:�d6S�qf�u|r��   �   ؿ��{�ί���E��
2m��I�:x%��Z��.ž<�����F��U�4}���k�n>B��%Z�k藽v��Z�"���b��2���
��Ξ�6m��"���,�_�5�}�8�)�4���*�{��m���澊������YmX��u�cнf���tD��3�&�b����ix��4I�E���ȾDD�@�'�~�L��p�E����Ó��Z���   �   �¿d��U��JW���[����{��.O���#���������}�h�)���ڽf#��އD�0I2���Z�D[���j����H�V��䉾힩�y]Ⱦ��R�����B��@�Ȝ��x�޾��¾�k���g��x�I�a4��i˽K���3�0����)����XKԽ�!(�r�}��[������5>%�SQ��7~�7���ȷ���u��Y����   �   ��翲�㿺Vؿ��ƿ�~���E��	�y��mF�^�O�ݾ�����P�.8�:j����P�������L�<Δ���Խ��d.<�Ti��(��[M��/6��0s�����kԳ����Ę�,�����[�#.�N������o�x����ϼ�Nؼ^�*��疽$+ ��vL�i����ܾes�?G��{�f2��Q����ȿ�mٿ�a��   �   ���<g�Y���v��.̿�i���K���g�<1�f)�@K���w���A���*�c���
��׼`����1�E\���$��p��P�d6�>QP�/�d��p�%t���m��G^��'G��l*�Ê
�@Խta���HA�8�ۼEj� =<� ����3��Z��� ���o�?q����X�0�NLg��t��m꯿ Ϳ��濒������   �   ��������Vj �a�俏�Ŀ�8���j��J/H�Zf��о�����4���۽�Jy��h�4I��̤���6���'���Q�i~���һ��x�k��`��L��VG��X�� �(���̽[����`�,n
����@�^� �;��ۺP����_@���½<*��ه���˾����F��́��ڢ���ĿL��� ����=��   �   �j"�
��4��3�C����<տ{D��W鍿�EZ��!���A(����F����X�����`:b� Tϻ� ��ji��3м|����Z������{���A��Ko���_���Q��T���zC`�5�8E��@ݻ���;�PO<�X<p-�;yy���L��ԽJ:��n���s޾��L�W�o֌�.a��+�Կ�p���=���(���   �   z�*�r�'��/�D+���~�߿&=��TB��@�e�?�)��^�/䢾�?R�p���e��d����7��:s�@��:��1��+�����K ���*� �O�D�j�H�y�B7z��l�p�O���'�(�Ɂ� [5���<6��<�+�<J��<��	<�7l�4V�>MསfD�����
Q�o�&���b�ٓ�p�����޿�����)���'��   �   x�	��j�o� �G��aҿ<���^���®n��6����.���	�����%�  Ƚx�[��A̼����:�s5; �@:����i$�����(����(޼�H��|���D��0Ҽ/���T3��A���Y<�ǡ<�%�<�=}#=Ь=1�<��;�3ټ4͗���a�o�}����P�
4��4l�`����߳�d�ѿ�R�b� ��i��   �   ���&=��D��9����ο俱�2����j�ƪ3���2���0;|��P"���ý$W�p�ɼ�����%���M: 
����~q��ᴼl��*H��u���!�ȑ���l��𗼘���V];��n<@�<N=��=U	=h��<0��;HiԼ
���;�pMk��^��.��1�Sh��>������ο���>���A��   �   $������E�s�ݿſ�%����^��i*��V���s��: n�)�����.�I���¼<�`�������x?1�xu��d��ƃ!���H�fj�C���D
��"h��t�v��W��[+���Hw� ǖ�=<:O�<���<x��<갫< Ս; �Ǽ)���r=�%�^�6��,��<(��]��D��Ǹ����Ŀ}�ݿ?s�W���   �   �_=�œ޿�̿\������������RL���>���Ơ��*X�[�	����6�p���p�M��3��_����Լ�w ���]����P��o�Ž��ؽ>����źؽ��Ľ�v��&���$@���XA0�p�;�5i<�z�<9{<��!;�b���s|����2K�F���ܯ�,|��HK�*L�������յ���̿4 ߿����   �   տzQѿ��ƿm���
ۡ�Ny��48d���4��	��Gɾ��On<��W��� ��P���玼hi���J��[F�驌�º���+����!�-�Ǆ6�J�7���1�d�$�ԟ�����俽@Ŋ��1�X᲼0������;`G�; �l�o��"&\���Խ��2��U����ƾU���4��}d�2܊�t���6��Boǿ-�ѿ�   �   W����������lw��^��N�m��pC��f�N�O���W^m�Y�.�Ž��k��%��Rż$+μ�b��C^�8O��0s߽�h�m4�f_U�$�r������O��,󌾬0��cP��;f�T�E��H!�.�������g��3���d��C���^л�ǝ�j�:��9��f�:�i�ݻ���꾀���D��\o��D���d������6q���   �   
�� 0��7L��?"��*�g��D��J!�2���7���a���4T?������Ǜ��<��H����d�H�b����
���
�%��U�vv��\J��hV��8���T�ʾ��;��Ⱦ�ϼ�\����+��]v�YC�°�.-νXS����@�8jl��r��t��Ϥ�����bT?����������X ��#�mG��i��4��&�������   �   �Vx���s�Txf��pR�c>9��
�B �:�Ⱦ�~��E�W�p���߼���h������ȯ��nS�:�������9.�V�i�|���^�����ؾO����`�J��2�����*�����>GҾ�}�����r!Z������ٽh�����&���м�X�������e��������]��F��N; �����n�;���T��:h�wt��   �   n�@�Q�<��P2�&i"�G}�v��-"þ�����Ea����b7ӽ4w��*�"��<弐6𼪳2��N���%���(��l�rѝ�gsɾ�����f���$��4���=�ʥ@���<��S2��k"������%þV����Ia����<ӽXz��П"�d?弬4�N�2��K��0!佋�(��l��Ν��oɾ<����c��$�o4���=��   �   R��΋����ͫ��BҾ@z�������Z����`�ٽd�����&���м�W��J��� f�:�������]�fI���;5����Z�;�1�T��>h��zt��Zx�.�s��{f��sR�.A9�a�< �_�Ⱦ���ۛW���!㼽�h�r�0��F���iS�N������5.�\�i�]�������L�ؾR���+^�s��   �   �;��ȾP˼�h���v(��Wv�'TC�Ȭ��&ν�N��*
��窼�al��r�����,�������FW?�����v���`Z �+#�G�*�i��6���'��|������2��N���#���g���D��L!���������D����V?�9���Gʛ��<�|I����⼄� �b������� �%� �U�gs���F��`R��ձ����ʾ�   �   �!-��M���4f�߂E�D!�\���2���g�J,�p�d� )���Sл�ȝ��:�"<��e�.�i�𽩾Ս�M�F�D�I_o�iF��Of��l���s���X��i ���«�
y��w_����m��rC��h��P�-���am��Z���Ž$�k�x&��Pżt%μ�]�p<^�bJ���l߽�d��4��YU��r�C���XL���   �   ��7�l�1�h�$�=��V���ݿ�P���:�0�Ҳ��r���ќ;PZ�;��l��p���(\�I�Խۈ2��V����ƾ� 	���4��d�m݊��u��V8���pǿ�ѿ�տ-Sѿ`�ƿ儶�Yܡ�mz��:d�Q�4�,�	�hIɾ����o<�H���X��ڷ �P��䎼tb��fE��TF�0���9���f���+��-�~6��   �   ���n�ؽ��ĽBp��`�@���漠%0� B�;�Ei<P��<<?{<@�!;�d��v|�A��z4K��������N}�HJK�M��¦���ֵ���̿�߿���`��>��޿O�̿l������������SL�������Ǡ��+X�A�	�����6� ���X�M�X�3�X����Լ$q ���]��z��GJ����Ž��ؽ����   �   fc��"�v��W��S+�X����v�����%=<"V�<��<���<���<0Ս;�Ǽ/���Q>�w�^�(��}���<(��]�VE��������Ŀs�ݿEt�h���$������F�M�ݿ@ſ<&��w�����^�dj*��W���t��#!n����������I���¼�8��ꍻ�{��(21��l�����b}!�f�H�(�i�Ҝ������   �   (��������藼x����];d�n<z �<�=ԑ=�U	=���<`��; kԼ�����;�INk�)_����A1��Sh�?��K��q�οu��S?���A���j=�EE�����4�ο/���[2���j�	�3�  �t����;|��P"�"�ýFW��ɼ��� �%��FN: �	�����@tq�$۴� ��D�dq�j�!��   �   ��Ҽ/�� U3��C��xY<Lǡ<z%�<~=S#=��=�0�<P�;�4ټ�͗�M����o������P�3
4�5l�v���೿x�ѿ�R�h� ��i�x�	��j�j� �8���`ҿ(���H�����n���6�ۅ�����拀�X�%��Ƚ�[�A̼� ���:�v5; �@:0��i$�@��������(޼PH��<����   �    ��d�����藼(�� �];��n<� �<% =�=5V	=T��<���;�gԼ�����:�Mk�Q^�� �z1��Rh�h>�������ο���M>��fA�v���<�;D�����W�οo����1����j�;�3�������@:|�P"���ýbW�<�ɼ(���`%� zN:��	����� rq�(ڴ�X�켾C�&q�:�!��   �   Cc����v��W�~S+����v�����&=<
W�<:��<���<L��<�;HǼ����<�0�^����C��u;(��]�,D��+����Ŀ��ݿRr�X���#�}����D�z�ݿ�ſ�$��C��^��h*�XU���r���n���:���$�I���¼�/��ۍ�po���,1�|j�����x|!���H���i�����j���   �   l��K�ؽ��Ľ-p��I��@�|��0$0� F�; Ii<���<�F{< �!;�\���o|����Q1K�D���~��A{��GK�lK��Ӥ���Ե�y�̿��޿?��^�<�^�޿ȁ̿(����������/QL����m�侖Š��(X���	����Ќ6�<����M�0�3��S��еԼ�o �$�]�Ez���I����ŽH�ؽ����   �   ��7�Z�1�]�$�4��A��~ݿ�&�����0��в��j��ݜ; l�; �k��f��~!\���Խ�2�KT���ƾ2��q�4��{d�ۊ��r��X5���mǿ�ѿ_տ�Oѿ�ƿށ���١�x��6d��4���	��EɾF��k<�����T���� ��F���܎�p\���B�tRF�6���]�����Ď�����-�\6��   �   �-��M���4f�ԂE� D!�2������0g�<+��d����P6л轝���:�Z6��F�b�i�����������D�0Zo�xC��c��݅��]o��2U����������u��\����m�anC�e�2K�~�� [m��V�D�Ž �k���@FżTμ�Z��9^�.I���k߽ d�H4��YU���r�+���FL���   �   ۡ;��ȾK˼�d���q(��Wv�TC�����&ν$N�����⪼�Rl��g��n��A�������jQ?����� ����V ��#��G�)�i�Y3��<$��������5.��_J��� ���g�k�D�\H!�����T���*����P?�\����Û��x<��;����^���b��	������y�%���U�4s���F��@R��������ʾ�   �   N��ˋ�~��ʫ��BҾ:z������Z����߹ٽ����6�&���м�L��V��\�e�.���(��J�]�YD��;��%����;���T��7h�tst�BSx��s��tf�emR�u;9�t�" �ȎȾ�{���W�:���ڼ���h�Z����*���eS��������.5.�ܳi�%���c���(�ؾ5���!^�l��   �   l�@�Q�<��P2�%i"�F}�r��&"þw���|Ea�f���6ӽv��ܘ"��2��'��2�LG������(��l��˝�lɾ����^a�/�$�P4�Y�=��@���<��M2�6f"��z���bþn����@a�����1ӽ�r��X�"�p.�(𼒫2��I������(���l�GΝ��oɾ����c��$�i4���=��   �   �Vx���s�Txf��pR�b>9��
�@ �2�Ⱦ�~���W�$���޼�҇h�$����v���aS�G�������1.�D�i�9���Я���ؾd���{[��|�p�����ʂ�̦�}>Ҿev������WZ������ٽ(����&��м�I�� ����e����t����]��F�� ;��}��b�;���T��:h�wt��   �   ��!0��8L��?"��,�g��D��J!�(���,���N����S?������ƛ��{<��=��,��L�8�b����������%��U�Np��2C��XN��t����ʾ4�;T�Ⱦ�Ƽ�X����$���Pv��NC�p���νI��0��ت�hGl��e�������������S?�R��������X ��#�`G��i��4��&�������   �   W����������nw��^��N�m��pC��f�N�A���(^m��X�<�Ž��k�<!��EżμvV�N3^��D��f߽l`��4�9TU���r��}���H���댾�)���I���.f�9}E�%?!����H����f�,#���d�����p%лH�����:�28����Жi�������t���D��\o��D���d������8q���   �   տ{Qѿ��ƿm���
ۡ�Ny��48d���4��	��Gɾ��n<�c�V��t� ��F���َ�|V��6>��KF�֟��Ե����Ί�r��-�)z6���7��1�Q�$�������+ֿ�������0�����@9��@�;���;�k��f��#\���Խ��2�fU����ƾI���4�|}d�0܊�t���6��Coǿ1�ѿ�   �   �_=�Ǔ޿�̿[������������RL���5���Ơ�_*X��	�?����6����HM��3�`M����Լ\i �d�]��u��>D��J�Žp�ؽd��
����ؽ��Ľ�i��`셽v@�����0�0u�;�Zi<0��<O{<@�!;�\��Zq|�@��}2K�(���Ư�"|��HK�(L�������յ���̿7 ߿����   �   $������E�s�ݿſ�%����^��i*��V���s��" n���������I��¼�.�@Ӎ��_��X!1��b���v!���H���i�J���� ���^����v��W�:K+�����v� ^���9=<�^�<
��<���<��<p�;HǼt���0=���^�#����<(��]��D��Ǹ����Ŀ�ݿ@s�Y���   �   ���&=��D��8����ο㿱�2����j�Ī3���/���$;|��P"���ýbW��ɼx�� H%���N: �	����� iq��Դ����@�m���!������� �����X����];o<�%�<"=��=TW	=���<���;lgԼ�����:�WMk��^��*��1�Sh��>������ο���>���A��   �   �BԿ��пj5ƿ�ﵿSE���牿�>c�:4���	��ʾ�鎾��B���FW���";���Ѽ�gg�H����򻀸���4�`�b�����4��Lܛ��Ɨ��F����R��E�� m9����; i�<l�<u�=n>.=��D=�,N=N�D=�"=���<��	�P $�pվ��)�fㄾ�I¾v����1��a�L��9ᠿ���-&ƿc�п�   �   ��п8FͿ��¿u�D������Y_�h1����Xƾ�1����>�m���x��>6� �̼Hmf�p�� D���*�`7_�􌼬&��8r����ɼ@ʼ����89��pi��d� ��:�65<$a�<�-�< =܅9=�hE=�{>=��=>_�<�&���PϺ���%����j徾t@���.�%�]�����G��%Ҳ��¿�LͿ�   �   �ƿouÿ%���;F���Ж�Հ�T���'����������N��~E3��i� T���'� �����e�`�3���G�`*���ΰ�|���P�By�L+�(2��0�p$���L1ۼ�m���K��Т�;@��<ڹ�<��=X�*=8�+=�O=�"�<�|\��
�*��ߐ�X%w�F��P���=&�C�R�����	����R��T�����ÿ�   �   �Q��5���쪿�����s�l��XB�z�����)֪�Ep�*�!��RϽ�u|�����g����l���j�Њ����ּJ��x�:��Xc�����B������F&������C����x��)G�4��ܕ���Rn�h�,<`;�<��<��
=P�<&��< �w9�\ �H7���ٖa�-���"@澫����A���l�nϊ������7��vF���   �   �m���y���1���\���>v�U�Q���+�L��8�;�����P�.�J����"R����+�����(٣���*��g��p���[��r�ӽʊ�|����l�L��2����[��Eý���e�����}� ��:8Gn<bƶ<B��<���< hy:ռW��] ���lF��b��	�˾�W�,-,��XR��.w��ዿ���� ����   �   �ǌ��(���傿']o��S�vF3�`���\�3٭��w{�М-��d��V���$�����>���\�������2������箽�{��[	��!�T�5���D��fM�uIN��G��M8�@#��	�̾ؽ#l��0	N���׼ �Ự]�;@6X<��=< �7:���a^�J�Ͻz"(�x�y�dB����b��3�4�B�T�K�p�f|��}���   �   j�z�e��0Y�z5F�V.�ť�����%���	��A�I��	��ͮ��KP�u�hx���ΐ�ĬҼ��)�+���|���5O��OO"�c�F���i�f��`Ə�S���EC��Y
��pd��Tx�7U�A_.�Z��F����|�F���DZ� ������;@H��8����0�"����6	��&M�vُ��ǿ�,���*��2y0��H���Z�iLf��   �   c~;�ݱ7�Պ-�����
����T|���,��|BZ�y�݅ʽ�fw�jI�Pћ��~p������b�zo�������M0���a��>�������]���)ɾV~Ӿ�G־*Ѿ֓ľ�����<��W?���uK���m�ֽ��������R���ʻ����0�`�������$�׽�"�+Ze��>��кþ���TW�JT �5/�[�8��   �   6��=n�V���msӾ
j��`����[�>Z��=ٽ�.���B� 𚼘�1��V���ϼ�3C�q�����*�0�d�l��:��_���iھ�����K��q�ˑ��p�gX��JwӾVm�����[��]��Bٽ�2��H�������1�V���ϼ�/C��m������ۆ0��l��7���[���eھ����OI��n��   �   1C־�%ѾƏľЬ���9���<��
qK�W����ֽ>���T���I��@�ɻ���p�`�^��W���׽ܽ"��]e�kA���þf�ﾌY��V ��7/�4�8�D�;���7���-�V�#�
�>��Z��/��>FZ��{��ʽ�lw�HM�X՛���p� ���l_�o������J0��a�<��h���;Z���%ɾzӾ�   �   �?�����"a��Nx��1U��Z.�|�����$�|�����.Z� "���ʂ;@;��આ��0�씧��8	��)M��ۏ�pʿ�����2���{0��H���Z�jOf�j�o�e��3Y�	8F�_X.����Љ�M(�����9�I�	�Ѯ��OP��y�<z���͐��ҼP�)��������PI���K"���F�1�i�^��Ï�׽���   �   �CN�MG�\H8��#�r	�z�ؽ�e���M� �׼P�� ��;�AX<p�=< �7:�"���d^�4�Ͻ�$(���y�xD�������?�4���T���p��}���~��uɌ�u*��7炿�_o��S�cH3����_�%ۭ��z{��-��g�Y��:$������>��xY��p��*�2�r� 㮽�u�NX	�b!��~5�e�D�>aM��   �   2�� ���>T��>ý������d�����}� ��: Zn<Ͷ<z��<B��< Ly:�ռ��2���nF�Td���˾Y��.,��ZR�/1w��⋿���}����n��5{��3��^���@v��Q�4�+�s����;k�����P���4���"%R�X��+��H���գ���*�g�Rl��NV��B�ӽ̓������h��   �   �e=�� �x�TG��� �����m���,<\D�<���<��
=*�<���<  w9D^ ��8��F ���a�v����A�ȟ�=�A�R�l�\Њ������8���G��S��Q��������Ƥ���l��YB�m����>ת��p�F�!�xTϽ�w|�ܶ�Lh����l���j�$�����ּ���l�:�,Qc�R���W���6��� ���   �   $����T#ۼ�`��������;��< ��<��=��*=��+=�P=�"�< �\�,�X+��ܑ��&w�E��� ��n>&�J�R� �������[S��!���z�ÿ��ƿ9vÿ㛹��F���і��Հ��T���'�����|���O��BF3��j��T����'�܄�� �e��3���G��%���Ȱ����&L��s�+�L2�v0��   �   �1��8i�@I黀]�:8B5<,f�<�1�<� =8�9=�iE=l|>=�=_�<�7����,к�?�%�����澾�@�o�.���]����,H���Ҳ�{�¿�LͿ9�п�FͿ��¿�󲿍���V���dY_��1�.�Yƾ�1��ؠ>�ԇ��Tx���6�<�̼�lf� ��A�@�*�H1_�����!���l����ɼ��ɼ�����   �   ��R� E�� i9� ��;i�<\�<Z�=\>.=x�D=�,N=$�D=��"=~��< �	�� $��վ��)��ㄾ�I¾�����1�?�a�L��Iᠿ���6&ƿh�п�BԿ��пa5ƿ�ﵿDE���牿�>c��94���	��ʾ�鎾r�B����W��h";�4�Ѽ gg����@����H�4���b����h4���ۛ��Ɨ��F���   �   t1��xi�H� b�:�B5<\f�<2�<� =|�9=jE=�|>=��=�`�< �&���κ�R�%����!徾B@���.���]�Q���G���Ѳ���¿LͿ[�п�EͿ,�¿�ߗ������hX_��1���'Xƾ*1��џ>�I���$w���6�4�̼0gf����<�@�*��-_�x| ��xk��t�ɼ��ɼ䑼��   �   �$�T���"ۼd`��0��p��;v��<���<��= �*=b�+=�Q=&�<�\����(����I$w����\���<&�x�R�
���w����Q������݌ÿ=�ƿ�tÿW���wE��AЖ�xԀ��T��'�#��������M��HD3��g轗R��p�'��~����e� �3���G�4"��xŰ�����J��r�+��2��0��   �   h%=����x�G�Է�D�����m�p�,<XE�<��<��
=:�<���< Jz9jY �h5����;�a�����>澿����A�I�l��Ί�����6��]E���P�����몿��������Ɋl�LWB�T��Ĥ��Ԫ�%p���!�\PϽNq|���`����l���j�h�����ּ*��F�:�DOc������������2 ���   �   ��؃��T㽬>ýw�����d�����}����:�]n<�϶<&��<���<�Nz:ռ���D����jF��a��@�˾�V��+,�1WR��,w�o���u���˼��0l���x��r0���[��]<v�d�Q��+�����;w���O�P�I�H����R�l��!�������ͣ����)�Hg�k��0U��V�ӽ��=����h��   �   �CN�(G�@H8�n#�\	�L�ؽ�e����M���׼���@��;�IX<��=< �8:���d[^���Ͻ' (�oy�f@�����ή�J�4��T���p�{��|��yƌ��'��i䂿~Zo�C
S�aD3�����Y��֭�Ht{�%�-�z`㽠S���$�T����3��$P��8��h�2�����~ᮽ�tིW	��!�9~5��D��`M��   �   �?�����a���Mx��1U��Z.�a��������|�����(Z� ��`�;@�������|0�N���$4	��#M�i׏�)ſ����7���v0�gH��Z�tIf�j�x�e��-Y��2F��S.�������"�������I�* 	��ɮ��DP��h�l��t���Ҽ�)���Q����G���J"�;�F���i�*���������   �   C־�%Ѿ��ľƬ���9��|<���pK�8��0�ֽȫ������E��@�ɻ�p��x�`�4������D�׽��"�.Ve�j<����þ���'U��Q �s2/���8�{;��7��-�_���
����
y���)��B>Z��u���ʽT^w��B��ě��ep�H����Z�o�:�����DI0�>�a��;��.���Z���%ɾ�yӾ�   �   0��8n� V���fsӾj��X����[�Z� =ٽ#.���@��ꚼH�1� V���ϼ(C�i������#�0�c�l�5��PX���aھ����F�il�����k��S�(�doӾ�f��r�����Z�kV�z7ٽ�)���:��⚼��1�hV���ϼv+C��k��D����0�a�l��7��x[���eھZ���AI��n��   �   `~;�۱7�ӊ-�����
����L|���,��^BZ��x�T�ʽ ew� G�ʛ��ip�Ю��<X�^o�����g��E0��a�9�� ���jV���!ɾ�uӾ�>־h!Ѿ��ľ����-6���9��lK�4��آֽ覉����X;�� �ɻ0d��(�`�.��������׽b�"��Ye��>����þd��@W�;T �5/�U�8��   �   j�x�e��0Y�z5F�V.�¥����%���	���I��	�Cͮ��IP�o�o��8��Ҽ��)�G|��F���QB��fG"���F���i�<������H���<��O���]���Gx�,U��U.�V�������|�����Z� ��� ��;����Ԟ���0������5	�f&M�5ُ��ǿ�������#y0��H���Z�fLf��   �   �ǌ��(���傿&]o��S�vF3�]���\�)٭��w{���-�d�%V��0$�ԑ��l4��N�� ��.�2��퀽Dݮ�$o�ZT	��!��y5��D��[M�L>N��G�C8���"�����ؽ^_���M��}׼`|�p��;XWX<@>< �8:����]^���Ͻ�!(��y�1B�����P��&�4�8�T�E�p�e|���}���   �   �m���y���1���\���>v�T�Q���+�J��0�;�����P�������� R�$���"��䃃�(ʣ�
�d�)�g�g��<P��m�ӽL|������d����{��FL�p7ý𣜽&�d����xn}����:�qn<׶<L��<���< _z:ռ ��^���xlF��b����˾�W� -,��XR��.w��ዿ����!����   �   �Q��6���쪿�����r�l��XB�x�����!֪�.p��!�vRϽ0t|�����a����l�8�j��|��p�ּ؄���:�\Hc�l�����|������蚽|7����x��G�����t���pm���,<�N�<\��<��
=�
�<t��< rz9HZ �h6������a����@澢����A���l�mϊ������7��wF���   �   �ƿouÿ'���;F���Ж�Հ�T���'���������yN��hE3��i轵S����'�p�����e�8�3���G�h��,������zF�fm�,+��2��0�j $�0���ۼlS���뷻���;���<H��<��=p�*=0�+=�R=l'�< \�:	�|)�����)%w�1��B���=&�@�R�����	����R��V�����ÿ�   �   ��п9FͿ��¿v�C������Y_�h1����Xƾ�1����>�L����w���6�0�̼hf����;���*�)_�0댼����f��ܕɼt�ɼL����*����h�p-� ��:xN5<�k�<�6�<�
 =�9=PkE=�}>=Z�=�a�<�	�8��Ϻ���%����`徾p@���.�#�]�����G��%Ҳ��¿�LͿ�   �   u;��N{��턒������l���I�$d%�Q���Ǿ�j��SZS����?o̽Y����L�2�t�v ������S��Ȇ���?��\F⼸�Ǽ�祿p4u��u�@@�p`�;�u`<@�<5� =�$=\�D=��_=��r=�z=��r=hW=$o"=vǝ<��*�L�R� �ٽ/�5�{���쿾�( ���#���H��;l�����/{���{���   �   ៚�W藿���}؃���h�sF��w"�lp ���þ𗐾�O�~���ǽ�8��>�F�j��2��T��� h�����@�zG����T�⼜�ļ�����\`�0�� ��9�<�@�<�j�<�=�'7=�mT=�i=�Es=Pfm=̡S=S� =���<(F �܁M��9ս�,2�{������&���*� �3'E�Jh�^������D헿�   �   �
���l���ꈿ~z���\���;���#2�B���e��L�B��Z�&(���:~���5��#�xz��p{�������b��¯����@�����������@���Sr�@�Ļ I{;�&j<xN�<�s=#2=��M=�X]=�B]=I=��=�6�<p��;>�rȽ�n(��~��벾�(�f��vY;���\�s�z����P~���   �   �+��׶��{{���e�X�J�	,������ݾB����4w��K/��R�õ����[��������2�XC��\�
�����L5�BI�paY���d���i��g���[�F�F�ڴ(�����K��С����;2"�<��<�=t8=�A=,�6=NN=�Ɵ<�m���2'��޴��k�U]h����Y۾�?��,�w�J��Sf���{��ل��   �   p�X�k�A	_�0�K�Q33�����~�¾�i��h�V���>�˽A3��X�0�lW���|ͼ��Ѽ�����I��Q?� &g�6]�����r������6��9պ�h5�����������c��#�h7��  ٻP�<^��<�[=�X=��=��=���<@!8�n��^Ŝ����o7M��$���l¾����y���#4�q�L��_��l��   �   W�M�-�I�4�>�u�-����r;��HҾ�z��#w�O�1��7���T���(L� �HD������'ż�O��5�Dp��𗽴߸�.�ؽ%%�������vp�Y�����.���!Խ~���k{��� �07�� �H�̫k<n��<tN�<�P�<��<��0�($߼+ς��{�c7/���x�t����Rվ������y/���?��mJ��   �   w0*��&�Ik��8�=����pӾ�/��uE���,���
�i��	�(���pk�,4��`BǼ���X%a�����ʽ��������-�$�A��ZP�Q!X��X�,�O�G@���)������������X�0漠*�� ��;�o�<ӗ<�uZ< �9�@���WS�󜻽����1N��Q��=����"پb
 �sY������'��   �   Ú����������e�ž�ҥ�j4���bL�����˽hˀ����|K��؝��s ��_g��cݼ��;�8Y����ɽ����
)���L���n��;��Ƃ��`���H���Ĕ�,ኾu�x���U�Q�.����JD½�W}����`R�@$�: h<��< ׹� ��Bk'��#���?齾*&��^� J���=��B$;=��[���m���   �   yо@�ʾ�|���
��?5��R�w��uD�ǀ��HϽ�-��b��3����u� ^�9 #K���h�K�F�l�Fȷ�ת�X�.�d5^�^������,���$�þ��;Aо��ʾ.������8��9�w��yD���NϽ�1��bh��<���v� ]�9 /K�p�h��H�R�l�'ŷ����Z�.��1^��������������þ̄;�   �   �E������,ފ���x�΋U��.�,���>½^N}����@�Q�@��:�r<p�< �ֹ�"�� n'��%��`C�N-&�x�^�4L��q@��v';���V��������Ȟ����H�⾔�žfե��6��VfL������˽�΀�$���R������x �0`g�Paݼ��;��V����ɽ<��`)���L���n�9�����?���   �   �X��O�d@��)����������X���p������;6v�<Jח<�yZ< ��9LD���ZS���������4N�xS�������%پ �g[�����'��2*�N�&�^m��:������sӾ2��h���xE�>������`�i�ҿ	�����k�x5��8AǼ����!a�E����ʽv���_��9�-���A��UP�BX��   �   	U�����&��]Խ����_{�X� �x'�� �B���k<��<�S�<�S�<l�< 1�\(߼т��~佅9/���x�d���AUվ�������{/���?�,pJ���M�_�I�I�>�[.�����<�HKҾ�|��w���1�6;���W���,L���,H�����'ż�N���5�Lp��۸�Z�ؽY��N��"��l��   �   U/�������� �c�F�#�@&����ػ��<2��<�_=�[=��=��=���<�08����Bǜ����9M�J&��vn¾������j%4�F�L��_��l�&p�`�k�+_��K��43�V��.��7�¾k��w�V������˽5���0�8[��0ͼ��Ѽ����(H�@O?�"g�mZ��-���Tn�����r1��SϺ��   �   ��F�R�(�f��,<���i��@�;�,�<ʳ�<:#=<8=�A=��6=�N=XƟ< v���4'��ഽ�l�'_h��[۾�@��,���J�aUf�0�{��ڄ�{,�������|{�[�e���J�,����2�ݾ\���P6w�M/��T�?�����[�X�����43�<C����
����J5�lI�z\Y��d���i���f�R�[��   �   �5���=r���Ļ��{;9j<`V�<w=�%2=ަM=`Z]=�C]=�I=��=6�<0�t=>�vsȽ�o(�&~�u첾*�*��_Z;��\���z����~��r��km��2눿z���\���;����3�gC��1f��'�B�V[�$)��f<~�8�5��$�d{���{�����������`��z��4<�L��������   �   p�� ��9��<�E�<0o�<��=B)7=0oT=,�i=�Fs=�fm=�S=]� ="��< I ��M�s:ս�-2����"��������� ��'E��Jh��������헿7����藿����؃�)�h��F��w"��p ���þ/����O�ż�v�ǽ�8����F���x�������g��~��@�8F�������$�ļ̚���Q`��   �   `>��`�;�u`<L�<3� =�$=H�D=��_=��r=�z=�r=>W=�n"=�Ɲ< �*���R�[�ٽg�5�0{���쿾�( �Ʃ#�ȇH��;l�����7{���{��w;��K{��愒������l���I�
d%�<��ƩǾ�j��!ZS�q��o̽8����L� ��s�f �T����S��|����?���E�\�Ǽ$祿�3u��t��   �   �� �9��<F�<�o�<�=r)7=foT=d�i=�Fs=Fgm=��S=� =
��<`C ��M�
9ս�,2�B��=��������� ��&E��Ih� �������엿����藿I��*؃�#�h��F�8w"�
p ���þv����O����ǽ�7����F�"��Ɣ�T����d�����>� E������⼈�ļt����O`��   �   `4��0;r���Ļ��{;L:j< W�<Gw=8&2=L�M=�Z]=�D]=�I=F�=�9�<@��9>��pȽ�m(��~��겾�'�����X;��\�s�z�T���}��1
��.l��ꈿ�|z���\��;�K���0�A���d���B��Y��&��8~�t�5�^!�u��|u������� ����j��p:�ģ�n�����   �   ��F�x�(����(;���f����;�-�<���<�#=�8=΢A=Ǝ6=�P=�˟<`W��4/'��ܴ�>j��[h��xX۾?��,�6�J�fRf���{��؄��*������by{�U�e��J��,�����ݾ㏨��2w�!J/�<P񽖳����[���l���H*��:����
�6��vF5�*I��YY�n�d���i�B�f��[��   �   �.��G��������c�ʀ#�`%�� �ػ��<���<�`=�\=�=�=`��<��7�������H5M��#���j¾Y���*��@"4���L�4�_��l��p�F�k�B_�V�K��13����� ��|�¾h���V�!���˽�0����0��N���sͼȮѼ����ZC��J?��g�}X��z����l�����x0���κ��   �   �T�E���&��Խ֝��h_{��� �D&�� �A�@�k<f��<*W�<�X�<��< �/�߼̂��w��4/���x����bPվ���G���w/���?��kJ��M���I��>�v�-�*���9�MFҾ�x���w���1��3��zQ��#L��� �(:��d��,ż I�`�5�D	p��뗽�ٸ��ؽ��������l��   �   JX���O�3@�ޝ)�b��ǽ�ֆ��Z�X�4�@������;�y�<Zܗ<�Z< [�9�5���PS�ʘ�����.N��O�������پ� ��W����u'�0.*�ճ&�i��6������mӾ-��\섾�qE�6��ڌ���i�ҵ	��@ik�l(��5ǼJ��ba���jʽU���o��p�-�&�A�\UP��X��   �   jE��f���ފ���x���U���.���@>½�M}������Q�@��:�|<��< bԹ���Hd'�O��x:齀'&��^��G���:��� ;���V���N��������������ž�ϥ��1���^L����ҽ˽-ǀ����P?������\ ��Fg��Uݼ,�;�3T����ɽ��`)��L��n��8��������   �   Zо)�ʾ�|���
��35��7�w��uD����{HϽl-��a�p0����u� �9��J�@|h��A���l���������.�-^�`�������������þ��;��Ͼj�ʾ y��V��<2���w�OqD�}��BϽ�(��*Z�0&����u� 4�9��J��|h�|C�J�l��·����X�.��0^�����f������j�þ��;�   �   ������������Z�ž�ҥ�`4���bL������˽�ʀ�����G��P��c ��Hg��Sݼ��;�R��R�ɽ���i)�b�L���n�.6���|�����=B��=���ۊ�1�x���U���.�W��8½�C}�����Q��k�:��< �< Թ��tf'�P!���=��)&�*�^��I��c=���#;��2���_���   �   p0*��&�Ek��8�4����pӾ�/��s�tE�ǚ�ː����i�F�	�`���Pqk�@*���4Ǽ���Ba�G�ʽ����w����-���A��PP��X�$X���O�E�?�J�)�A����ὰ����X����@������;"��<P�<x�Z< q�9�7��tSS�������1N�;Q������s"پH
 �`Y������'��   �   V�M�+�I�4�>�t�-����o;��HҾ�z��
w�0�1�t7��sT���'L�(� ��>������ż4H�H�5��p�'闽2ָ���ؽ:��o�� �;h��P�F������ԽP����S{��� ���� @;�P�k<���<]�<�\�<n�< �/��߼͂�Dz佴6/��x�/����Rվ������y/���?��mJ��   �   p�X�k�B	_�0�K�N33��� ��x�¾�i��Q�V������˽�2���0� S���vͼ0�Ѽl���B�ZH?�g��U��)����h��� ��#+���Ⱥ��(��J�����c��v#���� �ػ �<���<�d=`=Z�=R�=���<��7����Ĝ����6M��$��kl¾\���h���#4�i�L��_��l��   �   �+��ض��{{���e�W�J�,������ݾ:����4w��K/��R�i�����[���4����+� ;���
�Ƒ�D5��I�UY�Ҥd��i���f��[�L�F��(�����+���-���H�;�8�<޽�<�'=�8=�A=h�6=�Q=X̟<�Z��f0'��ݴ�"k��\h��𣾿Y۾�?��,�p�J��Sf���{��ل��   �   �
���l���ꈿ~z���\���;���2�B���e��=�B��Z��'��&:~��5�r"�|v��v�����*������������6����Ē�؅��)���%r�@cĻ`�{;�Lj<"_�<�z=0)2=©M=�\]=F]=�I=��=J:�<8�Z:>�|qȽ�n(��~�i벾�(�_��pY;���\�q�z����Q~���   �   ⟚�W藿���}؃���h�rF��w"�lp ���þ헐�~O�u���ǽv8����F����@�������d��Ĭ�0>� D� ��h����ļ$���`F`� �� K�9��<�J�<�s�<�=,+7=�pT=��i=�Gs=hm=.�S=p� =���<8C �0�M�@9ս�,2�n��������'� �0'E� Jh�^������D헿�   �   Pp^��jZ�h�N���<�Y$&����9��x#����T�}'� ��z��X������ƅ��	���ϔ�7Ɩ�թ���[���ր�&�_��H7��
�`���R0� �/:p�A<�5�<��=8*.=D�Q=$\p=�P�=���=���= v�=.F�=�X=yb=xAf<H���$en��b���3�ج��뼯�n��q��)�%�l�<�J�N��kZ��   �   �Z��V�z4K�w9��2#�}
�*��ȳ��d����P�̭��뽃���AK���΍��늽h����!���˔�M����D��M遽xjd�Vb>������ͼ�d���2��<���<���<�F!=F=0f= �=�Έ=��=@$�=�;=P�V=�=`fi<�4���*i�g"޽�o0���~�ķ���޾�V	�R�"��L9�84K���V��   �   e�O�S�K�\�@�7�/����"�J�־	ͩ��l����C����ڽ�����َ�3���Ġ��$�������V��[����������D[s�
�T��+1��!
�̏��x�W�@U �0�	<pϝ<�-�<��"=@�F=0�d=9{=���=`�=�t= 'P=��=`�p<ؽp�nZ�N�ѽ�O'��q�����mӾ�k�:z�-�/��@���K��   �   �B>��:���0�r� �W��X�]yþ(>����k�I0����t���n����v�fb�n b��,n�Z�ۇ��������������ч�o}�@fe��8H�&j&�`] �ʬ��8$����:x\<NH�<��=j�7=hPU=�ih=�m=B�b=D=p&=�&v<��G�ԵD�@����c��^�����!¾�iﾀ��o!�\�0���:��   �   C[(�/%�R��~������ VҾ]?�������ZL�	����ڽ
���Yp��E�H�6���;��"N��f�Q���	c��~���W웽Tힽō��=�����A?����n��!G����4�ż��)�� l;.��<���<Y�=4�;=��J=@�G=61==�=�=r<����+�`����X�^�E���w��K�Ծ�w������G�%��   �   4��m������G��Ӿ�����􏾇s`���(��i�������r�0)0�J]����BC�μ-�2�P���w��Џ������������n�̽�VӽD~Խ�dϽ�zý����9[���q��8-���˼ �� <���<=#==B#=�M=H��<�!\<Ps����7�<� +��Mg�ۓ������W�׾G6���-��x��   �   ���I�!�پ�8žܫ�䏾�8g�"�1���������w�z�!��EڼM�����ټ�m���A���x�N���丽�׽p��G9��������f���\�
�b����Խ�[���iz��b �,����9N�(R\<�%�<���<�s�<�Z�<��+< ����ƍ{��5ɽA����B�& y�Xk���^���<˾��ݾ�p��   �   #ܻ��鶾�z��v���tڅ�^��/�5g���>�x�v��$4����.����hz,�\���,�����<�H�ŭ��ڽ�Y����/��sA�{�M���S�A�R�ڱI��9�E#�����׽���hFO�@0߼�L�PS�;��j<+�<x<h<Д�;���\��6Z��ժ�V�^!���K�W�w��ϐ�l2���^���蹾�   �   �����銾�W���Cg��E��n!�+�����Z�l�����k�`B�p�; ��;�5��J��o开�D�C`���2˽WA�.�$�6E�D�c�̌~�D���쎾>���n슾\Z���Hg�>�E�'r!�&1��"�����l�̮��
l���� ̆;�o�; u���
J�(p�T�D��^��X0˽�?�Ɵ$�	3E���c�p�~��A��Jꎾ�   �   ɩR�k�I��{9� A#� ����׽M
���=O��!߼�4��y�; �j<1�<hEh< ��;p�����(8Z�zת�Y� !���K��w�Ґ��4��}a���빾!߻��춾�}������܅�^�i�/��i�X���l�x�N���=����.�p���`�,�蹖�����F�<�q탽2ĭ�h�ڽ�W�����/��oA�r�M�U�S��   �   q����
�h��2�Խ�U��6_z��Y �<��� �L��f\< .�<��<�x�<H^�<p�+<0뻼�����{��7ɽ���P�B�Py�Rm��a��J?˾��ݾ�s�Ҹ�2L��پ�;ž�ޫ�!揾<g���1�� �X����w�v�!�,Nڼ�S�����|ټjo��A��x��L���⸽�׽�}��6������fc��   �   �tý����U���|q�X/-��˼8b ��� <� �<+=~@=�#=�O=���<H#\<@x��`��Ò��>��+�BPg�����������׾9��/�z�Ѿ���<��:J�fӾ����~���Qv`�ć(�Lm�������r�F-0��`�����E���-�P�P��w� Џ��������������̽pRӽNyԽf_Ͻ�   �   X�n�\G����\�ż�e)� �l;nȊ<r��<J�=p�;=4�J=0�G=�1=�=�=r<�����+����?Z�0�E��Uy��=�Ծ:z�������Ą%��\(��%������������WҾ�@��􃆾�\L����o�ڽ<��D]p�^�E�8�6�n�;��$N���f������b��Э��뛽_랽3������풽5;���   �   bW �콬�� $��o�:X'\<�Q�<��=�7=PSU=�kh=��m=��b=�D=�&=�%v<�G�̷D�ֱ���d�G^������¾=k�}��&p!���0���:�%D>��:���0��� �X�UZﾦzþ3?���k��0�0��cv��Lp����v�� b��b��.n�|[��ۇ���:���摍�SЇ��k}��ae��3H�zd&��   �   �W�  ��
<�֝<�4�<��"=��F=p�d=�:{=N��=��=��t=�'P=��=�p<��p��oZ�� ҽ�P'�f�q�����nӾ�l��z��/���@���K�Q�O�6�K�0�@���/�L���"�0�־�ͩ�pm����C�@��H�ڽ����ڎ��������ᧄ�����LW���������������Ys��T�()1�B
������   �   @�2��"<�<.��<�H!=�F=�f=<�=-ψ=p��=�$�=�;=p�V=�=�di<�5���+i�F#޽2p0���~�H�����޾4W	���"�M9��4K��V�d�Z�~�V��4K�lw9��2#�E}
����jȳ��d���P�%��>�����K��@ύ�슽����V"���˔�b����D��遽�id�<a>�4��0�ͼp�c��   �   ��/:ЪA<�5�<��=@*.=D�Q=(\p=�P�=���=�=v�="F�=��X=4b=X@f<����en�,c�2�3����������⾄��<�%�|�<�T�N��kZ�Rp^��jZ�_�N���<�J$&� ����8��`#����T�c'�����y��T������ͅ�����ϔ�4Ɩ�ʩ���[���ր���_��H7��
����Q0��   �   ��2��$<���<���<�H!=�F=�f=p�=Bψ=���=�$�=><=��V=��=@ii<�2���)i��!޽:o0�c�~�v�����޾�V	��"�EL9��3K��V�n�Z���V��3K��v9�22#��|
���⾊ǳ�d���P�>���뽴����J��΍��ꊽ����2!���ʔ�P����C��"聽�gd��_>����0�ͼ@�c��   �   (�W�� ��
<�ם<l5�<�"=@�F=��d=R;{=���=8�=��t=�(P=l�=8�p<�p��kZ���ѽ�N'���q����lӾfk��y�p�/�A�@���K�{�O�g�K�w�@�_�/���k!�$�־̩�l����C����f}ڽ����b؎�倂�s�������q���-U��v�������צ��xVs��T��&1�Z
�X����   �   �U �@����$����:�)\<�R�<�=d�7=�SU=�lh=��m=��b=^D=�(=�1v<��G�"�D����Lb��^�l����¾�gﾒ���m!�5�0�Q�:��A>���:�H�0�M� �V��V��wþ�<����k��0�Ʊ�Zr���l���v��b���a��(n�lU��؇�狍�����k���·��g}��^e��0H�Zb&��   �   V�n��G�l����ż�b)�`�l;xɊ<���<��=4�;=�J=v�G=^ 1=w�=�Kr<�p���+�u���+W�(�E�'텾v��X�Ծ�u��_����́%��Y(��
%����%��)����SҾ�=��6���{XL�����ڽ[���Tp���E���6��;�~N�R�f����{_������蛽�螽爞�"����뒽�9���   �   �sý5���U���{q��.-���˼�_ �0� <2�<	=�A=G#=�Q=@��<3\<�L���	�;���7콜�*��Jg����������׾z3���+�Lw����̺�.���D�fӾL�����_p`��(�e��#����r��#0�$X�|���=���-�d�P�D�w�B̏�����~�����U�̽\Pӽ�wԽ^Ͻ�   �   ��U�
������ԽRU���^z�\Y ����� �L��i\<>0�<���<�|�<�c�<��+<p��l���B�{�1ɽ�����B�R�x�i��/\���9˾��ݾ�m�J���E� �پ�5ž|٫��᏾�4g���1����X��ƀw�D�!��:ڼ�A��� ����ؼ0g��xA�&�x�,I��&߸��׽�z�5�������b��   �   L�R��I�e{9��@#�����׽�	���<O�l ߼�1�Ё�;Жj<5�<�Ph<���;����x�<.Z��Ъ��P�$!��K���w�c͐��/���[���幾�ػ��涾�w������ ؅��^�t�/�'d��ڊx�b���'�� �.����c,���������r�<��都������ڽRV�:�U�/��nA���M���S��   �   b����銾�W���Cg���E�on!��*��ж����l�b��@�k� -����;p��; ¾��I�Lb�Z�D�?Z���*˽v<�.�$��.E���c�i�~��>��{玾����犾2U��?g���E��j!�|$�������l�J��8�k�@����;��;�{����I�da��D�^[��-˽>�\�$��1E�z�c���~�NA��ꎾ�   �   �ۻ��鶾�z��b���bڅ��^���/�g��󻽎�x�����1����.�0����m,����� ���|�<�都"�����ڽ�T���n�/��kA���M�s�S�ޤR���I�w9��<#�J��#�׽}���3O�߼��p��;�j<p;�<8Zh<�̶;���@y缾/Z�|Ҫ�,S�!���K�E�w�lϐ�2��r^���蹾�   �   }���H��پ�8žܫ�䏾~8g��1�n��Z��F�w���!�LCڼ@I�������ؼ�h��yA���x�VH��{ݸ��׽(w�Z3�P�����P_�V����
�����ԽNO���Sz�"P �d�����J��~\<�8�<��<ց�<�g�< �+< �����b�{��2ɽ
����B�(�x��j��c^��N<˾s�ݾ�p��   �   *��d�����uG��Ӿ������ns`�n�(�vi��S���&r�.(0��[����F@���-���P���w��ˏ�����}��{�����̽=Lӽ�rԽ�XϽUný�����O��Pqq�%-���˼B �`� <��<T=E=#=�S=��<�5\<�M������ :�* +��Lg�x���Y����׾6��l-��x��   �   >[(�+%�P��|�������UҾT?�������ZL������ڽ����Xp���E���6���;��N���f�����}_������曽瞽����.���蒽6���n�dG� ��Ķż�E)���l;�Ԋ<f��<��=�<=ԓJ=��G=�!1=y�=`Mr<0r��+�����(X���E�0ww���Ծ�w������?�%��   �   �B>�ު:���0�r� �W��X�Vyþ#>����k�60���at��rn�� �v�<b���a��*n��V�ه����Z���ώ��͇��d}��Ze�(,H��\&��O �p���$��=�:�>\<0\�<D�=�7=�VU=�nh=��m=.�b=xD=|)=H2v<@�G�>�D�
��� c�#^�H����¾di�q���n!�V�0���:��   �   e�O�S�K�[�@�6�/����"�G�־ͩ��l����C�t���~ڽ΋��pَ�Ձ��E���m�������U��������������fUs�N�T�r$1�n
��~��ȏW�����
<ߝ<2<�<�"=��F=$�d=@={=Q��=��=��t=V)P=��=��p<�p�XlZ���ѽ8O'���q�����mӾ�k�2z�&�/��@���K��   �   �Z��V�y4K�w9��2#�}
�)��ȳ��d����P�ƭ���j���K���΍�Y늽����!��˔�x����C��聽�gd�_>������ͼ`�c�@�2��+< ��<N��<bJ!=PF=f=��=�ψ=�=�$�=�<=b�V=��=�ii<�2���)i�"޽mo0���~������޾�V	�N�"��L9�64K���V��   �   �������
�k���{޾�������Oaz���F�:��(��{.彾 ٽc�ܽ�(�z��������� v������a����2ӽ�h��S;����3�@ɼ�NԻ��#<�:�<(9=�I=��p=��=���=�=�Ν=��=p�=X:�=0TO=�P=��<4c��(�p��׽�#�;sc������,���ܾUj��v�
����   �   ��$G�b����>bھs��б���_u���B��'�~{���߽d�ӽh\׽���� ���������D��Y�����tҽ����������8�ԯּ��
��^�;4D�<`�=�@=�7h=(2�=NK�=, �=�B�=X�= �=P�= M=��=��<�-��:�l�j�ӽu� ���_�1I����	�ؾ����a��P��   �   �_���(�|-뾨ξZ'������n�f�Jy6�������n3Ͻ�ý�ǽĵս/��x���<*����V�L� �LH콅sϽ`���zu���I�R� ��Up����:pP|<Р�<v�$=.eN=.q=��=N�=��=NX�=���=�`v=�F=��=��<��1b�ʽ�u��(U�q3�����pξ�r�ab�����   �   X���|�����Hp־�������?d��g"P��#��� �$nѽ�w��PJ���7��Aڼ�D�Ͻ���[�x��,/�����b��$	ͽ�����6��g��n'��Ҽ�]3� �J;��<�n�<�_"=lKI=P�h=�=�M�=��=�Ԁ=�f=49=���<Ht<l���JXS��	��PN�sE�;_��EB���=��n�׾��8����   �   ?��Lܾ7iϾ�9��|���bȊ��Gb�D<3��R��ؽHV��'t���������`w�����x�ýi/ս�nὨ���� (ܽZ�ͽ]���)L��ǻ���Yc�F=-�L���w�@����V@<l��<5'=<c6=,�S=$af=��l=��d=��M=�2%=\��<��;�]��?D�:����6�1��1f�0��c��\�����Ѿ�uݾ�   �   �����溾���gў��A����g��G;��o��}߽�w��j���<Q]�րO�`Y�
�t�RX���J���2��Ȱƽ�7ҽ 5ؽ2�ؽ��Խf̮̽���ܯ�Dɜ�������Z���#���Ѽhs3��@];$��<6]�<s�=T�3=4m@=�+>=��+=ϸ=�"�<��T;����\g9��@���署5��I�&Cw�����Ԥ�'۳�)���   �   .Z��>Ҙ��Ꮎ�{���^�E+8���h
�Q���Jo��R0�lR�P��4��j�,�D�T��E������&���`���IѽB!ݽ��x�软T�(����׽:�ƽf���8���h�D�#������4ڻ�_ <���<���<�=�=b =j|�<ȵQ<`b#������ 7��T���Dн�&
��2.���R�.Uu�gǉ�yQ������   �   �ky�,Mp���^��SF��)�A�	�0սw�����V�&���n���v�`�d� ې���ϼ�T��F��~���������ҽ��!� ���	�:D�p6����h�� ��3罶;ý �����`�
���\�� ���x�#<��<ң<%�<�BK<@';pi2����2�@�i���v����������1�� K���`���p�@�y��   �   o�>�� 5�jj%��F�� ���L����7� �Ҽ�4��֫� B[;�+K;@�պ��'����^��n�X��ɐ��(����޽�a����&�ڪ4���=�܈A��>�i$5��m%������B��4Q��`�7�H�Ҽ��4�@y��`�Z; �J;@Yֺ0(�$����F�X�?ʐ�3(����޽ ������&�2�4���=���A��   �   �e����-�<6ý������`�0��HO���̻�$<�!�<:ڣ<d,�<�OK<@6';X_2�l��R�@�����w������2��1��#K��`�Cq��y��oy�(Qp���^�(WF��)��	�$ս�����V�D���y����v��d��㐼�ϼ�X���F���~�~	��8��=�ҽ����� ���	�B��3����   �   ��ƽ����3���}h��#�������ٻw <�ˡ<���<��== e =ځ�<��Q< G#������ 7�HU��Fн(
��4.��R�Xu�$ɉ�lS����V\��bԘ��㎾�}��J^�6.8�����ུT���Po�tX0��W�*�������,���T��G��p���w���,���"Iѽ� ݽN���zQ�C�⽊�׽�   �   X���\�Z��#��Ѽ�X3���];��<�f�<��=��3=^p@=x.>=\�+=غ=�%�<��T;t���h9��A�����7���I��Ew������֤�(ݳ�L��.����躾���JӞ��C����g��I;��q�<�߽�z����6V]���O��dY���t��Z��M���4��b�ƽ9ҽ�5ؽ�ؽ#�Խ�̽�����ٯ��Ŝ��   �   �7-����v����Xk@<��<i+=�f6=p�S=�cf= �l=�d=t�M=W4%=r��<��;T^��R@D�p������1��3f�A1���d�����v�Ѿ�wݾM��R ܾ!kϾt;��
����Ɋ��Ib�&>3��T�ۈؽ�X��pv��񿋽����y�������ý\1ս@p�������m(ܽ�ͽl����J��¹��Uc��   �   dҼ�M3��$K;���<Xv�<c"=�NI=��h=h�=�N�=l�=rՀ=f=59=���<�t<�����YS���;O��E�`��[C��?����׾��������/�����뾾q־�������*e���#P�A�#�� �&pѽ�y��(L��z9��ܼ�*�Ͻr���\�0z��j0��f�����	ͽ����5��Rg�~k'��   �   Lp��݀:[|< ��<��$=lgN=@q=���=�=���=�X�=��=�av=TF=�=�<�\2b�ʽwv��)U�4�����mξ t��b����&`����(��.뾒�ξ#(��x�����f�2z6�t�����4ϽU�ýn�ǽ&�ս�������*�H���V��� ��H콒sϽ����t��� I�0� ��   �   ��
�i�;�F�<��=Z�@=�8h=�2�=�K�=� �=HC�=��=S �=��=HM=��=��<�.�� �l��ӽ�� �@�_��I�������ؾg���a��P�	�vG�Xb������bھjs�����v`u�0�B�#(�4|����߽�ӽ(]׽��彬��V���G��������,��xҽi���Z�����8���ּ�   �   �LԻ��#<�:�<C9=�I=�p=��=���=�=�Ν=��=g�=S:�=TO=�P=��<�c����p�$׽�#�ksc�ֿ���,���ܾpj����
����������
�Y��p{޾|������/az���F�*��#��v.�� ٽp�ܽ�(뽐���������!v����
��L���d2ӽhh��3;��d�3��ɼ�   �   ��
�0o�;H�<'�=��@=9h=�2�=�K�=� �=gC�=��=} �=�=�M=m =`�<�+���l���ӽ	� ��_��H�������ؾB��Oa�UP�c��F��a�s���aھ�r��Z���0_u��B�9'��z��.�߽��ӽ�[׽�� �����n�����������.ҽQ���f����8� �ּ�   �   �Dp���:h_|<Χ�<��$=�gN=�q=&�=B�=ڇ�=Y�=Y��=�bv=pF=��=��<잼\.b�jʽ�t��'U��2������ ξ�q��a�=���^�:��b'�M,뾖~ξl&������f�,x6��������1Ͻ��ý��ǽB�ս��轵���H)�����T�(� ��E�qϽ����s����H�Կ ��   �   <Ҽ�E3��<K;8��<*x�<�c"=OI=��h=��=O�=��=�Հ=4f=�69=��<Ȁ<@���TS�g���L��E�7^��A��Z<����׾D�w�����������d�뾯n־1���e��&c��� P�j�#��� ��kѽ�u��EH���5��ؼ��Ͻ��ZX�u��,��D���㽶ͽ(���3��H
g�8h'��   �   �4-�X����v��߾��o@<���<",=�g6=�S=�df=�l=�d=ܑM=A6%=���<�5�;TT���9D�����1�/f��.��oa��������Ѿ�sݾ��,ܾ0gϾ�7��ɑ���Ɗ��Db�:3�Q��ؽ�S���q��D���F����t�����U�ý�+ս�j��������#ܽ��ͽ񔺽�G��[���$Qc��   �   ������Z��#� �Ѽ�S3���];���<Th�<N�=��3=Jq@=�/>=��+=�=�+�< �T;t����`9��<�����,3��I��?w�&����Ҥ��س��������\亾ؗ��^Ϟ�@����g��D;�Om��y߽�t��_����K]�X{O�^ZY��t�U��`G���.����ƽd3ҽQ0ؽ&�ؽ��Խ
̽V���Rׯ��Ü��   �   ڵƽ@���2��^|h���#�К��P�ٻz <͡<b��<��=I=�f =F��<�Q<�#�@���P7�_P���?н$
��/.��R�MQu�Lŉ�9O������W���Ϙ��ߎ��y��:^�(8�R����M��rCo��L0�xL�~��2���,�R�T��A��}�������l����Cѽ�ݽ��:��@N轢��l�׽�   �   �d�� -罆5ýp�����`�n���M������ $<�#�<�ܣ<l/�<xXK<�e';@O2�����@�⩍��p��N�����w�1�"K���`�U�p���y�:gy��Hp���^��OF�9)�(�	��ս������V�.��Lb��@�v��d��ΐ���ϼ~M�>�F�d�~�������
�ҽѭ��� ��	��@��2����   �   ��>�X 5�j%�u��̦�
��lL���7�зҼ8�4� ���`S[;`BK;��պ��'�8��\��ҺX��Ő�#��И޽� �V��%�&�O�4���=�U�A�F�>��5��f%�2��֠�o���G���7�$�Ҽ��4� ����[;��K;�պP�'���������X�Ő�)#��ř޽�����)�&�Ӧ4�t�=���A��   �   -ky��Lp���^�XSF��)��	��ս+�����V�z��Tm���v�p�d��א�ئϼXQ���F�>�~����"����ҽ����� �x�	��>�P0���a�!�0'��/ýU�����`�P���?�� ���&$<�,�<��<�6�<�eK< �';�D2�t����@�ҩ���q��������N�1��K���`���p���y��   �   �Y��Ҙ��Ꮎ�{���^� +8����&
��P���Io�>R0��Q�N�����p�,���T��C��D�������V����Cѽݽ����HK����6�׽@�ƽ|	��>.��Bsh�D�#������ٻ�� <bס<>��<��=�=�i =ȋ�<x�Q<��"������7��P���@н%
�p1.�'�R�Tu��Ɖ�Q������   �   Ӌ���溾����Vў��A����g�hG;��o�|}߽�w��%����P]��O��^Y�x�t�AW��zI���0��6�ƽ�4ҽ1ؽ@�ؽ�Խ� ̽H����ԯ�����5���`�Z���#�ķѼ�83� ^;���<�q�<��=`�3=|t@=p2>=l�+=0�=>/�<��T;����`9��=����V4�͵I�Bw�����iԤ��ڳ�����   �   "��6ܾ)iϾ�9��q���XȊ�sGb�,<3��R��ؽV���s��m���c���v�����`�ý�-ս�l�*�����V$ܽޛͽ9���iF�������Lc��/-�x����v�@1�� �@<��<X0=Tk6=P�S=�gf=p�l=H�d=��M=�7%=Z��<�<�;�S��$:D������.�1��0f��/���b�����\�Ѿ�uݾ�   �   F���m�����@p־�������6d��V"P�ބ#��� ��mѽ�w��J��R7���ټ���Ͻӯ�Z�:w��_-��D������ͽ����\2��g�Ve'�|
Ҽ�63� {K;��<t�<Dg"=4RI=H�h=T�=P�=��=�ր=�f=�79=���<��<,����TS�#���M��E��^���A��{=��@�׾������   �   ~_�޳� (�x-뾣ξV'������d�f�Ay6����~��N3Ͻ��ý޷ǽ��սγ������)�?��vU��� ��F�oqϽ�����r����H�(� ��<p�@U�:i|<���<��$= jN=�q=�= �=���=�Y�=ܔ�=hcv=.F= �=��<잼�.b��ʽ5u�F(U�>3����Mξ�r�Wb�����   �   ��#G�b����;bھ
s��ϱ���_u���B��'�q{���߽P�ӽL\׽��彶 ����Y������������nҽb���Y�����8�ԩּH�
��w�;VJ�<H�=Ȍ@=*:h=E3�=LL�=!�=�C�=�=� �=~�=LM=� =X�<T+���l��ӽ4� �`�_�I�������ؾ����a��P��   �   R���F������������`Js�j�L��Y+�ޑ����je��ʣ�\.��(���@���X��m�k�z�(����z��Hl��U�M�8��q�xF���&�Y��LҼ hȺHW�<�=ԩP=|5=�=�=Ǔ�=jߤ=�R�=ڤ=�	�=�I�=��u=$�==z��<�8�;����XZ�=���Q��'7��pg�d�������~��O���   �   �G�������s��%���2��cn�|;H���'��2�p� ��A��s|����J%�&�<�|T��{h�;v���z�']v�(ch�`R��Y6����d6��=��ȆZ���׼ I(���<�S=�J=�Ty=�k�=�=�j�=I�=9��=`��=�'�=8�q=�/:=�q�<�p�;lի�.�X��!�������4���c��ۈ�G���m��nŷ��   �   XN��W���0ࣾ���,'��g'`�o�;���Ac�Q�i_�V����A��"A1���G�t[��[h���m���i�G5]��I��!/�������k���W^�l��`˿� e<NO�<��8=�yg=�=��=��=���=Nݛ=2?�=e��=�e=z�.=V��<p��;���ޚU��Ჽ{��n+-���Y��e��+��������.���   �   K衾�F������>��:m�~�I�K(������oeҽ�B˽�ս�7�Z�	�\��@!4�CjF��TS�nY�ǝV�'@L���:��|$���
�n�޽u�����g�D��)B�P�;���<c?=��H=�n=C�=J�=�Ǒ=��=�Ɉ=D�v=PTO=jM=���< 	�:a���IS�y���̘��j6"��xJ�%q�ଉ���k���   �   ���������K���k�QtM�'�-��v��3�N�Ľ���0�������ǽ[�R��bQ��,��&9�ՠ?��?���7�]*��P��(���ؽ�����={��%&�4q����q�8BG<�Q�<L=d�D=z�b=�w=�"�=8%~=`%p=�U=z	/=�!�<pm< m���Xڼ��U�����>���?8�KY�z?v��J������   �   ��r�\�j�>�Z�}JD���)����p��-7��{Y���C��V�{��f��:��޳���~۽&0�����<[���#�,�%�L6"�������"�����׽�����ԾU���ė�� �Z�/2<^��<�8=�}.=��E=8�Q=��P=*�C=�k)=N�=���<���;�DQ��a�lhb��ͣ�*(ڽ�a	���%�@�t�V��h��q��   �   ��G��0?��0����Ι���ؽ[O��$q����N�,�,���#��+3���W�4������Iƽ������@��������
������>8߽��Žor���H��J�]�\D��z���J��H�; z�<�f�<)�=v]=�X=h=�<���<���;��	� Oʼ�n.��N}��d����ӽT|�����g(�(�8�W�C��TI��   �   :X�����p����� ���j�a���%޼,&���p��p���<���`)��@b�u����ͭ��Ƚ�[߽2����f����������D{���NҽV⻽󶡽R(����H�nj��X���т����;p~<U�<� �<Xc�<�63< �:(7���ϼ�&�D�g�F������Tֽ���g�lx����#���#��   �   �D��v��@
Ľ�|���|��:5��漸Kq��i���\:��;�	��h5	��i��
��ܤ<��4y�����k���ͽ����i.�����L_��M��H����ྲྀĽ8����|��A5�H���cq�@��� �Z:`�;����HK	�4u����Ъ<��:y�G��n����ͽ�P���.�>�����]��K��   �   �޻�A����$��L�H��c��K��Т��0"�;`!~<�^�<@
�<�l�<�I3<@��:@7��}ϼ:�&��g����|����ֽk����g��y�I��#�D�#��Z����` �4��T�� �����a����1޼t1���{��Ж��(���Pf)�vGb�ڼ��5ѭ�@�Ƚ�^߽��n���X�����������y�@��Bҽ�   �   0F��p�]�J>��n���3��s�;���<p�<~�=�a=�\=l=0�<���<���;(�	��Gʼ�k.��L}�:d���ӽ�}������h(��8���C�}WI�^�G��3?�30�v��!���ؽS��yt���N���,�l�#��13���W�]7�������MƽZ�l�����0�����
�������U7߽B�Ž2p���   �   ��U����\��� mZ�hA2<��<�<=��.=6�E=��Q=��P=f�C=�n)=�=���<��;�:Q�`�vgb��ͣ��(ڽub	���%��@���V�h���q���r�#�j���Z�MD��)������j:��y\���F���{��i��K��,���h�۽�3�����]���#���%��7"����P������~�׽���
��   �   �"&��j����q��PG<�X�<rO=��D=rc=�w=R$�=�'~=�'p=��U=�/=*&�<�
m<�_��Wڼn�U�E�$��*��-A8��LY��Av��K�����񫎾H�#M��f�k�pvM��-�mx��6���Ľ�����2��������ǽp����&S���,��(9���?� ?���7�^*��Q�)��ؽD����;{��   �   �~�` B����;��<�A=R�H=\�n=D�=Q�=�ȑ=� �=�ʈ=�v=VO=�N=4��< &�:X`���IS��������M7"��yJ��&q�ʭ����4l��n顾H������?���;m��I�sL(�����뽈gҽE˽�ս:ｩ�	�����"4��kF�.VS��	Y�&�V�WAL���:��}$��
���޽H�����g��   �   @��𿿻`e<�R�<N�8=L{g=��=~�=P�=0��=�ݛ=�?�=���=�e=d�.=���<���;���p�U��ⲽ���(,-���Y�Pf��ۇ��Q���h/��,O��'����ࣾ����'���(`�f�;�ͨ�d����`������8��0B1��G��[�]h���m���i�)6]�tI�a"/������W���RV^��   �   ��׼�<(�t�<�T=кJ=pUy=Zl�=a�=�j�=��=���=���=+(�=��q=�/:=jr�<0q�;�ի���X�`"�� ��6�4���c��ۈ��G��en���ŷ�H������s����3���cn��;H��'�03�ڲ ��B���|�T���J%���<��|T�M|h��v���z��]v��ch�Z`R��Y6�Ʃ�|6��=��T�Z��   �   LҼ@aȺ�W�<�=�P=�5=�=�=ԓ�=lߤ=S�=ڤ=�	�=�I�=��u=
�==4��<�6�;(����Z�q��R��'7��pg�u�������~��V��T���D������������JJs�X�L��Y+�ڑ����}e��ڣ�o.�"�(���@���X��m�x�z�-���z��Hl���U�6�8�iq�HF��ЖY��   �   ��׼ +(� �<TU=F�J=�Uy=�l�=�=k�=��=���=���=T(�=�q=�0:=t�< z�;�ҫ�ȽX�"!��6��>�4�]�c�7ۈ��F���m���ķ�$G��4���s��� ��b2��Mbn��:H��'�P2�	� �A��|�p���I%���<��{T�{h��v�1�z�k\v�fbh�?_R��X6���5뽮<����Z��   �   ���@����"e< U�<4�8=|g=�=��=��=^��="ޛ=
@�=H��=�e=��.=��<�щ;�����U�(ಽ|��M*-���Y�e��d��������-��tM��r���Rߣ���p&��&`�I�;���bb����]�Ӗ����_��)@1���G�B[��Zh�2�m���i��3]�XI�� /�S��N��-����R^��   �   �z��B����;p��<2C=H�H=�n=oD�=��=&ɑ=!�=�ʈ=��v=8WO=�P=���<���:xX���DS�����ԕ���4"��vJ�#q�ƫ������i��硾�E��e ���=��8m���I��I(������4cҽ�@˽��սb5��	�����4��hF��RS��Y�̛V�,>L���:��z$���
���޽B�����g��   �   n&��c�� {q�xXG<�[�<�P=~�D=4c=`w=�$�=�(~=�(p=��U=X/=*�<Xm<�C���Mڼ<�U�P&�����=8��HY��<v�LI�������}vJ��m}k��qM��-��t��0�`�ĽL���c-��c�����ǽ<齜��{O��},��$9�}�?�?�-�7��Z*��N�_&���ؽ����,6{��   �   �U�������`JZ�H2<���<�==��.=�E=\�Q=��P=h�C=p)=*=`��<P&�;�*Q��Z��`b�xɣ��#ڽ"_	��%�#@�[�V�bh���q�f�r��j�,�Z��GD�!�)�N��Z�潒3��AV���@��|�{��c��
��i���{۽�+��g���X�&�#�t�%��3"�������}����׽*�����   �   �C����]�N;�dj���,�~�; ��<�q�<=�=Vb=�]=m=��<�<��;8�	��?ʼLf.��E}��_��l�ӽ�v������c(��8���C��QI�<�G��-?�a0�	��.��4�ؽ+K��km�� �N�ڟ,���#��%3�زW�k0��|���Eƽ�彗���y���~����
���#���l2߽G�Ž�l���   �   }ܻ�e���%#��6�H��a�TI������0)�;p$~<`�<��<�n�<�N3<��:��6��wϼ\�&���g�L��N����ֽ ���d�6u�X���#���#��T�ߛ�������	������<�a�����޼���Xd���~�� v���X)��8b�����ȭ���Ƚ*V߽R����*�������J����t�q��4ҽ�   �   vB�����	Ľ|����|��95�@�漘Hq��c���2\: ;�윺1	��f����8�<�>1y�@���h��/�ͽ>�D����*���~�nZ��H�T>��h�མĽ�w����|�25����00q� 7����]:@U;@J��	�\��p��r�<�~+y����Tf��B�ͽ���ɕ��&+�������[�mJ��   �   NW�d��V����P��������a�X���#޼�$��(o��ĉ��T����^)�&?b�S���Ṋ���ȽY߽�	����T���ި������~s�@��X�ѽ*ٻ�ϭ��x���H��Z�l<���k��pT�;h8~<li�<��<�w�<0a3<@��:@�6� nϼ��&���g�������&ֽ9����d�>v�թ��#���#��   �   ��G�H0?�0�������~�ؽO���p��N�N���,��#�<+3���W��3��_�� Iƽb�$���)��Z��6�Ѻ
��K����1߽��Ž�j��,A����]�r5��^��8�0��;쏊<�z�<��=df=�a=�p=z&�<쪔<�,�;pr	�x8ʼ$c.�vC}�,_��p�ӽ�w�����Oe(���8� �C��SI��   �   "�r���j���Z�>JD���)�q��,���6��@Y��rC��ܠ{��f�����w���T~۽p/��:���Z���#��%��4"�������~~����׽r������U�������� Z��Y2<6��<�A=8�.=|�E=��Q=��P=��C=Ls)=`=���<`>�; Q��X�B_b�Eɣ�	$ڽ�_	��%��@�E�V��h�N�q��   �   g��������K���k�+tM��-��v��3��Ľы���/��ع����ǽ� ��Q�m,�W&9�3�?��?���7��[*�bO��&��ؽr����4{�,&�(^���Gq� fG<`b�<�S=��D=c=w=�%�=+~=<+p=$�U=�/=�.�< m< 4���Jڼ��U�pۘ�Ύ��>8�JY��>v�dJ��U���   �   )衾�F������>���9m�f�I�K(�т�\��Keҽ�B˽��ս�7�>�	�5��!4�jF�HTS��Y�3�V�n?L���:��{$�>�
���޽\����g�py��B����;$��<�E=��H=P�n=zE�=��=ʑ=�!�=�ˈ=��v=�XO=IR=���<���:�V��dDS�	�������c5"��wJ�T$q���������j���   �   @N��E���#ࣾ���$'��Y'`�a�;���6c�<�R_�<����,��
A1���G�O[��[h�I�m���i��4]�+I�.!/�̰���n����R^����`����'e<�W�<��8=x}g=��=d�= �=���=�ޛ=�@�=ڧ�=�e=��.=��<P؉;�
����U�Zಽ¾��*-�=�Y�ze������f���{.���   �   �G�������s��"���2�� cn�s;H���'��2�k� ��A��m|����J%��<��{T��{h�"v���z��\v��bh��_R�<Y6�<���5��<����Z�x�׼�%(��<�U=�J=�Vy=�l�=��=ck�=��=榢=�=�(�=��q=01:=4u�<�}�;ҫ���X�)!��M��l�4���c�nۈ�G���m��aŷ��   �   �c�z�^�:�R���@�7�+���T��%���A��J����"S5���[�P����e��鏯������5̾�0о6̾���Ꮾ�rǗ���|�~�G�(�R̽�Or�xǼ`��;�y�<��A=1|=�d�=O��=���=�(�=��=�j�=�L�=�+�=��]=��%=�)�< ��;����90��#��E�ͽ���( #�)=���Q�f�^��   �   ��^��aZ��NN�ަ<��1(������
�.�0� ����\1��W�����d���9���?��9sȾ�h̾�ȾI;�������@���x��D�)����ɽ8�o�d�Ƽ�;��<�L>=�}x=pi�=��=:|�=\ԩ=m!�={��=7J�=��=�W=en=��<`K`;\ט�ZW2����Jl̽
H�M!�NZ:��3N���Z��   �   �R�D	N��!B��
1�^��
����hB��y޽^����	�~�%�h�I���r�𮎾⌢��в�d���f{�����,z���𢾪�����l��I<�T���½��i��{Ƽ`\;
��<�F4=�$m=�V�=4�=�ˠ=:��=�d�=t4�=b.�=�p=�$C=�=xГ< ���ϱ�2�9�݆���	ɽX} �5��[2��lD��O��   �   �z@��;�BS/�K ��x�<���`׽3OŽc�½��ѽ���x����4�J�Z�q��T~������������������Ky��Q����炾0b[��V/��]�UǸ��>b��˼���:x��<Wk"=�MY=�̀=�*�=�4�=Ob�=�)�=�܈=�Wu=��O=w� =�m�<�U$<������t�H������eŽ|���r�Mu&�(�5���>��   �   ^�)�K�#�����J� �}ͽz���z���랽E���U˽u���|��<�h�_��y���0�����bq��cw��ّ��f����j��:F�& �/���ɮ� ^�hBۼ �N�4��<�$=��;=|�b=�|=�[�=���=n~=Nh=HzH=��=��<��X<����O��D/�"Ld�A嚽UIĽ.�����k���$�*��   �   %e��	�F�����ݽ`��ğ�#e����p���k�캁�*[��	�Ľ�����9��&9�RV�l�n���������"�z��sg���M�<*0�����B�XЧ���a�������"��L<���<:=t�8=��P=p�[=��Y=<zK=�W1=F�=�)�<�!)<@
}�@�����:�N�w��:��Zɽ��潀� ��
�J��*��   �   b���߽V�ƽA������a�R5�n�.��|y(��U��{�������`�da*��@�[�O��X��<Y��PR��D�>�1�������ֽoԦ�"�r�F��L�����T���7<�+�<�4=��=p$=�*=!R=f �<tÂ<�}S;� 5�ּ�?)� �e�t|��l�����U�ֽ���H�������%;�>g���   �   ��ǽX^���O��r�p�,�7��y��_��@ֆ���v� ���(����,��zw��¦��Խ�����0�D!"�%�+��-/���,��{%�����H��u��^Aҽ6<���I��*'N�Zo
����p�����;���< �<���<�~�<`7�<P��;�i˻Ǭ�\����\�����ث���Ľ�mؽ�����p������m�Pw�;�ڽ�   �   tr������6S�@V� }���9�@�	�`Hm;0_�;��;P饻6����J�����/����Խ8�����e
��������1�� ����ؽrt���t��󍇽vS��[�������9� -
�`�l;�5�;�=; ��4��������J��	��l4��pս#�k��	h
��������2�  ����ؽ�r���   �   �H��j#N�k
�����퐻��;��<��<���<���<B�<,�;6˻���������\�檎��ԫ���Ľ�jؽI�����o��Z����m��x�b�ڽ��ǽ;a���R����p��7�V��j��8ᆼ�v�ص������,��w�UǦ��Խ	����3�$"�ޢ+�l0/� �,�~}%�����I�vv��8AҽK;���   �   P�r����������T���7<`3�<�8=y�=}$=�.=�V=T
�<\΂<`�S;X�4���ռ(9)���e��y���ꩽ���7�ֽ���ժ������)<��i��a��N�߽��ƽ�����a�5������(���U�O��������� �@d*��@�h�O��X�p?Y�uSR��D�� 2�8������ֽԦ��   �   ��a� ���@�"��W<���<E=��8=$�P=��[=0�Y=�}K=�[1=��=T3�<�5)<��|���2���N�ou��9���ɽ��� ���
�w�����f�Ƽ	������ݽ�����ǟ��g���p�f�k�޽��i^����Ľ���<<��)9��TV�x�n�������i����z��ug�@�M��+0�����C�sЧ��   �   �^�X@ۼ��N�0�<�&=�;=��b=R|=D]�=���=\~=<Qh=�}H=>�=���< �X<����H��t,�Jd��䚽jIĽ��u��d���$��*���)��#�(��
L��"�5ͽ��<}��V����R˽zx���~�E�<���_�\{��P2�������r���x��Qڑ�h����j�L<F�
 �0��'ʮ��   �   �>b��˼ Ԇ:H��<�l"=lOY=�̀=�+�=�5�=Mc�=�*�=�݈= Zu=0�O=,� =s�<�_$<@�����b�H�����]fŽN����r�;v&�H�5���>�|@�U;��T/���z�����6b׽BQŽ��½��ѽ\�����y�4�.�Z����~������궬���������\z��<����肾Xc[��W/�^��Ǹ��   �   ħi��zƼ�!\;���<�G4=�%m=�W�=�4�=>̠=Ⱒ=�e�=75�=-/�=��p=<&C=��=xӓ<���α�¬9�����n
ɽ�} ����\2��mD���O��R�H
N��"B��1��^�b
�n����C�`{޽
����	���%���I�-�r����������Ѳ�R���P|��s���z����7�����l�,J<�����½�   �   �o�ЊƼ��;0��<6M>=\~x=�i�=g��=�|�=�ԩ=�!�=ޡ�=�J�=z��=�W=$o=�<@S`;�֘�XW2����l̽QH��!��Z:�4N�o�Z�D�^�mbZ�>ON�Z�<�,2(�C�f�����.�� �r	�V]1�jW����Se��5:��]@���sȾi̾��Ⱦ�;��Q���#A��h�x�A�D�N����ɽ�   �   vOr��Ǽඝ;6z�<�A=41|=�d�=e��=���=�(�=��=�j�=�L�=�+�=��]=��%=�)�<���;��:0��#��~�ͽթ�@ #�)=�ʝQ�r�^��c�}�^�5�R���@�2�+�
��Q��%���A��_��'��CS5�̘[�d����e�����������5̾�0о6̾ܝ��ُ��cǗ���|�\�G�
��Q̽�   �   �o���Ƽ`�;��<�M>=�~x=�i�=���=�|�=�ԩ=�!�=���=�J�=���= W=�o=��<`c`; Ԙ��U2���Vk̽�G��!��Y:��2N�C�Z��^�?aZ�NN�J�<�.1(�Z����
�X-��� ���P\1�;W�I���d��Z9��n?���rȾh̾��Ⱦ�:��z���e@��#�x�4�D�u��i�ɽ�   �   ңi��tƼ F\;B��<$I4=�&m=�W�=�4�=z̠=��=�e�=n5�=o/�=0�p='C=��=�֓< 	��ȱ���9�섑��ɽB| ���Z2��kD�ŚO���R�	N�� B�y	1� ]��
�8����@�ax޽����	���%�a�I���r�B�������ϲ�w���oz�����4y�������g�l�+H<�
�c�½�   �   \9b�4˼ 9�:螷<�n"=�PY=$΀=�+�=�5�=�c�=�*�=(ވ=�Zu=�O=`� =>v�<h$<P�������H������bŽ:���dp��s&�a�5��>��x@�8;��Q/����nw������]׽�LŽF�½��ѽ���1��X�4���Z�u��<}������\���f���P����w��
����悾`[��T/��[�Bĸ��   �   @�]�86ۼ��N���<�(=��;=
�b=>|=�]�=L��= ~=�Qh=�~H=P�=v��<x�X<�w�,B��6(��Dd�aᚽLEĽ��콣��6��n $���)�-�)�,�#�����H���f�̽����x��6鞽�����˽�q��'{���<��_��x��j/��}����o���u��wב�te���j�U8F�� ��*���Ů��   �   p�a������"��c<(��<�=��8=,�P=��[=��Y=�~K=�\1=��=�5�< <)<`�|��������b�N�~r��\5��xɽ���� ���
�������b���	�ݔ����ݽ�h����a����p��k������W����Ľ�����7�R$9�$OV�8�n���P��,����z�Hpg�?�M�='0�&���=��˧��   �   ��r�ޥ�0��� NT��7<�6�<�9=��=D$=�/=mW=��<TЂ<��S;��4���ռ`6)��e�0w���穽j�����ֽ.�车������b8��a��6�� �߽��ƽ������a��5�8�"��Fs(�f�U��w���칽,�콯	�f^*��@���O�]�X��8Y�PMR�n�D���1����	��(�ֽeϦ��   �   �D���N��f
�����ې�P�; �< �<���<���<�C�<�2�;�.˻����0����\�����,ӫ�|�Ľ�gؽ� 罦���j��z���4g�q轼�ڽ��ǽbY���J�� �p�|�7��r��R���Ɇ���v�������弎�,��rw�7���vԽ�����-��"���+�F*/�L�,�&x%�	���E��o���;ҽ�6���   �   =o������S��S��x��ȯ9���	��Wm;�e�; �;�㥻|툼`����J�����.��S�Խ������d
�U�����R/�� ����ؽ�m��Zm��Ȇ��tS�BN�hn��0�9��w	���m; ��; �; ���4ሼz���J�� ��0*����Խ��񽸿�vb
�v��$��@.�f �b��ؽ�n���   �   0�ǽ1\���M���p�h�7�Bx��]���Ԇ���v�̨����6�,�>zw�i¦�!Խ����|0�� "�H�+��,/���,�z%�~���F��p���;ҽ 6���C���N��b
����P��� 7�;��<�&�<t��<D��<�M�<�^�;��ʻ0������̑\�����'ϫ���Ľ\dؽ��潀��ti������g��r轮�ڽ�   �   ��J�߽��ƽF���3���a�v
5�������x(���U�Q{��}𹽌��"�a*�z@���O�R�X��;Y��OR���D���1�,�����ޙֽWϦ���r����P����T�88<>�<�==A�=$=�3=�[=H�<�ڂ<@JT;��4���ռ�/)���e�1t��a婽[���X�ֽ���������K9�Bd���   �   :d�d�	�<�����ݽ��hğ��d����p�N�k������Z����Ľ�����9��&9��QV��n���������>�z��rg�,�M��(0�*���>�Ç��a�T�����"��m<���<�!=ԝ8=&�P=�\=B Z=B�K=^`1=�=�>�<hO)<`F|�\󚼶����N��p��4���ɽ���X� �>�
�������   �   ��)�ą#�.��<J���&ͽ9���z���랽���(˽�t���|��<�J�_��y���0��扗�0q��#w���ؑ��f���j��9F�� �-,���Ʈ���]�$5ۼ�xN�,�<�*=��;=R�b=�|=�^�=���=�~=�Th=܁H=��=���<��X< :� ;��%�<Bd�����EĽ\��%��
���$�0*��   �   Bz@��;��R/� ��x������_׽OŽA�½��ѽ���h����4�6�Z�d��E~������������������y������炾ba[��U/�}\�Ÿ�:b� ˼ L�:���<�o"=0RY=�΀=�,�=�6�=�d�=�+�=?߈=0]u=��O=� =�{�<�r$<pw�����R�H�S����bŽ�����p�Rt&�\�5��>��   �   ��R�	N��!B�t
1��]��
�ė��LB὿y޽G����	�s�%�]�I���r�讎�،���в�S���R{��|��z����u���t�l� I<��
�*�½��i�\uƼ�H\;0��<�I4=�'m=PX�=~5�=͠=���=vf�=6�=90�=ԩp=�(C=��=�ٓ< ��LƱ���9�����ɽv| �s�3[2�glD���O��   �   ��^��aZ��NN�Ѧ<��1(�������
�.�,� ����\1��W�����d���9���?��2sȾh̾�Ⱦ8;��搫��@��Àx���D������ɽ��o�T�Ƽ`�;6��<N>=,x=j�=�=�|�=թ=*"�=R��=&K�=
��=�W=�p=h �<`q`;�Ҙ�U2����Ok̽�G��!��Y:�W3N���Z��   �   L��((��u��ӽ�eĽ��H(��o5ӽT|���
��L�z��Oˤ�PɾH��Z�����L���� �B�����VC�.쾲�ž%j��B(q�e1,�	�߽��t�����DU<�_=H\g=��=S��=2�=4R�=���=|�=ZS�=fˆ=Xsg=\�:=��=$Н<�͂;��M�(H���1F�G��D���F�Ƚ@�߽���   �   �K�TF�HUݽ�ͽLH��ٶ��|�ͽ2=���c��5H�(r������J~ž�o�X��A����������dA�u����>_¾Q���m��<)�;ܽ�$p�����=W<
=�te=�,�=�;�=ZU�=豩=�j�=�g�=`9�=2?�=�]=�m0=ҿ�<Ԩ�<��:xn�x��]J��鈽�@��0 ǽ+�ܽ�`��   �   ��W۽j�ν�ﾽ;q����췪�``���	�z��t;��kq�7=���i���ܾA���s
�����~����1�
�����)ܾv}��hד��)a��� �&�нX�b�|���0�Z<\f=@X_=A�=�̘=f��=޺�=��=x|�=l̅=��h=ڶ?=�=��<p]<F���
�������W�E"��H�����½\lս���   �   �#Ͻ>Lƽ�>�������W���Ɛ�lӒ�9ң��nǽ� �	�'��BY�����%���Ⱦ�h���������23�<������L�ɾ|H���Ї�O����O��ʺO�@�x�`�Y<b�=��S=:6�=�?�=�6�=n#�=��=���=lga=h�9=�=��<�< ���d���V4��5:�xr�]Q�������ɽ�Y�ʽ+�н�   �   f;��:묽W���Q\���rx��ef�vwh��	���Ģ�ս����:��gn�0I���g��wɾ��ݾ�������5ྠB̾�精�h����q��
9���X�����:�H�]�heJ<=P	B= /k=�!�=|�=���=^Rl=d�L=�$=���<@�<`�>;x�+��l������E�vls�q���������ƿ���T��|쿽�   �   KR��2V���0~���W�zr7��#�>�"�P	;���q��ऽ�+�t��-�D��Uu����R���p����Ǿ<m̾3�ɾY���֮�}���ǁ���Q��!�ڇ�����)��SU�x[#<^��<`(=K=�'\=�Y\=�L=��/=-�=PU�<���;06�� ������O���~�	k���}��k���*�� ���w������&t���   �   q���`6s���D������D5���Ѳ�U׼���>�b��"��xg潆+��4B�)Qk������ ��򒢾<��Z���%靾E���Y��v�Z�S�2�X7�T�̽J扽��� �l�P͵;�ŭ<l,=�{!=��+=�S$=�=��<؆:<�g���-��z!���h��������	AƽRս�Dݽ�E߽O�۽B�ӽ�ǽ�(�������   �   �t��d�J��p�,_���fW���ջ���� �廰o�4�� Q� V��T�ܽQ��K2�d�Q���k��)~�b���;S���z|�� j��Q�V�4��x�9��е�6�������� 鲺��F<b�<<��<���<���<�Hy<��;Zl����t$d���|�ɽN��D��0�l���������9�����66ݽ:I������   �   �{��3.�8-Ѽ��3��l:��<��H<ح7<�:�;�ӻpټ�~&5��9��Z!Ľp������v�-���=�m.G�S1I�.D��8���(�z��,��,�ҽ�U��^�{�>5.�2Ѽ��3���:��<��H<��7<��;��ӻ輼/5��>��'Ľ���#��>�-���=�@2G��4I�zD���8�H�(�9�������ҽuV���   �   x����̤�� ����F<�h�<���<ھ�<4��<0_y<�";�;l���td��	��h�ɽ�ｸA��-�k��ߙ�P���7�����4ݽ�H������u��J��s�Pf���vW�ֻ�ȉ��������!��Q��Z����ܽFT�CO2�b�Q�9�k��-~�����OU��|~|�=$j���Q�|�4��z�9
��ѵ��   �   �扽���(�l��ڵ;tʭ</=�~!=�+=X$=��=��<��:<�,������p!���h�Q��G����;ƽ�ս�@ݽB߽��۽��ӽ6�ǽ�(��D�������n9s�:�D����<
�@>���۲��_׼���<�b�'��al�o.�M8B�Uk�������O���r>������:띾��0[���Z� �2��8�ɟ̽�   �   �6 )�HRU��_#<���<p!(=�K=�*\=�\\=��L=�/=o�=Ha�<� �;�����|��ƦO��~�xg���z������r������;���W��u���S���W���4~��W��v7���#��"�~;���q�:䤽�/����D�CYu����ET��
s���Ǿ�o̾|�ɾ [���خ����dȁ�u�Q�=�!�����   �   a�����:�8�]�hJ<K=�
B=�0k=�"�=X}�=7��=�Ul=x�L=��$=��<TK�<�:?;n+��`���}���E�8hs�ڛ����\��������U�����<���쬽=���F^���vx��if��{h�5��FǢ��ս���:��jn��J��ri��~ɾ�ݾ^��H������7�cD̾
鲾�i����q�N9����   �   B����O���x���Y<)�=��S=�6�=�@�=�7�=�$�=6�=* �=�ja=$�9=�= ��<X�<�ׁ������0�<3:��r��P��p���5ʽ�'�ʽL�н=%Ͻ�Mƽ�@��U���fY���Ȑ�AՒ�;ԣ�#qǽO ���'��DY�B���$'��{�Ⱦ�j�ܗ�����r��4�����{�澏�ɾ�I��Tч�<O�����   �   ��н��b�����@�Z<�f=�X_=��=\͘=��=���=��=q}�=�ͅ="�h=t�?=�=��<�g< 3�����Z����W�"��g����½mս��$��8X۽��ν��~r��e��A����a��@�}���u;�mq�>���j��F�ܾ�����s
�6��<����̩
�����*ܾ2~���ד��*a�V� ��   �   qܽ"%p����� >W<d=>ue=�,�=�;�=�U�=N��=Fk�=jh�=�9�=�?�=`�]=Ho0=d��<8��< ;�:n�����\J��鈽�@��� ǽ��ܽa�L��F��Uݽ)�ͽ�H���ٶ��ﹽX�ͽ7>��Qd��6H��r������~žXp龷�B����I������A����l辔_¾����nm��<)��   �   ��߽x�t�0��� FU<%`=r\g=)��=h��=A�=DR�=���=��=hS�=eˆ=\sg=X�:=p�=�ϝ<�̂;��M��H���1F�e��b���b�Ƚ[�߽��\��/(��u��ӽ�eĽ��Y(���5ӽ�|���
�=�L����kˤ�8Pɾg��h�����S��ģ �A�����NC�.쾚�žj��(q�;1,��   �   �ܽ�"p�h����BW<H�=�ue=-�= <�=�U�=j��=^k�=~h�=:�=�?�=��]=�o0=���<���<@W�:h�m�v�� [J��舽�?��6�ƽ2�ܽ�_��J�nE�nTݽ��ͽ�G��Zض�3ݠͽ�<��`c�l5H��q��C����}ž8o��eA�G�����&��A���T辦^¾ͯ��4m��;)��   �   ��н��b�hz��`�Z<�h=,Z_="�=�͘=J��=λ�=��=�}�=�ͅ=��h=�?=l=�<0m< %��0�������W�$ ��)�����½Wjս��*��<U۽��ν���o���������
_��(佮���s;�ojq��<���h��$�ܾ%���fr
�؜��}�:����
�����(ܾk|��~֓�U(a�~� ��   �   T��ʵO���x���Y<~�=h T=~7�=�@�=�7�=�$�=z�=k �=Vka=��9=�=T��<�<�ȁ�ԇ���-�|/:� �q�$N��W����ƽ�^�ʽN�н!Ͻ�Iƽs<��d����U���Đ��ђ�IУ��lǽ� ��'�;AY�����$����Ⱦ]g�D���������;2�]���;�澮�ɾG��Lχ��O�����   �   ����z�:�8�]�hwJ<=�B=^2k=`#�=�}�=���=�Vl=�L=>�$=���<PM�< O?;Xg+�`\�� {�f�E��cs�#������ϻ��Q���追�7�� 謽Y����Y��hmx��`f��rh�k�������ս
���:��en��G���e���ɾ��ݾ�뾼��Y�쾦3྇@̾�岾g����q�j9�ҡ��   �   ֑��h)�;U��p#<ֶ�<�#(=(K=�+\=�]\=��L=��/= �=�b�<�'�;X�������^�O��~��e��Ox����������������q ���o��QN��~R�� *~���W��l7���#��"��;��q��ݤ��'�5��|�D��Ru����P��un��L�Ǿ�j̾��ɾ�V��kԮ�d���?Ł�?�Q��!����   �   �ች��`�l�P��;�Э<X1=^�!=P�+=�X$=��=@�<p�:< '�����o!�B�h�f�����[:ƽ�սS>ݽ?߽.�۽t�ӽ��ǽ�#������"���j.s�Z{D�J������)���Ʋ��I׼���x�b�����b��(��1B�kMk�Ն��i���}����9��Ҕ���松����W����Z�߉2�S4��̽�   �   w��p��D��� ��@�F< m�<��<<��<��<(by<�-;9l�P���d�	����ɽ�&A�-�|��������6�"���@0ݽ�C�����ep��"�J�8i��Q��NW���ջ�v���y廐W����TQ��Q����ܽ�M�H2�]�Q���k��$~������P���u|�fj���Q���4��u� �p˵��   �   �|{��,.��"Ѽ0�3�  :�<��H<8�7<PA�;��ӻ$ؼ��%5�49��� Ľ����I���-�+�=��-G��0I�(D���8�x�(����6����ҽTQ���|{�~+.��ѼP�3���:8<x�H<��7<�h�;��ӻ�ʼ��5��4���Ľֆ����n�-�a�=��)G��,I��D�߾8��(��������.�ҽ�P���   �   �p��6�J�l�`X���\W� �ջ`���p���l�����Q��U���ܽ�P�pK2�(�Q���k�)~�����R���y|��j���Q���4�Aw�z��̵����6��ؖ���ױ�X�F<�r�<���<���<Ԯ�<�vy<@�; l� ��4d�����ɽ�
��=��)�t�������4�>���X.ݽ�B��k���   �   ���,1s��~D�"�����L2���ϲ�pS׼����b��"��:g�h+��4B��Pk�ֈ��� ��ɒ���;������蝾���"Y��6�Z��2��5��̽�≽�����l�`�;�ԭ<�3=0�!=��+=�\$=��=t�<(�:<�P���f!���h�G��ު��?5ƽ�ս :ݽr;߽R�۽v�ӽ��ǽS#��Y����   �   �O��T���-~���W��p7��#�l�"��;�(�q��ऽd+�[���D��Uu����R���p����Ǿm̾��ɾ�X��_֮�����Ɓ�j�Q���!�$��(����)��;U��s#<P��<v%(=TK=T.\=�`\=TM=��/=��=�m�<�Z�;���������>�O�"�~��a��u��`����������0���� ���p���   �   R9���鬽,���u[��Dqx��df��vh��	��ZĢ���ս����:��gn�'I���g��lɾ��ݾ�����쾲5�bB̾@精kh���q�
9����'����:���]�0xJ<�=B= 4k=\$�=�~�==�Yl=��L=��$=n��<4X�<��?;�N+�,P��(u��E�_s�J���N��򯽸����Q���鿽�   �   _"ϽKƽ>�����<W��iƐ�/Ӓ�
ң��nǽ� ���'��BY�����%���Ⱦ�h��������x��'3��������ɾ=H��?Ї�nO��������O���x� �Y<��=(T=8�=�A�=�8�=�%�=��=��=�na=h�9=Չ=���<@�<0������0*�V,:���q�`M������ƽ���ʽ:�н�   �   '��aV۽�ν6ﾽ�p�����ķ��D`��z	�n��ut;��kq�2=���i���ܾ<���s
����~����(�
�����)ܾQ}��;ד�w)a�W� �'�н>�b� |���Z<�h=�Z_=r�=Θ=Ʋ�=m��=��=�~�=�΅=��h=��?=#
=��<8x<@��t������2�W����
�����½�jս���   �   jK�F�UݽR�ͽ+H���ض��j�ͽ&=���c��5H�&r������H~ž�o�X��A����������`A�p����,_¾;����m�P<)��ܽ�#p�����hAW<%�=�ue=,-�=%<�=V�=���=�k�=�h�=�:�=x@�=�]= q0=J��<l��<���:��m�f��8ZJ��舽�?��C�ƽl�ܽ�_��   �   P{M���J��kF�>^G�D�U�2|�$���ݽ�L�<�U��Ð�Å���\򾚦�,�/��G�D?[���g�u�k�s�g��/[���G��/�n���p����,����6�o�߽X�[���$�O�<V,A=���=@�=E��=�=���=M*�=Ǐ=8X�=d<]=��6=��=X"�<0�f<�.q;p�ڻ�0��P�ּ����4*���>�lZJ��   �   ��J��<F��@���@�B�N��s�(���8�׽u��^Q��ٍ��ٺ�o����c�,�<hD��hW�z�c���g��c�hW��>D�g,����V�龳L������$v3��B۽<�U�������<d�@=��=�:�=�1�=fϤ=���=ȁ�=�U�=PKt=ԁO=��'=p�< �< &*< �`9� �l����s缌���-���?��?I��   �   �B�>�9���0��.�>L9��[�Ǧ����ƽ3��C��e��4������
��]#��":�ICL���W�0\�dX��nL�s::��2#�;d	�Ƚݾ"֪��Ty�i)���ͽ��D����Xw�<�>=��}=L�=��=�a�=�=_f�=0�s=R�N=6�%=���<H �<0�< �z�p�*� N��������}&��8��C�z�F��   �   l�8��\(�Lr�ھ����6�:Js��q�������.��hp�(����=̾s���Y�*���:��E���I��E��O;���*�/�������ʾ�<��f�c���?.����+��|�����<�:=<<r=��=8��=�_�=�)�=d�b=�z;=:o=�<�.6< mι0�5�$n��d�����H_+��2=�I�ζN�4�M�r�E��   �   �0�¨�t����޼ �߼����;�����:xͽ�w���N�ے���T����ܾ$����h�$���.��2�u/���%�����7���޾	t�����H�H�	�17���� ��H��<�1=d`=��v=R�x=Ԝh=6ZI=4J=H�<�eF<�]�諆�d[�(�&�\{L�b�h��{��U��/��:��>�s�2�a� �J��   �   �#/��J��Ǽ ۖ�����0���0���D�G�z��������(��e��&��Ҍ��,wݾ����:��){�n���-��I��� ����E+��bi����k��6+�;4�΅�0m���;��<�F"=@#F=\R=�YH=�`+=���<P��< (\��������[��?��N��������½�pŽ�5��\(��O���v���툂� XZ��   �   ,�8� ��H����&�0չ���ջ(�c�}�?V�W����E��84�L�m��V��k����ξ��侢����4��"u�p:Ծ'_��m6���~���C���E��4�Y����� a�;H �< #=��#=�"=�%=��<���;�<�����rh���Nн#+���g	�T8��-�Dz�%�
�X��*���d���l���Ry��   �   z_Q����x
���]����;��;���:�f�dX�f^��a��b����2�-Ud�\����栾�貾���&ľ)����\��֨��ǔ��{���L�/��W�,ƙ�@0�<���`�y;��<��<���<���<<т<��:���9�?�� �Խ�	� 0%���<�\M�eGV���V��bO���@�h!-���]!���cƽ�����   �   �Sz�L_���q�@)�:(EH<dv�<8�<(�<`���Kм�)V�&Q�����
�#��J�I n���������]��j]��5ꌾ�ȁ��8f��oD��� ��>�������Pz�^��q���:�<H<�p�<� �<��<0L�� [м3V��V��j���#���J�n%n�y���㮏��`��/`���쌾.ˁ�j<f��rD�e� �sB��S���   �   ș�B0�\�����y;��<���<x��<t��<�ۂ< 2:@ޤ���9�J��2�Խ�	��+%���<�<WM��BV�E�V�H^O���@�1-�V��l���`ƽǥ���]Q�8������]�@��; ��;�*�: |��e伨^�g�����W�2��Yd�񭊾y頾�벾1��I)ľK����_���ب��ɔ��|���L�-1��Z��   �   ;G����Y�컬�`a�;T�<�$=e�#=��"=I*=<�< ��;P�<����gh�製�Gн�#���c	�q4�7*��v�"�
�D��%���a���j��dPy�N�8���� "��X�&�`칻�ֻ@�c�0��FV�����VH��;4�W�m�PY���m����ξ����������Fx�?=Ծ�a��j8���~��C�����   �   �6彊υ�p� �; ��</H"=l%F=LR=�]H=de+=��<���< $T�T锼��B�[��9��2~�������½�kŽM1���$��]���]��������VZ��#/��K�DǼ�ߖ��������8�����G�疝���콤�(�8�e��(��<����yݾ��������|�-��@/��K��� �Z��L-���j����k�L8+��   �   )��8��x ����ܶ�<�1= `=�v=@�x=|�h=�^I={O=hT�<�F<�������TI�
�&�drL��~h��{��R��| ��*
����s���a���J���0�
���w����޼��߼6��;�O���k{ͽ�y�Z�N�n���V��6�ܾt�l����$�2�.��2�/�%�%���� 9�~�޾�u������H��   �   ��s/��J�+� ���$��<�:=d=r=r�=H��=4a�=,+�=@�b=v;=et=T��<G6< :˹x�5��a��������Z+�/=�vI�6�N�|�M���E�2�8�X^(�t���F��6��Ms�)t��������.�kp�����P?̾f���v�Q*��:�v�E�?�I�g�E�5Q;���*�"������ʾ�=��Ȟc��   �   %j)�u�ͽ��D���绌w�<��>=��}=��=���=�b�=�=�g�=2�s=��N=��%=���<p�<��< �y���*��G��<����h|&�@�8���C���F�ڶB�Z�9��0�`.�.N9�^�[������ƽ%4�6�C�ff�� 5��̴�
��^#��#:�CDL���W�.\�YX��oL�>;:�o3#��d	���ݾ�֪��Uy��   �   dv3�/C۽t�U������<��@=��=<;�=a2�=�Ϥ=C��=v��=@V�=�Lt=��O=l�'=d�<��<x-*< �b9� �����q���̘-���?��?I�.�J��=F���@���@�l�N�Z�s���2�׽��-Q�Zڍ�rں�,��'��߃,��hD�	iW��c��g���c�xhW��>D��,�0������L��蹃��   �   ��6��߽ʤ[���$��O�<�,A=���=\�=W��=*�=���=]*�=Ǐ=9X�=p<]=��6=��=D"�< �f<@-q;жڻH1����ּ����4*��>��ZJ�t{M�ΧJ��kF�\^G���U�\2|�R��/�ݽM�x�U��Ð�녾��\򾰦�B�/�*�G�Q?[���g�y�k�q�g��/[�~�G��/�n���O����,���   �   \u3��A۽4�U�`��T��<��@=�=r;�=�2�=Ф=c��=���=\V�=0Mt=�O=��'=$�<��<�/*< nc9 �����o�z���-���?��=I��J��;F���@���@�2�N���s�������׽(���Q��ٍ��ٺ���x���,��gD�hW��c��g���c��gW�>D��,�������L��9����   �   +h)���ͽ��D�����{�<�>=��}=:�=
��=�b�=K�=�g�=��s= �N=R�%=���<�	�<�<��y��*� D�����V���y&���8�H�C��F��B�J�9���0�>.��I9���[�������ƽ\2���C��d��Y3�����1
�E]#�
":�kBL���W�6\�lX��mL��9:��1#��c	���ݾժ�KSy��   �   ��a+��Z�+��^��<��<�:=�>r=��=���=�a�=p+�=��b=�;=�t=���<�I6< �ʹ��5�p^�����8���W+��+=�lI���N���M�R�E���8��X(�dn�P��N���6��Fs�p���}��~�.�gp����K<̾Ȓ��]��*���:�ȵE���I���E��N;�Z�*�~�����2�ʾv;��)�c��   �   ���3��P� ��@��<h 1=�`=f�v=4�x=0�h=@_I=P=�U�<H�F<������,G��&��pL��|h��{��P��d�������s�Χa�J�J��0�F��$j����޼��߼�}�p;�R���euͽ v���N������R���ܾ�
������$���.�[2���.� �%����6�N�޾r�������H��   �   |/�.ʅ�\`༠A;P��<K"=t'F=�R=�^H=0f+=p��<(��< �S�蔼�V�[�/9��g}�������½*jŽc/��O"������l���g����OZ�Z/��D�HǼ�Ж�0����y��L���ĞG�J�����콌�(��e��$�������tݾ�������ty�����+�RH��� ����(��Bg���k��3+��   �    @����Y�����0��;�
�<�'=}�#=#�"=P+=��<� �;�<���pfh��磽Gн�"��pc	��3��)�v�-�
��������^��Ig��bIy��8��������&�0�����ջ��c�|q�f8V�K���(C��54���m��T���h����ξn��.󾋻������q�I7ԾG\���3��a~��C����   �   ����70��x�� $z;��<t��<���<\��<�݂<�c:�ܤ�(�9�����Խ�	��+%���<��VM�BV���V��]O� �@�-�������]ƽp����VQ������~��7]�0Ɇ;���;�^�:�O�K�j^�]��h���2��Pd�ި���㠾�岾����"ľ�����Y��Ө��Ĕ�A�{���L�v+��Q��   �   �Fz��U�Ȋq��д: TH<�{�<��<�< ��hJм()V��P��N���#���J� n�����૏��]��,]���錾�ȁ��7f��nD��� �
<������fJz�`W�X�q���:�ZH<���<��<�<�蝻�<м� V��K������$�#���J�8n�󚅾����Z��fZ��H猾(Ɓ�|3f�#kD� � �8������   �   RTQ���(�~��M]�@��;p��; ��:@b��V��^��a��B��l�2�Ud�L����栾�貾����%ľ�����\���ը�2ǔ�,�{���L��-�HU�[Ù�$:0� {���%z;�<l��<<��<���<��<��:Τ��w9�|��`�Խ�	�_'%�2�<�&RM�V=V��V�0YO��@��-�S��L���ZƽW����   �   ��8�������(�&�@�����ջȹc�8{�j>V�����E��84�6�m��V��k��z�ξ��侌��������t�0:Ծ�^��
6���~���C�����B��8�Y�L���`��;��<M)=Ç#=I�"=j/= $�<P3�; b<�����[h��᣽.@н����_	�0��%��r��
����6�཮[���d���Fy��   �   �/�E�Ǽ�Ԗ�p������ �����G�4���u����(�Ӫe��&��Ɍ��%wݾ����4��"{�f���-��I�l� �����*��
i����k��5+�Z2�̅��d� 3;h��<L"=$)F=4R=�aH=Xj+=��<�Ć< L��֔���r�[�[3��dw��z��к½�dŽ�*��H���������ւ��8NZ��   �   .�0�B��\m���޼��߼���;�u���xͽ�w���N�Ԓ���T���ܾ"����g�$���.��2�n/���%�}���7�f�޾�s��M����H�O��5����������<� 1=`=8�v=��x=l�h=<cI=�T=a�<@�F<�[�h���t5�z�&�|gL��sh��{�`M��}�����ޭs�֥a���J��   �   .�8��Y(��o�$��t��(6��Is��q�������.��hp�$����=̾n���V�*���:��E�ލI��E��O;���*�!�d�����ʾ�<���c�>�%-����+��h��X��<�:=�?r=��=���=�b�=�,�=D�b=�;=�y=X��<�a6< �ǹ�q5��Q��l�����R+�z'=�hI���N�n�M��E��   �   `�B�2�9�"�0��.�|K9���[�������ƽ3�޼C��e��4������
��]#��":�ICL���W�.\�bX��nL�n::��2#�1d	���ݾ֪��Ty�-i)��ͽh�D�����z�<�>=(�}=��=���=�c�=5�=�h�=2�s=$�N=��%=4��<��<�	<��x�p�*��<���������w&���8���C���F��   �   Z�J��;F�P�@�N�@��N���s����#�׽p��ZQ��ٍ��ٺ�l����d�,�:hD�~hW�z�c���g��c�hW��>D�e,����J�龥L�������u3��B۽x�U����l��<Z�@=
�=�;�=�2�=NФ=ο�=��= W�=�Nt=��O=��'=

�<��<�7*< ^e9�
 ������l缂��h�-�z�?��=I��   �   �Ốs񻈼%��D������T�S�?����D	�Y�M����5 ̾�<��0,���R��4x������䙿1S���<��jS��*ڙ�V���8�w�ĮQ�a~*�˳��ľ^���ZE2�H0ʽ�&�@5+;�
=`�b=fՌ=�J�=�X�=�\�=$o�= h�=�e=trA=\�=�
�<��<��o<�a<��Z;�XY� ���PQɻ�𻐙���"��   �   @'� ����/�� �r�K�ç�����vI������4Ⱦ����)��
O�\�s��X��J��m����y������I��@���ds��N���'�lY�-:���$��f�.��aŽ�� ��Z;�\=�a=^�=���=b��=���=��=�x=T7U=X)/=C�=<��<�p�<�<< �_;����������(�(6��������   �   8���9黨��H W��,ȼ�5�N	��e��Bu<�$U��sּ�����2 �<D�!dg�qY��U��������r������#я��d���8g�T�C�������Yݶ�.2��$�Ɓ���$�@߯;/�=�-\=���=b/�=�%�=D�=d�r=x�M=�#=���<�"�<�d< D>9 ���G�8~�����𙼀l���E��h�h��9��   �   Ѝ<��C�Ȼ���T���2��7.����ٽ"(���u�F��?侾��N]3��S�z�p��߃�vD���ލ��i��3���Lq�x+T��]3�\��
���Ʀ���g�$���)��8F��<c=��R=��x=,�=�ny=��]=��5=��=T�<�C�;���tR����� ��)!�`�(�l'������ ���4������   �   Dr����0뒻Pŗ�`	5��Ѽ2aN�+��F�TS����^�Ǿ�, �����;�`�T��i�N�v�#�{��Yw��[j���U��;�G��Ŋ �+Ǿg���J��.������į� �;<E�=��C=�?\=�Z=�dA=�e=l��<'�;0�0�@�fC6�
�o��$��W����������}䘽�v��8�o���D�:$��)ؼ�   �   �ͼ��N���� 2��@�Z��fg�)��5�����
�,���v��8��#3ؾ�������|5��iG��S�UJW�שS��H���6�7� ��r��۾�?��{x�E�)�xҽ\&V���_���h<=<�,=�M5=S"=$��<0G]<`��� !�>�Q������jý���D@����5M
���������ݽ,ۼ�f1��Lj���$��   �   �������W�� �$;@�|;�*�а���2������%��.B�H�������پ���	��8�#�ն-�c1��~.��T%�l���L���޾���µ���AJ��	�1���r���ֻ�ށ<�+�<�;=��=�<г�;�h��^�,����s�ҽi���R%���<�ePM���U�j�T�S�K��;�*�%��W����s����t��   �   �`�̕�����gp;x <x�<`��Զ����P��i��c$J��/������˾���pC��c	�����b
��2��f��Ҿ,ⰾ覎�g0[�k��,Խ��w��׼��w�΁<4��<XX�<���<�:�E�� 7R�+��>� �V�*�pET�0�y�-��������ğ��N��X���~�k���F�F ������a���   �   �`��ƍ0��Q�� 7';��b<�K�<h�F<����� ����]�e�����>	B���x�
N��5���H,þa?оw�վ��Ҿ�Ⱦ�ȶ�z��M3����Y�*�&���｣]���0� N���;';��b<�F�<�F<@o��,/���]�}������B�v�x�<Q��ǚ��!0þgCо��վ��Ҿ� Ⱦ"̶�}���5��n�Y�"�&����   �   �Խ>�w��׼ �w�@ρ<��<�^�<D��<���:5���,R����C� ���*�@T�#�y�����|��u��q���K��������k���F��B ����8^���`�(��P��@cp; <��<����±���P�P�����(J�H2������ ˾��龛E�-f	���-e
��4�vj�;Ҿ�䰾����3[�����   �   �	�����p��Вֻ�ށ<P.�<_>=��=��<���;4W��r�,�������ҽ����M%�b�<��JM�v|U��T�Q�K���;�E�%��T�`�⽎���v�s��������T�� �$;��|;�P*�(���F�2�0���k(�<2B�����ə��͒پ���-����#�<�-�pe1�
�.��V%�l��NN���޾<	�������DJ��   �   6*��zҽ�)V���_���h<�=D�,=�P5=�!"=���<�c]<�T�����tQ�����;cý����;�B��I
���������ݽ5ּ�{-��n�i���$� ͼ؂N� ��� ����[�Ptg��-��8�����Ε,�S�v��:���5ؾ6������~5�JlG�S��LW�/�S�E�H���6��� �@t��۾xA��3x��   �   �J�1�������ǯ�h�;<Ӆ=p�C=
B\=�Z=iA=�k=�< h�;�[0��缸76���o�n��������~��Rߘ�xr���o��D� �T$ؼ$o��H���pЗ��5���Ѽ�eN�.��H��VS�������Ǿ�- �3��X;�`�T�A�i���v�^�{�\w��]j�|�U���;����܋ ��Ǿ�����   �   h�g�$���*���H��<jc= �R=p�x=h�=�qy=��]=��5=��=��<���;�U��@��̥��0!!�\�(�@'���x��p��`/��T����<��C� Ȼ8��������%0����ٽ�#(�֣u�� ���@�� ��^3���S�+�p�����dE���ߍ�rj��
��uNq��,T�_3�B��p���Ǧ��   �   ,3��$�����`%�Pݯ;h�=�.\=���=10�=�&�=��=� s=^�M=]�#=��<$-�<p{< D9P�߻��G�,t����D陼@f���@��P�h��9���� ;�X���$W��/ȼV�5��
��g���v<�V���׼�C��� �=D�Deg�Z�� ���j���1s��-����я�je���9g��C�;�����޶��   �   %����.�bŽ�� � �Z;�\=a=��=��=���=���=d��=�x=�9U=�+/=��=���<@v�<�G< �_; ��� 㥻 ���p#� 2���� ��'� ���x0��$���K���������wI�v���u5Ⱦ`��z)�DO��s��X��sJ��˙��Yz��
���lI��c@��+es��N�E�'��Y�x:���   �   <���$E2��/ʽ��&�@<+;Z�
=��b=�Ռ=�J�=�X�=�\�=5o�=h�=4�e=�rA=u�=�
�<��<��o<Ha<��Z;�aY�0���0Rɻ ����0$�0
�u�@�%��D��`���ȌS������D	���M�5���e ̾=��0,���R��4x������䙿8S���<��iS��&ڙ�O���"�w���Q�I~*������ľ�   �   e$����.��`Ž�� �`�Z;�]=�a=��=?��=��=���=z��= �x=�9U=�+/=�=@��<�v�<8I< �_;����pݥ�`������-�(����� �@��(-��P�輖�K�D������dvI�����x4Ⱦ����)�T
O���s�JX���I������y��Z����H���?��ds�N���'�Y��9���   �   w0��$����X!� ��;f�=0\=��=�0�='�=��=� s=��M=��#=<�<�-�<H}< �D9`�߻p�G��q��H�� 晼�b���<����h�(�9�0�� $�@���W��(ȼ�5� ���c��_t<��T���ռ������ �P;D�1cg��X����������q��ྗ�Џ�Fd���7g�Z�C�������Aܶ��   �   ��g�d���&���=��<9f=��R=��x=��=`ry=D�]=`�5=��=��< ��; R廠?��H����!���(�Z'���Ԇ�����(��@���{<� $� �ǻ؄�L���
��o,����ٽ� (�ӟu����=����+\3���S���p�߃��C��
ލ��h��R��JKq��)T��\3�>��9��zŦ��   �   k|J�e*��<���D�����;<�=��C=�C\=Z=�iA=l=�<�k�;�Y0��$76��o����\�������}��1ޘ�q��Ĉo�~�D�2��ؼ<f��x��ǒ�@�����4��Ѽ�\N�e(��`D��QS�������Ǿz+ �?����:���T��i�-�v���{��Ww��Yj���U�@�;����v� �Ǿ�����   �   [�)�qsҽV��_���h<�=��,=tR5=�""=$��<�f]<�P���
�ntQ�k����bý>�罼;�����H
�s��������ݽ�Լ��+��:�i���$�Tͼ�mN����� ����Z�(Tg��#��2����὚�,���v��6���0ؾ������z5��gG�VS��GW�y�S�˃H���6�M� � q��۾U=���x��   �   �
	�g������@Uֻ��<�5�<�@=��=0�<���;�U���,�����t�ҽڽ��M%�6�<��JM�*|U���T���K��;���%��S�p�l�����s���H�@&���%; 	};��)�����z�2����� #�r+B�<���|���m�پ���� �#�{�-��`1�J|.�VR%�I���J�Z�޾��n���>J��   �   GԽ.�w�h�׼ �u��ف<H��<�c�<���< ��:�3���+R�Z��(� ���*��?T��y�����|��T��F����J��A�����k���F��A � ��� \��,`���8����p;�, <��<�W�䩱���P�"踽J��x J�D-�������˾���TA��a	�]���`
��0��b�N Ҿ�ް�2����+[�þ��   �   
X��܀0��>����';X�b<HR�<��F<����x��ԝ]�"�����$	B���x� N��*���:,þL?о\�վ��Ҿ�Ⱦ�ȶ��y���2����Y�A�&����r[��V�0��C�� �';X�b<�U�<`�F<�������X�]����c���B���x��J������}(þ\;оX�վ��Ҿ�Ⱦ$Ŷ��v��i0����Y��&�����   �   �`��Hz�@�p;�( <X�<���(�����P��츽I��I$J��/�������˾���lC��c	�����b
��2��fﾺҾ�᰾�����/[����GԽ��w���׼�Kv��ف<ܪ�<i�<���<@f�:�$��b"R�N��r� ��*��:T�4�y����@y�����𘙾�G��b��k���F�r> �����X���   �   ؙ�|��� %; �|;��)�����Ш2������%��.B�>�������w�پ�����6�#�Ѷ-� c1��~.��T%�Z��yL�z�޾���s���*AJ�	�t�������eֻd�<t7�<C=��=�!�<�$�;�E��б,�����#�ҽ����H%��<�@EM��vU�L�T���K�H�;���%�YP��y�/�����s��   �   x�̼�gN�����  ����Z��^g��'�"5��b���,���v��8��3ؾ�������|5��iG��S�SJW�өS��H���6�&� ��r�i۾d?���x���)��vҽJ#V�p�_� �h<�=:�,= U5=�&"=\��<��]<���(���hQ���[ý,�罅7����}D
����\���Q�ݽJϼ�\'����i�h�$��   �   Tb��ȷ��ǒ�����h 5�(�Ѽ6`N��*���E��SS����Y�Ǿ�, �����;�a�T��i�O�v�&�{��Yw��[j���U���;�8���� � Ǿ2����~J�-��O���(�����;<�=��C=�E\=�Z=�mA=q=��<`��;860�����+6���o������������x���ؘ�wl���o�Z�D���|ؼ�   �   �v<�� �0�ǻp�� ������-����ٽ�!(���u�A��?侼��M]3��S�z�p��߃�wD���ލ��i��2���Lq�r+T��]3�P������Ʀ���g�����(��(B���<�e=X�R=��x=��=4uy=�^=��5=i�=p��<0��;��X.��P����*!���(��	'�
�v���|"������   �   8���"黀��HW��*ȼZ�5�	���d��5u<� U��pּ�����2 �<D�dg�pY��V��������r������#я��d���8g�O�C�������Dݶ��1��$�8���<#���;�=@0\=d��=1�=�'�=��=�s=�M=��#=��< 8�<8�< NJ9��߻��G�Pg������ݙ��[��(7����h��9��   �   �������-����"�K��������vI������4Ⱦ����)��
O�\�s��X��J��l����y������I��@���ds��N���'�hY�":���$��H�.��aŽ� ���Z;g]=�a=�=���=y��=D��='��=жx=�;U=,./=��=���<h|�<�T<�`;@E���ʥ������0(���� ���   �   p��<�J�<�6<@�źྼ�k��ܽ�&6�������ʾ���S9��k��������Pi��_�ο��ٿ�Pݿ_�ٿ�uοc2���B��fs���<i�p7�
'	��$þ�0��04�h��8������< O4="�x=EJ�=8�=k�="��=�pd=4�>=7>=���<Dc�<X�O<�=�;��;@�D;��S;0*�;��;`2<@k<p�<�   �   l��<8݆<Q5< �v������$c��]ֽ 2�Nވ�v�ƾ;�	��5�U�f������ݤ�eE��I!˿��տd�ٿ��տ�˿[!��m�������Je�'�3�6�������N���uҜ�����ώ<�3=�u=$�=��=�r�=N[v=H�R=��)=`s�< �<�P<��;��:�/!��9e�`j1� ȹ EJ;�;��<<�by<�   �   ��W<��j<��0<��:���t�L��Ž�1&������d������S,�n�Z�m���z����$���C���˿%?Ͽ��˿"f���2������5��M�Y��*��>��L����p�����_�����|5�<�/=�=i=�6�=�Ā=B�l=|1I=cM=P �<0�_<`�;@��ؙ��썬�D"�����xp��PΆ�O-��]��`	;;8�<�   �   �;ȸ(<��!< |+;xG_���)�Sƫ�8���Dg������l�>��KH���t��ݏ�ۢ�cӱ�w��Sݾ������$���)�������t�=�G��8�@��Ф���Y�d~�`Rz��2[���<o�&=�ST=�`=2#R=��.=��<�G}<��������` �b|3���Y��ep�@w�~;n��W�D�5����hF��ДI�`��   �    ����r;0��;pm�;�	�� ������d��TyF��Q��ĭξ�
�ԕ0��~X�r����] ���֦���� �����).��z���0Y�W�0���	��;�<���<��Gܽ��J�@=��,(�<��=��4=1/=��=�Ȫ<��D;�֏��T!��y�����^ƽ/*޽E��}�S��Zc̽���߷���U�������   �   �貼��̻�|R; �; ���렼HaM�Մý5�!��@t��7���(�%���g8�p�Y�W�w�ٶ���\���������V���Xy��[���9����Η�隭�dcr�j]�@b���H� 8���<��=j	=��<�gG<���g	� �}��V������В��-�t7=�_uD��C���9���(���gg��u��m��\-��   �   �3�X&��𞁻@Ɖ;�(K;�0���������;���?�4���󃼾���P���13�ufL��l`��pm�
5r�>n���a��WN��]5�w+����(���7���C�������� ʼ� L;�+�<@`�<���<t�;8[����9��T������#��L���q�9܇�#���YM����������@a��`�Ⱥ:������۽�ϕ��   �    ��.6��Ql� >e:P��; ��:��o��:/�oX�����Q�2��.������c�>�!�Z2�t=�qA�e�=�p
4�|F$�%����
ľ����/\���;�����:���a�0��;�h}<�Ac< ?;�3��>�P�4ι�:�RB���z�z���Ή��`zž3�Ҿ�ؾ�Ծ��ɾ����⠾�Ć�dW� �"�i��   �   �iٽ�y~�ĉ�p%��Ь�;�<< �Z:�����K��ڻ�Ӥ��R����_H��#LվE�����b����`�1�	��/���ܾ�q����[c�n�#�feٽ�s~�|��`�� ��;�3< �Y:�����K��໽Ĩ��R�����L��jPվ�������d�̬�4c���	�q4���ܾg�/���`c���#��   �   ���ə��B�:�p�a����;o}<�Oc< �;$$����P�dǹ����zB�d�z�ٽ�������už��Ҿ�ؾ��ԾT�ɾ�𷾲ޠ�����m_W���"��*��"1�pFl� ve:���;�y�:�o�B/�k]����T�Q��4��������Vf���!� ]2�{=�~A�_�=�>4�
I$�N'�q���ľn���L3\��   �   �C�n���*��`ʼ�L;�-�<�e�<���<৺;�I��d�9��M�������#�7�L�!�q��؇�k󑾕I��ᇔ�^� ^���`�+�:�6����۽p˕��3��������ǉ;�K;p=�����Ō�/A����?���������V�����y43�JiL��o`��sm�>8r�.An���a�:ZN��_5�w-�8������9���   �   +fr�V_��d���K��V��	�<��=�	=P �<��G<p��8\	�v�}��N��H��������-��1=��oD�DC�e�9��(����:`��o���h���-�T߲�`�̻��R;�;���򠼠fM���ý�!�lDt�:���+����i8���Y�*�w�\���Y^��k!������gX��9[y�<�[���9�p��Z��Ҝ���   �   �=����<�Jܽ2�J��E���(�<m�=��4=5/=6�=�֪<@6E;����xH!�"�y�	���Vƽ�!޽��꽲t�m��#\̽8������h�U����D������@�r;���;�g�;`������{!���g���{F��S���ξ+ 
���0���X���Q����!��[ئ�+���A"��Ԟ��_/������2Y���0���	��;�   �   �Ѥ��Y�R��Tz��6[���<��&=�UT= �`='R=��.=!�<f}< �������U ��p3���Y��Yp�tw�t0n�ܑW�h�5�~��\:��0�I����0μ;�(<`�!<�m+;O_���)��ȫ�έ��Fg�z����n�X?�*MH�X�t��ޏ�)ܢ��Ա�Fx���޾�竻��%���*�����
�t�t�G��9����   �   ���t�p�p���`�����5�<p	/=�>i=�7�=�ŀ=��l=�5I=BR=��<��_< W;��������~��X�������c��4Æ�8<-�`?���6;;P�<��W<�j<X�0< o:���L�ȴŽ�2&�В��f��V��xT,���Z����9����%���D���˿@Ͽ��˿�f��x3������6��"�Y���*�~?���   �   ΋��YO�@���Ҝ��� Ў<R3=^ u=��=ק�=�s�=p]v=ĘR=��)=�y�< �<P+P<�ʹ;��: � ��e��91� �ƹ@hJ;0�;(�<<Hfy<h��<|݆<P5<��v���� &c��^ֽ�2��ވ�)�ƾ��	���5���f�歷�Lޤ��E���!˿��տܶٿ��տ˿�!��������>Ke�o�3�i���   �   �$þ�0���3���(���P��<pO4=��x=dJ�=48�=>k�=9��=qd=`�>=\>=<��<dc�<x�O<�=�;p�; �D; �S;0)�;@�;�2<hk<�o�< ��<�J�<�6<��ź ᾼDk�Yܽ�&6�꺋�թʾ��T9��k����Ȯ��ai��m�ο��ٿ�Pݿ]�ٿ�uοX2���B��Vs���<i�R7��&	��   �   ݊���M�H��Kќ�P���Ҏ<43= !u=��=���=�s�=�]v=�R=��)=�y�<H �<�+P< ̹;��:@� ���d� 31� {ƹ�rJ; "�;8�<<�iy<d��<�߆<(U5< Qv�l����#c�P]ֽ�2�ވ�*�ƾ�	���5���f�P����ݤ�E��� ˿�տ�ٿ�տ-˿� �����v��=Je���3�ǵ��   �   /��Ւp����^�������:�</=(@i=8�=3ƀ=��l=�5I=zR= �<x�_<�Z;���Љ���}��4��L���b�� ���h7-�4���O;;x�<0�W<��j<��0<�(:����\L���Ž�0&�i���&d�����R,���Z�艅�ޭ��2$��C��=�˿K>Ͽ�˿Ne���1��U����4��6�Y�1�*�=���   �   SϤ�n�Y��|�@Mz�@"[����<��&=hWT=�`=�'R=:�.=�!�<Hg}< w�`����U �\p3�,�Y��Xp��w�p/n���W���5�̴�`6���yI�`�� �; �(<��!< �+; ;_���)�Zī�����Bg�ܳ��kk� =�jJH��t��܏�ڢ�Lұ��u��$ܾ������#���(�������t���G��7�Z��   �   �:��J�<��Cܽv�J�P���0�<8�=h�4=T6/=�=�ת<�=E;���(H!��y����gVƽT!޽N��@t����t[̽Y�������U�F���	��@෻`�r;@��;���;��������h���`��:wF��P���ξ�
�P�0��|X�O
�͞�����զ�K�m��"����,��Q���.Y���0�V�	��;�   �   �_r��Z��]��.B�����<�=!	=#�< �G<����[	�"�}��N��$������x�-��1=�boD�
C��9���(�f��&_�n��g���-�tز��̻��R;��;�H��ᠼ|[M�>�ý�!��=t��5���%�|���e8��Y���w�g���A[��F������uU���Uy�c�[���9����˔꾅����   �   C�ݎ��<����ʼ`�L;7�<l�<Т�<в�;�G����9��M�������#�$�L��q��؇�[󑾁I��Ň��:��]��(`���:����V�۽�ɕ�B
3����0j��`�;�|K;��R��+���7����?����@���E��F���/3��cL��i`��mm��1r��:n���a��TN��Z5�A)�=��!���05���   �   P��������:���a����;H�}<�[c<��;�!����P� ǹ�����yB�P�z�ҽ�������už��Ҿ�ؾ|�Ծ3�ɾ~�|ޠ������^W���"���}��P-��4l���f: ��;���:��o�P3/��S��x��Q�|/�������쾫a���!�NW2�~=�gA�b�=��4��C$��"�x��-ľ(���+\��   �   �^ٽ�h~�Lq輠ߧ����;�M< �[:X�`�K�Lڻ�����R����XH��Lվ@�����b�
���`�%�	��/���ܾ�츾1���$[c�Ķ#��cٽp~�Xz�@����;`S<�h\:�皼��K��Ի�&��v�R��|���D��Hվ����~��Z_�S���]���	�	+���ܾA鸾E����Vc�<�#��   �   *��v'�h&l� -g:���;�I�:�o�L9/��W��i�ԾQ�2��&������c�;�!�Z2�r=�mA�`�=�h
4�pF$��$�|��z
ľ����/\�A������R�:���a����;��}<hfc<� ;�����P��������uB�k�z�^���΁���qž	�Ҿ3ؾ��Ծ��ɾ�췾�ڠ������YW���"�� ��   �   d3�d��0U�����;�qK;$����Q���};����?�(���ꃼ����N���13�tfL��l`��pm�5r�>n���a��WN�r]5�f+�������[7��>C�]���>���	ʼ kL;�7�<p�<L��<�ߺ;d8����9�G������#���L���q�&Շ���E����������Z����_�а:�����۽ŕ��   �   �Ͳ���̻��R;��; i��格�_M�Y�ý�!��@t��7���(�$���g8�o�Y�X�w�ٶ���\���������V���Xy�މ[���9������꾻����br��\�a���E�@�麬�<Z�=�#	=�+�<P�G<��ZQ	�X�}��F��L�������-��+=��iD�YC���9���(� ���W�h��6b�� �,��   �   @����s;0��;0��; ���d���R���c��8yF��Q����ξ�
�ӕ0��~X�r����_ ���֦���� �����(.��x���0Y�L�0���	��;�<����<��Fܽ<�J��%���/�<�=z�4=�9/=ʙ=��<��E;�����<!��y����VNƽ�޽����k����T̽���쫎���U��������   �   ���;x�(<��!<`�+;8?_���)��ū����Dg������l�>��KH���t��ݏ�ۢ�eӱ�w��Tݾ������$���)�������t�6�G��8�*龭Ф�]�Y�~��Pz�*[�d��<(�&=�XT=d�`=D+R=��.=\-�<�}< g�����K �e3�J�Y��Lp���v�($n�J�W���5���h)��eI��}��   �   �W<��j<��0< :H����L�òŽt1&�򑀾�d������S,�n�Z�l���z����$���C���˿&?Ͽ��˿#f���2������5��J�Y��*�v>��:��U�p����^_�� ��89�<$/=�@i=�8�=Hǀ=اl=z9I=�V=��<h�_< �;�x��z��hn��4���￼�T��x���H#-� ��@�;;8�<�   �   8��<���<(V5< Mv�����,$c��]ֽ2�Lވ�t�ƾ:�	�
�5�S�f������ݤ�dE��J!˿��տf�ٿ��տ�˿\!��k�������Je�%�3�2������N����1Ҝ����Tю<3=0!u=2�=j��=pt�=J_v=��R=0�)=��<�&�<�9P<��; �:�� � �d� �0� Ź��J;3�;�<<�ny<�   �   X�=���<L9�< ;8J�8�����!Xr���������v9�5	t��ə��4���7ٿ1���\@�xP�D��zO�2�;\�� �ؿ�M������Bjq�ʊ6��a����H[a�{��(�V���.�Th�<d�Q=�}=h~�=�}=�ra= �:=
=���<(�c<֮;@Y��p`�˻����]��0��; </<G�<0��<\j�<�   �    ��<�:�<0�< C!;��ݼ�Ք� a��@m��U��l��6���o��,������տ�����
�q�

����z��'տ�T���'���Ym�4_3����@����\�eG���P�@2��S�<�rM=lsu=T�}=��n=d4O=;�$=u�<��<0>�;`R�H�#��!e�h�v���Y��.� �7���;� Q<��<`��<�   �   H�<��<\��<`mP;DTüI���n�}^��ë�4���gf,��_c���������O˿��U����b����Dw�ѿ���1��"˿\����܎�l�a��&*�zN���~���O��m�~0=� 3���<��?=�*^=�\=��B=خ=\3�<G<����������,��*�*�>�,�(J ��t�8�ļ^� D!� ]<H��<�   �   �+<<�<�at<��{;Ի���]j���؂G�~O��`��N?�6P�d������� ��uӿ����-򿰄���z�l�ӿ�_�� ���c����N�ٵ���޾iC��N�:�+b˽�� �@��: ��<�$(=�6=1=#=$2�<@�a<����D�ü8�0���x������?��}j���������(��t{y�0�9�̆���S� ��:�   �   �&��`J�;&< Ks;Ib�T�;���ý��*�5����ƾ�
��f7��i�J���y������Ϳ�ؿ
ܿ��ؿV�Ϳ�Ӽ�� ���s��Zi�,7��S	�7�þ]����� �3ꪽ��� i�;<��<�	=`W�<���<�6;�Ȥ�4p;��;����˽Q
��Z��F% ��K&���$��F�0q��:��X���*��<�4��Ǻ��   �   ��＀W"���:`i;	�pi	������
�PO^�<���+�辂��ΰF��&s�����-⡿4Ѱ�{���������|���n㢿�߿t���G��:�0#����
�Z�����F��D3�����;���<��<�7-<�c ���
�Yᆽd�н���5�LYW�:�r��Ă�V����ք�=.{�BNc�D`D��)!�����(2c��   �   b w�L���H�5�����O��P����Z�d7ѽ�.� L��l)��������"�	OH���l�gX�����>T��
[���כ�Y����~����n���J�ݶ$��/ ����Q��.�?�̽�|G�`�k�pܜ;�x)<@�g;��n���/�!��v��� �2�Vih��q����������ž+�ʾҳǾ\���#���Cm����x��iD���H�Ƚ�   �   |˽� l��O��`��,m���:�����̐�����y�G��А��}ž�����e���;�ajV��gk�(y�|#~��z��Fm���X��>��!�.x���ɾ����^�M�G=��Z��"j�H�� ;@-��\3��V�:�������X�J�����*9���Ͼ���B����L��	�݄�����s%־__���w��x�Y��8��   �   ����⸽�gD�PR��`���O[�����,�Yƨ��D��R��%��<ο����T�E$���4�ť?�'�C��@�.�6��&�F�����VƾU"��#]����.޸�@bD�M����� t[�T���� ,��˨�RH��$R��(��8ҿ�s�� �^$��4�D�?���C���@�s�6��&��������ƾ4%��|#]��   �   �M��?��]��xm���� ;����p&��޵:�<�������J�"�5��3�Ͼs��f����I���������� ־�[���t����Y�'5��v˽�l��F��Y��5m�p�:�v���А������G�WӐ�}�ž���gh��<��mV��kk�y�`'~��z�2Jm�@�X�Թ>�N!�6z��ɾf����   �   �R���.���̽��G���k�P�;�)< �g;0fn��/� ��������2��bh��m��j�����ȴžA�ʾ�Ǿ��������i��p�x��dD���F�Ƚ��v�����(�5�@v�`Y��P����Z�<ѽ.�FN��r,��������"��QH�ވl�5Z�����BV��]���ٛ�:���������n�G�J���$��1 �l"���   �   ������Z�L���H���6��P��;,��<4�<�P-<A �r�
�Eچ���н���5��RW��r���������@ӄ�:'{��Gc��ZD�%!������鱽�(c�����E"��U�: n;��:m	��Ø�<
��R^�����9��v��2�F�c)s�r����㡿Ӱ�
}���������R���墿 ���l�t��G�O<��%��   �   �þ����+� �쪽���`i�;p��<�=a�<0�<`�;`���c;�E4����˽s ��}�� �"F&��$�nA�rl�P2��Q��%����4�����`��� c�;�+<�Gs;�Pb�$�;��ý˄*�σ��ƾD
��h7� i��	��L{��M��MͿqؿ�ܿj�ؿ�Ϳ!ռ��!���t���[i��-7��T	��   �   N�޾]D����:��c˽� ����:D��<:'(=.
6=�A#=�>�<0�a<�9��\�ü��0���x����08���b��q���Jx���!���oy�(�9�`v���S� 7�:(9<<�<�dt< �{;����
aj�:�҄G��P��G�⾎@��P�Y�������!���ӿ��^/�9���r|�n�S�ӿa����Jd����N�˶��   �   fO��4����O��n�\1=� 7����<p�?=-^=�\=��B=�=�?�<0c<@i��ܞ��L��b��H�*���,�A ��l���ļ��]� � �0m<`��<h�<��<���<�cP;�WüqJ���o��~^��ī�����\g,�ac�����X���P˿� �n���tc�&���w������2忠#˿���~ݎ�D�a�m'*��   �   ��	A��.�\��G���P�`/�U�<tsM=�tu=~=��n=�6O=<�$=|�<��< a�;��Q�h�#��e�Ыv�`�Y����]7�p(�;�*Q<@�< ��<���<�;�<�<�9!;��ݼ�֔��a��Am�1V����T6���o�W-��+��{�տA��j�H
�Nq�L

�$�%{�-(տ�T���'��7Zm�v_3��   �   �a�㜲��Za���v�V���.�i�<��Q=�}=�~�=`�}=sa=`�:=:=��<��c<�֮;@V��@p�˻�����`��p��;�;/<�F�<Ȟ�<�i�<�=d��<�8�< ;\K�o8�����vXr���������v9�c	t�ʙ��4���7ٿG���d@�|P�F��xO� 2�.\���ؿ�M��姘�jq���6��   �   Z�$@����\��E���P���(W�<,tM=0uu=T~=�n=7O=Y�$=L|�< �<�a�;@�Q��#��e��v�h�Y����X7��+�;�,Q<d�<d��<x��<�=�<\�< Q!;�ݼ4Ք��`�|@m�@U��<�z6���o��,��c����տ?�����
��p��	
���*z�N'տT��V'��.Ym��^3��   �   M���}��S�O�Vk��,=� �����<��?=.^=��\=L�B=(�=�?�<�c<�h��������.���*�N�,��@ ��k�(�ļ��]� � ��q<���<P�<h �<@��< �P;Pü�G��2n�|^�ë�>����e,�_c�o�������N˿��Z���\b�
���v�þ���0��!˿����F܎�I�a��%*��   �   �޾B��B�:�_˽ȱ �@��:ԭ�<)(=f6=�B#=�?�<��a<�7���ü��0���x�����8��~b��6����w���!���ny��9��s��S��m�:8A<< �<qt< |;8����Yj�?�P�G�oN�����U>�� P��������i��6ӿ#��\,�.���ty�@k濹}ӿ�^��	����b���N�����   �   �þ����6� ��檽�����;0��<�=�c�<�<`�;�����b;�+4����˽` ���|�� �F&���$�EA�:l��1� Q��V$��<�4������뷻�z�;P:<��s;�7b���;��~ý��*�䀆�
ƾ�
�*e7��i���tx��#���Ϳ�ؿ>ܿ�ؿ��Ϳ Ҽ���9r���Wi�8*7�ZR	��   �   ������Z�����B�� &��0��;�Ƙ<��< W-<(= �ܨ
�چ���н���5��RW��r�����}���0ӄ�'{��Gc�ZZD��$!�����豽�&c�H��x9"� Շ:`�;@���c	�9����
�fL^�B������͚���F��#s�X􎿃ࡿcϰ�"y������$��������ᢿ폿�t���G��8�) ��   �   �N���.�ܢ̽jtG��k�P�;P�)<`h;�_n��~/����S�����2��bh��m��g�����ôž8�ʾ��Ǿ����榫�}i���x�\dD�A�(�Ƚ�v�@����5� #�0!��걼��Z��2ѽ�.��I���&��5��l�"�nLH���l��V�����FR��Y���՛�m���}����n�ڃJ�z�$�. �����   �   �M��9�hU���a���� w; :���!��^�:��������ʳJ��5��/�Ͼp��e����I���
������� ־i[��_t��%�Y��4�yu˽�l�(?�`E���l�H�:�����ǐ�Ф����G��͐��zžt���;c���;�gV�Qdk�ay��~�z��Bm���X�ѳ>�"!��u�;�ɾ����   �   ����׸�8XD��<���ǖ� �Z��,��Ũ�WD�jR��%��7ο����S�F$���4�ĥ?�%�C��@�(�6�ݒ&�9�b���,ƾ$"���]�/���ܸ��^D��C���Ж���Z��瀼x,������@��R��"���ʿ�+�ﾳ�M$�U�4�T�?���C���@�֓6�ʏ&�|�����Kƾ���]��   �   �o˽>l��4��:���l��:�����ː� ���Q�G�yА��}ž�����e���;�cjV��gk�(y�z#~��z��Fm���X�߶>��!�x���ɾņ���M��<�&Y��f� ��`�; ܋�����:����������J��E1����Ͼ]�ﾞ��"��F���4�}���3־rW��q����Y��0��   �   z�v�����h�5���#�����Z��6ѽ�.��K��d)��������"�
OH���l�hX�����?T��
[���כ�Y����~����n���J�ζ$��/ �����P���.���̽jyG�p�k���;��)<�Ih;�Dn�0u/�A�����f�2�y\h�Mj��E��r����žT�ʾ$�Ǿ%󼾬����e���yx�_D����Ƚ�   �   L�Ｘ$"�@7�:��;���lf	������
�(O^�0���%�辂��ΰF��&s�����/⡿5Ѱ�{���������|���l㢿�ڿt���G��:�#�������Z���XE���+�����;Pɘ<���<�l-<p ���
��ӆ�~�н���	5�6LW� �r�:�������vτ��{�Ac��TD��!�����ZⱽNc��   �   𾷻 ��;�B<��s;;b��;�.�ýT�*�&����ƾ�
��f7��i�J���y������Ϳ�ؿ
ܿ��ؿW�Ϳ�Ӽ�� ���s��Zi��+7��S	��þ8���8� �骽�	�����;���<H=�k�<���<�E;�����V;��,��/�˽�����w�- �w@&�{�$�<�fg�()�I��(��L�4�<����   �   PQ<<L!�< wt<�|;ܶ���[j�
꽴�G�rO��[��N?�4P�c������� ��xӿ����-򿲄���z�l�ӿ�_�� ���c����N�ӵ���޾LC���:�_a˽x� �@^�:l��<�*(=.6=�F#=�J�< �a<��H�ü��0�.�x�����o0���Z�������p������by���9�,b�ȞS���:�   �   �"�<�#�<,��<��P;Qü�H���n�}^��ë�3���ff,��_c���������O˿��U����b����Fw�ӿ���1��"˿[����܎�j�a��&*�mN���~����O�$m�/=� 2����<��?=�/^=@�\=��B=��=�J�<�}<@,��܍�������D�*���,�n7 �dc�Ёļ��]�`� �Ѓ<�<�   �   (��<�?�<��<�U!;�ݼ\Ք��`��@m�U��k��6���o��,������տ�����
�q�

����z��'տT���'���Ym�1_3����@����\�'G��P��"��V�<ZtM=�uu=l~=��n=09O=��$=t��<%�<���;��Q��|#��d���v���Y��� 7�`F�;�7Q<��<��<�   �   ��=��=` �<����'��oͽr�>�c蜾zR�,R,���k�C���C����迀�������&�j0�PO3��0��&�����&�Ǭ�j���-���G�h�4)�g���,����0�KQ����Ƽ�ȃ<��&=�pZ=��h=�[=�,:=�=L��<�< E��08�dV���Tv��Dۑ��=� �G�P5�; j�<��<ܿ=�   �   �
	=P/ =��<@����"��`Ƚʳ:����꾷,)���g���������(��e��Q�$�"-��:0�>-���#�0%��
�<�����g�d�&���便C��;�,�f��X�� �<��!=·Q=�[=@�I=�K$=��<�&l< =\:�P=�屼��D�����C�T}��Z?� �2�Ȳ/<�G�<()�<�   �   �6�<h��<�e�< ��L
��鹽��.����W�ݾ? �տ[�2��������ڿ������$���f$��k'���$�p�������qٿ�ų��֎��?Y��m�}ؾ�ъ� "���������8v<,�=$A6=��3=:�=H�<H�< ����Լ<�)�(�\�����^�����w�h)P��z�`����K��;pA�<�   �   ��<8�<�SO<@N��9�.���A3��|��Zɾ<����H�y�����}�ȿ��鿤������8�h���r����\��R��ȿ�����^���:G����d�ľ?X{��P��9��캒��W<b�<�=���<��h< ��<�ּ�PK��䔽y����oU�����������[ҽ��:q��l*,�LЮ��9g��   �   8�U� �:���;`*e���ּU7�����Xa�W(��ԥ����0���i�`{��5Ų�	�п�) �x���U	��(�"� �O)�ɊѿLQ������hKi��20��`��;��p-Z�+����i�psp��<�(�<��<�B;P���dA:�E��έ��l�/�B�G�!�W��y^��[�l N�,�8�m��n��6���p�z�����   �   ��3�t+�� �� t��G��
�Y�=׽Z�9��!���2׾4��
G��|�%���I᳿�˿WHݿ\(鿘����鿑w޿'b̿Z)��=�����}���G�����־���J 5��)˽,�:��4K�`�e;#�;P���M���~���Ͻ���ZrE�ft�4Z���X��Ě��X��eG��o������������R��#��"��T���   �   ���P
D��ļ�b�0���.7#�]ˣ�����h�En��Q��#��%P�'�~�1����T��4踿�ÿ�ƿ\�ÿ� ��[Ѫ�)�����)R��u$�����T7��Sih��/��1��Ve�(LE�@�����o��|�8���	�ro2��!r� ~��n;��ճؾ�R�����B���� �4��>�ݾ����֠��K��?�0-��   �   �x	��X���~;�@żP����)鼾"g��ӽ5�.�V��粽�\ ���$�%�J��co�r ���锿�O��n�������� x��J|r�ܐM��''�>�~���2?��)�1�b�ս�Re�T]ؼpXk�(.��� �瘽����ٯA��̇��6������������n*���4���8�)�5��R,��b�	����V��'���JL��   �   �TG�B���\���(b�����d�����#���Ǔ��dX@���1ÿ�@)����4�7�ͤQ�Rf�f�s�w�x���t� mh��fT�A�:�Ώ�����ľhJ���PG����������^�����i��T����������]@�!��8ǿ�=.�������7���Q�0Vf���s���x���t�qh�{jT���:����������ľ1M���   �   sA��I�1�k�ս�Ve��_ؼ8Rk� %��� �Wᘽ������A�"ɇ��2��x����b~�Kk*��4��8�u�5�O,�����	����&R�����`EL�'u	�T�� y;���ļ貓�P0�J)g�#�ӽ�.����k���� ���$�z�J�|go����씿8R��qp��i������z���r���M��*'�H	������   �   �9���lh��1�v4��Jg� IE������|o�Xs�s1��� ��i2�r�z���6��x�ؾ�L����*���� �y��|ݾG���&Ҡ�WE��?�R)�4 ���D��ļ�b�\���;#��Σ�f���h�q�����#��(P���~�1����V���긿&ÿ��ƿɹÿ1#��yӪ�	�������+R��w$�����   �   ��־����t"5�,˽n�:��3K�`�e;�I�;�U�$9��.~��Ͻ\���kE��^t�V��8T��
�������B���������������R�ߦ#����N��ƌ3�������m�@K��b�Y��@׽>�9��#���5׾���G�
�|�⯙�C㳿-˿�Jݿ�*���*���y޿3d̿-+��ϯ����}�ɱG�C��   �   �b���<��l/Z����,�i�tp��<,0�<H$�<@�B;x蔼@4:��<�����2��G�/���G�-�W��r^��[��N�0�8��g��e��ŝ����z����0�U� �:���; (e���ּ�9����L[a�U*��������0�ɓi��|���Ʋ�ݧп	�@ ����W	�*�*� �,+�l�ѿ�R��쩓�LMi�f40��   �   �����ľ�Y{��Q��:��������W<\g�< =��<��h<�Ë�x�ּVCK��ܔ�脿�����K����C������pSҽ����j���,�������f��<��<YO<`S��;�5����4��}��ɾm��(�H�r�������ȿ9�鿂��t���9�b���s����"��S�2�ȿ}����_���;G��   �   En�IؾaҊ�� "�$�4��<v<�=�C6=��3=�=h�<��<�i�D�Լv�)���\����hX������w��P��q�p���`1��;`I�<0<�<ع�< g�<@��"�b빽��.�������ݾ( ��[�����s���ڿ����`�����g$�\l'�`�$��V�����rٿiƳ�Q׎�X@Y��   �   X&�K���C��l�,�������p�<��!=L�Q=�[=��I=�N$=,�<x7l< o]:�;=��ٱ��	�\y��}��8�hs��PH?���1�(�/<�L�<�,�<�	=�/ =�<����h�"��aȽ��:�eÙ����I-)�c�g����v��#)�Hf�\R�h$��-�<;0��-���#�v%�J�y
俅���?����d��   �   )�*���,��L�0��P��p�Ƽ�Ƀ<Z�&=�pZ=,�h=<[=�,:="=Ե�<�	<�?�808�0V����Lv��lۑ�=���G�P4�;�i�<h�<��=H�=Z�=��<�����'�pͽ��>��蜾�R�WR,��k�;C���C����迎�������&�p0�RO3��0�ڽ&�����&����O�������h��   �   �&�.��'C��[�,���,����<��!=܉Q=h�[=��I=�N$=T�<�7l<�s]:h;=��ٱ��	�Py��}��8�s���G?���1���/<tM�<�-�<V	=�0 =8�< ���D�"�&`Ƚ~�:������|,)�X�g�k������+(忸e��Q��$��
-�t:0��-�.�#��$����	俿��������d��   �   �l�,ؾ�Њ���!�l�������Ev<��=�D6=L�3=|�=��<P�<pi�0�Լf�)�|�\����[X�� ���xw��P�*q�d����.�`�;LK�<�>�<��<Pk�< ����m蹽ҳ.�j���{�ݾ� ��[�����鸴�-ڿ����,����f$��j'���$���*�ӭ��qٿ�ĳ�֎�k>Y��   �   �����ľ�U{��N��6��\����W<�k�<^=Ș�<��h<0����ּ<CK��ܔ�焿�����K��ּ�'������5Sҽm���j��,�h�����f�X<H�<�dO<��26���1��{��ɾU��c�H�������R�ȿM��޺�����7�r���q������Q꿻�ȿh����]��9G��   �   ^��9���*Z������i��[p��<h5�<�'�<��B;D甼�3:��<��~��1��H�/���G�*�W��r^��[��N��8��g�%e��4���L�z��� �U� �:`Ô;��d���ּ�4��,�/Va��&������e�0���i�/z���ò�b�п$�" �`���T	��'�� �T'���ѿ�O��h���2Ii�110��   �   �}־󤐾"5��$˽n�:��K�@;f;�`�;�G� 7���~���ϽO���kE��^t�V��6T���������B������}���y��m�R���#�9�N����3���`��0C�4<���Y� 9׽��9�
 ��a0׾����G�q�|�����w߳���ʿFݿ &�-��a��Bu޿�_̿h'��������}�P�G����   �   w4��eh�Y,��,��]��-E��^��qo��q��0��� ��i2��r��y���6��z�ؾ�L����*���� �q���{ݾ0���Ҡ�E���?��(� �����C�P�ļ8�a���0#�$ǣ����T}h��k�����l#�F#P��~�S���hR���帿Hÿ
�ƿ�ÿ���*Ϫ�,��O���!&R�qs$�����   �   z<���1�!�ս�He�DLؼ�7k����4 �����6���h�A�ɇ��2��v����d~�Lk*��4��8�s�5�O,�����	����R��ᑍ��DL��t	��R��pu;���ļ$���(�8g���ӽ��.��������M �&�$��J�`o�m����甿�M���k����b���u��vxr���M�&%'�������   �   �KG�������T��򨼠X��֌������2X@����+ÿ�>)����6�7�ФQ�Rf�h�s�y�x���t��lh��fT�8�:�ď�������ľ>J��EPG�r���$����Y�L���V��|�����/���T@�"��|����$��5���7��Q�Nf�(�s��x�J�t��hh��bT�ȭ:�͌�����Ͷľ4G���   �   �p	�oM��|n;� �ļl���,�\g�ߪӽ��.�C��ڲ��Z ���$�&�J��co�s ���锿�O��n���������w��C|r�ӐM��''�0�Y���?����1���սZNe�\Qؼ6k����� �ۘ������A��Ň��.�����5��4{��g*�V�4�V�8���5��K,��	��	�����M�������?L��   �   ����,�C�P�ļp�a��~���2#��ɣ�(��ɀh�5n��K��#��%P�)�~�3����T��6踿�ÿ��ƿ]�ÿ� ��[Ѫ�&��	���
)R��u$�����.7���hh��.�90��F`� /E��K��x\o�Zi�+�����d2��r�v��2��I�ؾ'G�������� ����vݾm����͠�M>�1�?��$��   �   ��3���� ��4�=��~�Y��;׽�9��!���2׾3��
G��|�&���K᳿ ˿YHݿ](鿙����鿑w޿%b̿X)��;�����}���G�����־ꦐ��5�(˽�:��K��Rf;��;0�p$���}���ϽI|��eE��Wt�R���O��_�������=��t���Z������R�X�#���G���   �   �{U���:�۔;��d�8�ּ�5��~�JXa�K(��Х����0���i�a{��6Ų�	�п�* �z���U	��(�$� �O)�ǊѿJQ������cKi��20��`���:��-Z����ʮi��`p��<�:�<1�< C;PԔ��':�X5��n����T�/��G�J�W��k^��
[�2N���8�,b��[��a�����z�*y��   �   X!<Ȭ<(mO<`��6�<����2��|��Qɾ:����H�y�����~�ȿ��鿦������8�j���r����\��R��ȿ�����^���:G����N�ľ�W{�8P��8��L���ؽW<o�<�=���<�i<@|���}ּ~6K��Ք��|�����AB���������r�Jҽ����c���,�x��� Nf��   �   |E�<���<(n�<���f�&鹽��.�����S�ݾ> �Կ[�3��������ڿ������$���f$��k'���$�p�������qٿ�ų��֎��?Y��m�nؾ�ъ���!������	��Ev<t�=�F6=`�3=�=�'�< <@I���Լ|)�8�\����QR������w��P��g��������G�;|T�<�   �   "	=2 =��< ���$�"�R`Ƚ��:����꾷,)���g���������(��e��Q�$�"-��:0�>-���#�2%��
�=�����g�d�&���侶C���,���8��H�<��!=��Q=[=��I=tQ$=��<�Fl< �^:�'=�ϱ���뼀s��w��-缸h���4?� �0���/<LS�<|2�<�   �   F�=\�=8ď<`22���m��k�V�p��þ�!��T��C������]�鿔��N$�b*:��uL���X��;]���X��PL���9�\�#������翙u���T���zP�+��^�����e� ����>� �:\p�<^u7=z�G=�b8=q=P.�<�W<@n���������R�pg �"���w�x ̼@�b�����X�@<�}�<��=�   �   �9=@B�<�=�< �1��h�|�l��ܿ��a��8P��ƍ�3_����z
�@�!���6�\�H�,�T�Y���T�(�H���6��� �,�	��C俼��������L��R��$����`�I�r:���v:�C�<�5-=x�8=�.$=p��<8}< V1��π�L����(�ƫH�6�V��>R�&�;�PT��1Ƽh'����;���<ls�<�   �   D�<,��<tP< �4�.�Y��(����]�/۴�g	��8E�錆�gC���ڿ�������-�>�l6I�^9M��bI�K>���-�4^��W�O�ٿGۭ����'pB�w��`Ư��S� �߽�Z.� �9<j�<��=��
=x��<�u)<8���伦C��셽_H�����Xy��x绽/Ŭ�����2�e���J���qʺ�'P<�   �    �7;��"<���;� C��D�v�ڽ~�G�xɣ�`����4�v������ɿ����U�*e�v&.��8���;��T8�&�.���������ɿ�8����t�62�����?����?�,�ȽhU��J�L7�<�V�<X6m<@��x���XCG�9��%�ӽT����w$�R�)�� '�Z����	��^�و����s��`�qP��   �   t�ʼ`p������0l��,�ް���>,��W��_�ھqL�ּY�Yӎ��`����ؿ������`��:E#��e&��#��}�^���L���7ٿL���Ω��}�X��#���׾N��Ӌ%�Gܬ����@�����;�p�:��e�2� �BÒ��2߽%�ՠ?��Lc����o��+*��Ί�������j���H�6D"��)���\���M��   �   &����m���N��*��⚽t�E�l��|��%���69��Ut��(��?���%�ٿNT��0������{�J�Zm��'���rۿ����Ku��O9��w�F#��5i��h	�u�������VI�8@9���м<UX�O⺽����D��|~���������cɾ1�־��۾�_ؾU̾����]������O����W�Ͻ�   �   �|�>���&n$�������w��n߽�$<�xb���	پYe�I�DL��^��U޵��BͿ��߿���S����Y�/'Ͽ���c霿�ʀ�;�J�ZA���پ�R����:��dڽ�8i�4���4���Ħ	�F3y��5ӽ��"��g�SX����¾�u���@�œ�}"��}���bV	�S���nȾN۟���q�#S,��   �   �61��f�!7���)�����B��Φ����^a��/���
��pK�)�x�qP��V����
������¿ҿ��y��L|��� ��
|��M��� �n�������c�>l����Н<��9��p��~�0R׽��)���y����r�ྂ����&�|�>�G�Q��{^��+c��_��	T�q�A���)�]���h澋������   �   ��|�J�&� %ͽh�q�"��b?��j��<ǽ�I"��Fw����B��J��F�>�5�a� ����⌿8씿�엿t������&��fOe�["B�	������������|�ބ&�� ͽ��q�H��B���j�Bǽ�M"�ELw����#��N����>�X�a�n���6匿�[�����c��^Se��%B�ْ�,�������   �   ���e�c��n������<�<8��k���~�cK׽��)�:�y����P��n���&���>���Q�$w^�%'c�t�_�^T���A�3�)�n��d澻	�����21��`㽐3���})����̶B�SҦ�����ba��2��S"�����"K�%�x��R��۸��������¿¿�Կ�Y|���~��#���|�&�M�� �8���   �   ��پ�T����:��gڽb;i�����\���|�	�*(y��-ӽp�"�k�g�,T����¾!p꾱��<����"�z����3S	����jȾaן���q�iN,��u低����h$�X��*���w��r߽(<��d��Tپ�g��I��O��`���ൿIEͿ��߿���V���쿛\῱)ϿH���R뜿m̀�ПJ�XC��   �   Ty�L%���7i��j	�߾�����hKI��)9���м�HX�,ں����<�D��t~���������U^ɾp�־��۾Zؾ�O̾����Y��
���j�O������Ͻp�����d��HL�����䚽����l�������89��Xt�g*��N���~�ٿ�V�����V��R}��K��n��)�� uۿ�����𚿛u��Q9��   �   B%���׾TO��K�%��ݬ��� ���@�;@D�:��e�� �n���U)߽k��3�?�7Ec�����j���%���Ɋ�����j�j�>�H��>"�� ���U���M�`�ʼ [�@����.l�8�,�p����@,�=Y��ȜھN���Y��Ԏ��b��p�ؿ��������F#��f&�h�#��~�����N��j9ٿ�����;�X��   �   B2�^���8��� ?�a�Ƚ�U�@!�H=�<H`�<�Pm< ��H����5G�1����ӽ.���	��q$�j�)�3�&������	��U�3���4�s��V��QP�@88;��"<0��;�!C�D�Ыڽp�G��ʣ�z���4��v�����ɿQ���V�<f��'.��8�$�;�V8�@�.����ґ���$ɿ�9��_�t��   �   �pB����ǯ���S���߽[.� |9,n�<��=,�
=���< �)<������ �B�_慽jA��n�� r��@໽]���F����e����:��@�ɺh;P<P�<x·<�wP< �4�0�Y��*��)�]�Tܴ��g	��9E�����GD�� �ڿ2������-�>�b7I�V:M��cI��K>�r�-��^�BX��ٿ�ۭ�����   �   ��L�S�)%���`�t��zr:��w:F�<~7-=��8=�1$=Ġ�<p&}< H,��Ā�t?���(���H�$�V��7R���;�`N� 'ƼH�&���;��<�w�<�;=�C�<,>�<� 2�h�h��|�l�Xݿ�b�h9P�bǍ��_����X{
���!��6��H���T��Y� �T���H���6�2� �d�	�6D� ���'����   �   �zP���"���:�e����6�>���:<q�<�u7=��G= c8=jq= /�<Y<l��@���,��.�^g ����w�� ̼��b�������@<,}�<b�=��=��=LÏ<�42���m�.l���p�&�þ"�T��C�������鿤��.N$�r*:��uL���X��;]���X��PL���9�L�#�|�����|u���T���   �   �L�fR�9$����`����:p:� ow:�G�<8-=2�8=�1$=��<�&}< L,��Ā�p?����(�ĤH�&�V��7R���;�HN��&ƼX�&��;@�<�x�<<=|E�<l@�<�1��h��{��l�^ܿ�ja�s8P��ƍ��^�����z
���!�.�6��H���T��Y��T���H�2�6��� �ֵ	�JC�?�������   �   oB����9ů�:�S��߽�V.� J9�q�<�=��
=���<8�)< �������B�a慽sA��s�� r��>໽K���0�����e���9��@�ɺ�>P<t!�<�ŷ<�P<��4���Y�u'����]�uڴ��f	��7E�l����B��H�ڿ��f��\�-�J>��5I�j8M��aI�,J>���-��]�2W�P�ٿrڭ�����   �   �
2����������?�ܖȽ�O�@��DB�<Dc�<�Tm<��������5G�1����ӽ0���	��q$�h�)�.�&������	�yU����s��U�hMP� P8;��"<p��;C���C��ڽ�G�]ȣ������4��}v�� ��[�ɿH��U�2d�\%.�j 8���;��S8� �.���������	ɿ�7��*�t��   �   V"�I�׾`L��F�%�Hج����ζ����;�~�:8�e�H� �J���B)߽j��5�?�?Ec�����j���%���Ɋ�����Z�j�$�H��>"�J ��/U��¢M���ʼ Q��j�� l���,������<,�0V��l�ھK�
�Y�3Ҏ�_��ӂؿ���������C#�d&���#�@|�*���J���5ٿ����}���`�X��   �   *v�� ��P1i�0f	�����<���7I��9���м�GX��ٺ����0�D��t~���������W^ɾt�־��۾Zؾ�O̾���sY������3�O�r��A�Ͻ������\���@��~��qޚ�&�(�l�bz������49�bSt�'��`�����ٿ�Q��؞�n��\z��H��k��$���pۿ�󻿑횿?u��M9��   �   <�پ!P��.�:�_ڽj/i��������:�	�8&y�D-ӽH�"�X�g�'T����¾#p꾴��<����"�z����.S	�����iȾEן�h�q�N,��t�2�d$���编��v�w��i߽n!<�@`���پVc�iI�I��\��ܵ�0@ͿB�߿��,P����Wῒ$Ͽ����Q眿ɀ�Z�J�?��   �   ~����c��h�)���<��0��f���~�wJ׽��)��y����N��n���&���>���Q�&w^�&'c�s�_�\T���A�-�)�d���c澜	����� 21��_㽦1���w)������B��ɦ�V���Ya��,��6���ZK�v�x�LN��񳥿`�����¿CϿ�w���y�����|���M��� �$���   �   �|�i�&��ͽ��q����d8���j�M;ǽ>I"�hFw����>��I��I�>�7�a�"����⌿:씿�엿t������$��`Oe�S"B��������������|�J�&�ͽ��q�Ċ�7���j��6ǽ�E"�cAw�M������|����>�H�a�쉀�V����锿'ꗿᕕ�%�����:Ke��B�����~��ث���   �   |-1�Y�d-��Xs)�~����B��̦����]a�s/���	��qK�-�x�sP��Z����
������¿ҿ��y��K|��� ��|��M��� �P�ﾗ���c��k����<�<�40��b�6�~��D׽F�)�D�y������྇����&���>���Q��r^��"c���_�T���A���)�Q���^澆���
���   �   <m��鋽�]$����P��h�w��l߽5$<�Xb���	پXe�I�FL��^��V޵��BͿ��߿���S����Y�.'Ͽ���a霿�ʀ�3�J�PA���پ�R��a�:�cڽZ3i�̻���z��6�	��y�L&ӽ��"�&g�AP��&�¾�j꾎 �9�n��"�Vv����O	�־��dȾ$ӟ���q��H,��   �   ������R��<��މ��������l�v|��"���69��Ut��(��A���)�ٿQT��2������{�J�Zm��'���rۿ����Ju��O9��w� #���4i�?h	�7��������0I��
9���м�<X�gҺ����"�D��m~�;~��
��Xɾ��־�۾KTؾ$J̾y���T�����ΦO�N��G�Ͻ�   �   ��ʼ 8� L���l�8�,�\���Y>,�tW��S�ھqL�ռY�Zӎ��`����ؿ������`��<E#��e&�
�#��}�^���L���7ٿK���̩��v�X��#���׾�M��F�%��ڬ�����ȶ���; 0�:@�e�(w ����7 ߽���ړ?�>c�����f���!���Ŋ������j���H��8"����xM����M��   �   `�8;H�"<���;C�N D�_�ڽ-�G�eɣ�W����4�v������ɿ����U�*e�x&.��8��;��T8�&�.���������ɿ�8���t�/2��������|?���Ƚ�Q����HF�<�j�<�km< �}�<x�� )G��)���ӽ8�����k$���)�d�&�M��y�	�OL� y��(�s��J�@+P��   �   �)�<d˷<h�P<�}4��Y�I(��q�]�#۴�g	��8E�ꌆ�iC���ڿ�������-�>�n6I�`9M��bI�K>���-�4^��W�N�ٿFۭ����%pB�q��MƯ���S�>�߽zX.� �9�s�<\�=p�
=��<�)<Px���� �B�-����:��W����j��
ٻ�d���ő��<�e�� )�� �Ⱥ�TP<�   �   D>=�H�<�B�<��1�֜h��{��l��ܿ��a��8P��ƍ�4_����z
�@�!���6�\�H�,�T�Y���T�(�H���6��� �,�	��C俼��������L��R��$����`��q:� Rw:hH�< 9-=��8=�3$=��<�5}< �'�$����3����(��H�6�V� 1R��;�H�xƼ��&��=�;,�<`~�<�   �   �=��<P�:<�K�� ���%�����b?꾗40��z����o�ۿ����%�B�`�]���u��?��|4���;����u��i]�T$A��#����=ٿɍ��0w��-�>�便Ό�
��M[��p�U�8��<�
=��)=E=���<�qK<�n�(Ӡ����O;��D[��h�ޘb��xI����TcӼ�0� j�;͕<+�<�   �   ���<@��<h
$<����!��?�!�UՎ������,��\v��զ��ؿ����N"���>���Y�q������d��j���6�p�UY�`�=��U!��n��տoդ���r�n�)�Հ�x�����E���P�X�l1�<�z=��=�>=�)�<��n;h�e�"g��LB�2zv�F������e���j��\�V������� ���Ȁ6<�x�<�   �   ͂<� �<���;���ի��� �&�����ؾ��#��i�a|���{Ϳ �BF�d�4���M��c���q���v���q��Kc���M�Fc4����������˿�圿ƪf��!�<Ծd2��Z�� s��p�e��b<H��<��<�0k<`���;��<��5��2���x�ֽ���߿��+���F޽
3���X����Z�� ��y0� A�;�   �   �i��@�;�~��9��b����Y	�,_s���ľ�$�ٜU��j�������뿠��.�%���;� oN��[�x�_� �[��O��h<��%�Z���;��!��Uc���S��%��'��Xl��+��7n����`	�;`.(<��;x�|���%��֏�0 ѽ��I%� [<���K�ҘQ��M�cr@�� +��u�#��{���zH�8�¼�   �   Z���@��Hq�|�ټ�`q��&�IzS��٫����@<�
����i4ҿ,���o��s&�P6�z�@���D��;A�.7��d'�+����tҿ(৿O���;��z������M��d��X�຤�@�����G������1s�Дƽ*��E�>�5�l����Р��C��������ɧ�I���,>��#Gt�`�F��F�W�׽ R���   �   �E��:�K�6]����Č[�P�ɽsr0�b�tܾ
����[��1��!"����ڿ���fk��j�j%�vK(���%��k�����O �gܿ���B�����[�N��.۾�K���,���� �G��1�,�ټ��0�KU��F�����2��s�8H���Z��$ھ��/� ����z�ڧ����ݾ����䟾�8|�x�;�Й��   �   y��J��i�R�1�ƒO����%T���f�P,��B�"R4�bLn����������տ����>�	��|��e
�~���S�(3׿�H��?З���o��15��c������e�TA��y���bA�d� �R�T�Jt���@�)K��ۍ�������]�RG!���1���<�L�@�=�^�3�"�#��%�ﾕ���T��n�R��   �   �'Y����Y9���Yq�<R��+���^ٽ��0�����l�ʾc���=�ݵp��̒�.��"q¿�Կi�߿����i�տmxĿ #��k���Y�s��*?�dR�M�̾G����{1���ؽ�ǅ���I���e�5����!
� S��B����ϾD���,'��F��qb���x�����6�������z�Ae�m�I��"*���	��dԾ����   �   +5��H&M����%{��x�e��(d������, ���I������qվM���m8�Ԙb�󛅿=����ѥ��������ԯ�G0���P��;g����e�D>;�J���ؾ?2��>"M�j��wx��V�e��+d�H����/ �X�I�״��Evվ&��q8��b�X���曗��ԥ��������ׯ�3��yS���i����e��A;�����ؾ�   �   ��̾�����~1���ؽ�ȅ���I���e�����
��S��>���ϾD��@)'��F�mb���x�s����3��Q����z��<e�h�I�@*��	�e`ԾN����"Y��� 5���Uq�BR��-��cٽ��0�f���(�ʾ���!=�Ĺp�Jϒ����	t¿�Կ��߿Z��=��w�տ={Ŀ�%��������s��-?��T��   �   :e�Y����e�)C�.{���aA�� � �T��m��^<�K��׍�������{��C!���1�5�<��@�u�=�J�3�e�#�������	��Q����R�q�#E��Zi���1���O�%"���V�v�f�5/��D��T4��On����������տ�������	�J~�2g
����V�5׿�J��җ���o�45��   �   �O�1۾sM��͔,�����(�G�8+�P�ټ��0�<N��������2�(s��C���U��6ھ���η ����v������ݾ����#���i1|�ŷ;�z���?����K�XX�.����[�+�ɽ
u0�h� wܾ��l�[��3��($����ڿۥ���l��l�2%�DM(�h�%�Xm����P ��ܿ�������@�[��   �   J;��{�Y����M�df㽞�X�����@�����G�L����#s�ƽ�����>�r�l�,�����L��������ħ����9���?t���F�MA���׽�K�����84���q�T�ټ^cq��)��|S��۫�U���A<�KÀ� ��M6ҿK.���p�Nu&��6�@�@�|�D�H=A��7�"f'�0,����vҿv᧿P���   �   '�S��&�)���l��,��8n���� $�;�C(<�[;Hs|�,�%��Ώ���н�z�C%��T<��K��Q�$�M��k@���*��p�+��{���H��¼ 5���;�]��9�������Z	�jas���ľ�%���U��k��8	��<�뿖��R�%��;��pN�`[��_���[�>O��i<� &�&��=��"��%d���   �   ��f��!��<Ծ�2�����0s��p�e��b<X��<���<�Jk<�>�ܹ��R~<��.������^�ֽC��J���ñ��>޽�+��R����Z�8 �8\0��n�;PՂ<��<��;�������������ؾ�#�J�i�2}���|Ϳ� � G�D�4�ʯM��c��q�>�v���q��Lc���M��c4�$��ݍ����˿朿�   �   ��r���)��ྜྷ�����+���0�X�4�<�|=R�=8B=2�<��n;@�e��`�HEB�frv�4�����a��4g��n�V����$���0l����6<�}�<��<T��<0$<䪱������!��Վ���徆�,��]v�;֦�+ؿV��`O"��>���Y��q�惀�4e��������p��UY���=��U!��n�[�տ�դ��   �   �w��-���侌Ό�����Z����U�H��< =�)=lE=���< sK<`n��Ҡ�ܢ��O;��D[���h�ؘb��xI�����cӼ��0�`h�;�̕<l*�<��=��<`�:<,M�����%������?��40�X�z�%�����ۿ���%�&B�r�]���u��?��}4���;����u��i]�B$A���#�Ќ��=ٿ�����   �   ��r���)���������佈���X�,6�<p}=��=tB=d2�<@�n;8�e��`�PEB�jrv�9�����a��2g��`�V�n������pj����6<�~�<<��<���<0$<\����
����!�"Վ�}�徵�,�l\v��զ�BؿƇ��N"�2�>���Y��q�7���d�������p�zTY���=�RU!�tn�|�տ�Ԥ��   �   ��f�!��:Ծm1������p����e��b<���<T��<�Lk<@;�����F~<��.������n�ֽL��W���ʱ��>޽�+���Q��H�Z�� � Z0��t�;`ׂ< 	�<��;$���d������������ؾa�#�,�i��{���zͿ� ��E���4�حM��c�r�q���v���q��Jc���M�nb4���ы����˿�䜿�   �   Q�S��$�(&���l�*��1n�����:�;�J(< l;�p|�޿%��Ώ���н�z�C%��T<���K��Q�$�M��k@���*��p�����z���H��¼�)���.; *�D0�����X	�T]s���ľ�#���U��i�����H�����.�%�x�;��mN�0[���_�h�[�^O�bg<���%�n��@:뿤 ��Kb���   �   �;�jy������M�)`�r�X� ��� ���H�G�����#s���ƽ�����>�|�l�2�����Q��������ħ����9���?t���F�'A�w�׽K��4�� /����p���ټ�Zq�"#��wS�%ث����~><����=���2ҿ*��Tn�rr&��6�ĩ@��D��9A��7�Nc'��)�� ��sҿ�ާ��M���   �   L��+۾�I����,����H�G���yټ��0��M��~�����2� s��C���U��=ھ���ҷ ����v�~�����ݾ������>1|���;�*���>����K�0T����N�[�%�ɽ�o0������qܾN��r�[�o0��R ��w�ڿ�����i�di��%��I(��%�j�"��NN �ܿ�������[�[��   �   ~a����2�e�>�Qt���XA�� �^�T��l��<��K��׍�������{��C!���1�8�<��@�v�=�J�3�c�#���t���	���P����R����C��*i�P�1�b�O���XQ���f��)��|	��O4�^In�Ō��^���jտ������	��z��c
�ڼ��P�o0׿)F��6Η���o�/5��   �   ��̾s����w1�/�ؽ0��I��e�K���t
�KS��>���ϾC��B)'��F�mb���x�v����3��Q����z�~<e�d�I�:*��	�J`Ծ)���"Y�o��3���Oq�2R��&��YٽM�0�A����ʾ#��=�F�p��ʒ����_n¿�Կ;�߿���Ɉ�L�տ�uĿ_ �����p�s��'?��O��   �   �.��M����;r��n�e�� d�����+ �8�I�o����qվK���m8�ؘb�����A����ѥ� �������ԯ�G0���P��9g����e�<>;�?����ؾ2���!M�����u���e�jd�*���T) � �I�~����mվ���Dj8��b���������2ϥ�3�������ѯ�k-��8N���d����e��:;�j����ؾ�   �   �Y���� .��Jq��R�(��x\ٽN�0�����W�ʾ^���=�ߵp��̒�1��'q¿�Կj�߿����i�տmxĿ�"��h���Q�s��*?�WR�&�̾
���{1�W�ؽą���I���e�ꋭ��
�L	S�{;����Ͼt���%'��{F��hb�ѐx����E1������z��7e�8�I��*��	�{[Ծv����   �   ���=��:i�H�1���O����@S��f�/,��:�"R4�bLn����������տ����@�	��|��e
�~���S�'3׿�H��;З���o��15�sc������e�Z@��v���YA� � �~�T�6g��8�hK�ԍ�V����꾶x��?!���1���<���@�%�=�(�3���#�T������M����R��   �   �7��B�K�N�(����[��ɽ�q0�2��sܾ����[��1��""����ڿ"���hk� k�n%�xK(���%��k�����O �eܿ���@�����[�N��.۾�K��)�,�����κG�(��nټ�0�FG�������2��r�`?���P��ھW��~� ����Js�����ݾ�����۟��)|���;�~���   �   ���� ����p�D�ټ�[q��$��yS��٫����@<�����k4ҿ,���o��s&�T6�|�@���D��;A�07��d'�+����tҿ'৿O���;��z����5�M��b�~�X�|���0k��ؗG� ���(s�3�ƽJ��6�>�	�l�����|���n������������읾�5���7t�!�F��;�u�׽D���   �   �� �; ���-��p����X	��^s���ľ�$�ٜU��j�������뿢��0�%���;�"oN��[�x�_��[��O��h<��%�Z���;��!��Sc���S��%��'���l�N+��3n�����L�;8\(<��;�L|��%�dǏ��нvu�H=%�ON<�@�K��Q�^�M�xe@���*�.k����s��L�G� �¼�   �   �<��<�+�;d�������% ������ؾ��#��i�a|���{Ϳ �DF�d�4���M��c���q���v���q��Kc���M�Fc4����������˿�圿êf��!�<ԾD2������q��0�e���b<��<���<Pck<`��0���Js<��(��������ֽ�����f���6޽6$��GK����Z� ��90����;�   �   D��<���<$<襱��
���!�IՎ������,��\v��զ��ؿ����N"���>���Y�q������d��k���6�p�UY�^�=��U!��n��տoդ���r�k�)�̀�j�����������X��6�<|~=��=�D=D9�< ?o;��e��Z��>B�kv�Q����ꓽ�]��Wc��8�V�����뭼�C��П6< ��<�   �   H��<̣�<��;�IK���A�����x���}I�����cb��'h������<��K_�S!���a���ښ�x����՚��A��5р��F^���:��������3��j䌿v{F�e�Ve���T:��@��$�ϼ�	><|��<��=�<`R�< mW;��l��W��fD�T�x�����|��Gz��!聽$TT�Z�G�� �0��Q<t+�<�   �   ��<���<�Me;�L������ >�f������E��@���,��T���P�$�8���Z�h�|��9��fd��E	��k���.��:y|�0Z�X�7�
 �I�1&��)���2C�í��E����6�+=���iѼ�"<�k�<���<,��<(�5<Qջx�ռ`B:�䀽ȅ��`v��o���{���K��w���?N�Ε��tM���;p�<�   �   h�&< �8<�����5�D����J3� ������%\;����س������dI/���N���m�h[��'������ƍ�΃��v�m�"�N���.���\���=��0���v�8��Z��.C��},��Ϧ�t�׼���;��<���< M�;�[����}�{���W�߽�U��s�)0���n����h}��x���V[/��ס�@$���   �   �%j� ��@�+����k����"���������*���s��;��Wֿ<_�x� �0�<�2�W���n���~��H���1�ȅo�j[X��0=�� ����$տo4����q�!)�|�߾8a��N���՚�P�輠=����U:������\Re��綽r�����#��D���]��n��`u���p�Bla���H��)��U�i-Ľ_
������   �   0�N��L���RȼX��2�����w��ƾ=�n>W�����V���P��R?�VL'���=���P��]��{b�vI^�<�Q���>�d(�����!n���%��V���#+ľ�2r�6
��0���L�䱜��ż�6����{����I,��Fa�E�����������Q���F�ž�¾�ö�Ѥ�y썾_Vh��m3�rF�MA���   �   Sͽ�Ƃ�>�6�V�8���ӻ󽑅O����y���B7���z�]�IͿ�i����ܠ"���1�H<���?�ؾ<�h�2���#��)�_���3οSW��E�z�L�6�����p���v=L�d��k3���"'�m#�Jp��U��'\��JT�8m��`����!ھ����%J���Q����A���/��<޾S����\��Ǡ[����   �   �_)�U�޽孓�*�i�����{̽�'��׆�`ξb��UtN�Uᇿ��t�ο�"���j��#�$-����&��	��_���пc^��ǫ���LO�$���
ξ�Q���?&�6�ǽ	��t�[����Mս1�#��lo�>w��q�ؾ\���!��9�n�K�u�W��O\�r�X��VM�
5;���#�ܻ	��Cݾ�]���"v��   �   6c}�H)���ܽ4㘽�����Ъ�TT��P�-��7N�q#��xX�	G��D=ÿ	:ܿ������� �{���m��1S޿�Nſ赨����grZ�ul$�P������@Q�:�਽
E��j9��ϧֽkp%�h+x��'��$P��H�W�?�p#c�XA���������$���kP��K���=���<f���B���)m��Mw���   �   �p���p����l�ɽ	.��-t���Kǽ����m�]4�������&%�qBS��_���(��!H��p(���wƿ<Kʿ�?ǿ�����������$�U�*?'�����Hm��ep�տ�W�ɽ]-���u��Pǽ���	m�8������ *%�iFS�Rb���+��K���+��6{ƿ�NʿBCǿ0�������������U�%B'�D����   �   ��k����Q��]ᨽD��#6����ֽ�k%�%x�E#���J�E�H�?��c��>��Ѧ��%���/����M�����������f���B����h��js���]}�j{)��ܽ�������� Ӫ��V�'�P�2"��sR�B #�||X�:I����3@ÿI=ܿ��s���]� �������XV޿oQſU���
����uZ��n$��   �   ��Vξ�S���A&��ǽ�����[�ߑ��!ս�#��eo��r����ؾ�X���!��9�ǪK���W��J\���X�dRM��0;��#���	�h>ݾ�Y��Lv�[)��޽!����i�'���V!̽��'��ن��ξ���SwN�9ㇿM��$�ο�%�L��J��%�(/�������	�}b�t�пw`��w���lOO��   �   6�6�7���:����?L�]��}3��t'��e#�,
p��M���V��CT��h��;����ھʹ���F��	�.M�������#)��f޾[����X��U�[����Kͽ������6���8�����z�O��	�������7���z�>�LͿ<l��b���"���1�h<�&�?���<�R�2���#�<+�����5ο�X����z��   �   �V���,ľ�4r�1
�N1���J�`���H�ż� 6�����M���ZC,�?a�ޛ������&���������ž¾����)̤�0荾Oh��g3��A��9����N�x>��Kȼ������<���	w�G�ƾ�>��@W�c������n��@��M'���=���P�>�]�~b��K^�&�Q�\�>��(���a#�0p���&���   �   �q�)�Η߾b�� ��֚�D��  ���JW:���|��De��޶�������#�D���]�V�n�(Yu��p��da��H� �)��P�%Ľ������Hj�p䪻��+���m�� �"�F������T�*���s�=���ֿ&`��� ���<�ԷW���n���~��I���3���o��\X��1=�� ���&տY5���   �   �����8�i[���C���},��Ϧ�P�׼��;��<�ć< ��; �Z������}�����߽Q��n�P+�\�j�l��v��/����P/� ǡ� Y����&<آ8<@y��B6�����L3�"�������7];�����س�������BJ/���N���m�(\����������ƍ�{�����m���N���.�j�(�濃>���   �   X���rC����E���6�=���gѼ��"<�o�<D��<���<x6<�$ջ��ռ�::����e����q��� ��w���G�������8N�܏��`M�P!�;P�<(��< ��<@Re;�M�o����!>��f��y�s�E�A��*-���T���P���8�� [�.�|�:���d���	��pk��2/���y|��0Z���7�D ���o&���   �   K䌿C{F�>�e���T:�Y@����ϼ�><T��<V�=��<S�< sW;��l�\W��fD��x�憍� |��Bz��*聽<TT���pG����0���Q<�*�<���<��<�;���K��[�A�橨����~I�Ƿ���b��Ph������<��K_�_!���a���ښ�x����՚��A��*р��F^���:���������3���   �   �����C�K���D����6��;��ddѼ��"<\q�<$��<��<�6<`$ջ��ռ;:����h����q��� ��
w���G�������8N�Ə�8`M�0#�;�<D��<���< ge;�K�����p >��e������E�x@��Z,���S��RP���8�l�Z���|�R9���c������j��m.��~x|��/Z�ޱ7����
�%���   �   ����m�8�Y��B��i{,�ͦ�L�׼p�;l�<(Ƈ<���;@�Z������}�����߽$Q�o�Z+�b�j�h��	v������P/�<ơ� A����&<�8<�-���2������I3�x������x[;�S��d׳��迖���H/���N�d�m��Z��c�����Qō����4�m��N�,�.�>�K��=���   �   �q��)���߾�_��4��4Қ���輠����W:h��<���Ce��޶�������#�D���]�`�n�4Yu�
�p� ea��H���)�rP��$Ľd������j��Ҫ��+�ؔ�i���"�����\����*�F�s��:��"ֿ|^��� ���<���W�4�n���~��G���/��o��YX�:/=�� ��g#տF3���   �   �V�>��(ľ4/r��
��,���D����Ԫż��5�����"���RC,�	?a�䛊�����/���������ž¾����'̤�*荾�Nh�wg3�|A�s9����N�09���Bȼ|��������ew�@�ƾ�;��<W�ҕ��ܛ��|��2>��J'�*�=���P��]��yb�LG^�<�Q���>��(������
m��S$���   �   �6�"��������9L�ŀ콆.��('�b#��p�&M���V��CT��h��?����ھҹ���F��	�2M�û����")��a޾P����X�� �[���Kͽd���N�6��y8����.�󽙂O��������O 7���z����GͿ!g��f�.�"���1�6<���?���<�n�2�8�#�@(������0ο|U��P�z��   �   ���:ξ`O��	<&�G~ǽ���"�[������սȩ#��eo��r����ؾ�X���!��9�˪K���W��J\���X�fRM��0;�	�#���	�X>ݾ�Y��v��Z)���޽꧓�Dyi�񰅽r̽��'��Ն�uξc���qN��߇������ο������
��!�$+����F�2	��\�K�п\��穈��IO��   �   �뾤����Q���
ڨ�H?��3���ֽrk%��$x�2#���J�E�J�?��c��>��զ��)���1����M�����������f���B�����g��Hs��%]}��z)���ܽ�ݘ�����}˪�7Q�~P�a��fJ��#��uX�E���릿�:ÿ�6ܿ���3����� ��������O޿�KſS���Ѧ���nZ��i$��   �   ni���p�z��y�ɽZ'���o��.Iǽ���0m�A4�������&%�rBS��_���(��%H��t(���wƿ>Kʿ�?ǿ������������U�"?'�����m���p���h�ɽ�(���n���Eǽ�����l��0��
~���#%��>S��]��o&��IE��Y%���tƿ�Gʿ�<ǿى�������왿E���&�U��;'������   �   �V}�dv)�O�ܽ�ژ�膇��̪�(S�g�P����"N�m#��xX�G��G=ÿ:ܿ!������� �|���m��2S޿�Nſ嵨� ���^rZ�kl$�,�뾘���uQ���+ܨ�?���0��3�ֽ�g%�-x�T���E�[B�r�?�Pc�><�����G���A����J��������� f��B�K���b��o���   �   �U)���޽q����ti�����T̽�'�Z׆�<ξ]��StN�Wᇿ��w�ο�"���l��#�$-����&��	��_���пa^��ī���LO���j
ξ�Q���>&��ǽ#����[�	����ս6�#�v_o��n����ؾ�U��!�l9�>�K���W��E\���X��MM�,;�,�#�O�	��8ݾ5U��2v��   �   1Cͽﺂ�t�6��v8���O��фO�~��c���A7���z�_�IͿ�i����ܠ"���1�L<���?�ھ<�h�2���#��)�_���3οRW��A�z�C�6�_���1����<L�̃�n/��2'�L\#��o�F���Q�w=T��d��X����ھN����B��VI�����d"��`�ݾ'���TT��H�[�@���   �   &�N��(���8ȼj��4�����vw��ƾ =�n>W�����Y���S��R?�ZL'���=���P��]��{b�xI^�:�Q���>�d(�����!n���%�� V����*ľ�1r�>
��-���C�D�����ż�5�H�������^=,��7a���������𥴾(����žj ¾.���5Ǥ��㍾eGh�(a3�f<��1���   �   8�i�@���~+�z���i����"�у�������*���s��;��[ֿ>_�z� �2�<�4�W���n���~��H���1�ȅo�j[X��0=�� ����$տo4����q�)�`�߾a�����wӚ�P���� �X:�s��伊6e�nֶ�����#��D�v�]���n�kQu�Z�p��]a�G�H��)�8K�Ľ���l���   �   x�&<X�8< ����1�⵳�pJ3��������%\;����س������fI/���N���m�i[��(������ƍ�σ��v�m�"�N���.���]���=��/���s�8�{Z��C���|,�:Φ��׼p(�; �<Dχ<@��;8�Z�x��,�}��汽��߽�L�Rj��&��
��e��}轂n�������E/�$���@\���   �   ���<Џ�< }e;�J������ >��e������E��@���,��T���P�$�8���Z�j�|��9��fd��D	��k���.��:y|�0Z�X�7�
 �H�0&��)���0C�����E����6��<���eѼ��"<�s�<��<���< 6< �Ի�ռH4:�C܀�D}��hm��Q����r��VC�������1N�b��xJM�PG�;L�<�   �   @��<�E�< @9$��ܽ��X�������>�]�A���bpҿd��(�)���O��5y��t�������ѯ�� �� ̯��q���&��=x���N� �(�����п�󚿶$[�5~�{x���R�^�н6x��*�;^�<��<���<��]< -d�H鸼B"*���o�Fٓ��,���O��{����n��z�|���9���ܼ��p<0�<�   �   tܫ<T�<��ɺ�g$�rzؽ�T�fn�����,�Y�0ٙ���ο����&�t�K��"t�D���ٟ��˫�����ѫ��Ο����n]s�&�J���%�*���3Ϳ�`���TW�N�������N��cͽ�+� hi;�Ե<(��<��<�k�;�9g��F���e�Kn��}"��*M̽�Խs�νpռ�l���	v��"���� \����g<�   �   p�;07�;��㻺�&��rν��H��(����	�-QN����C�Ŀ�6�����A���e�@N���W���X���O���z���~��X���e���@��������Ezÿ�ߐ��>L�.����ocC�[Ľ.\�@��EB<�m0<�q��V����?�����vϽ� ��l��l!�h^&���"�T�����ؽح���3T��!ۼ0ػ�   �    ˪�@�4��,����-����$7�yX��2��y<�������)�j��p�0�x�P�hdp����e_���ؒ�Ɲ��TB��� q�f,Q�B�0�̰��X鿘+��;��G�:��?����t02�g������XF��˻�����5��#{ս·�H�9�s�\��x����)���&R����{���`�tZ>�b��Aགྷ��Ƶ.��   �   v�v�@��*���>�u����M!�X����ܾ*�%���l�ޠ�U�пH!�����8��Q��#h�ew�}�Zx��i�^�R���8�h�<@��п�}����k���$�
ھ"����^�����P.�l��.�l�b��l��A~�bC�N}����������Ⱦ�3־~۾�"׾F�ʾQ߶����\v���H�"*��$Ž�   �   {v�yG��`�\���^����.k
�9h�	����u� �I�Eቿ�ʳ����Vl�P��(�2��/D�T�O�\T�^�P�,8E���3�����Q��s&��4�I�_���V��
�e�~�TC��d�P�zUM�d������(���n�jC���7ɾN?����#�>�#��$'��?$��;�[��������̾����� u��_.��   �   q/>�����嫽�I��jܜ����=��T�����K%���c��[������)��������d"�<m+�x�.���+�fU#�����M/��ü�s���Cd��%�����蕾�;� �SG��ZɄ��U��������9�DL��S���O�� �ɵ2�DLL���`��m��r�'{n�-�a�#N�V�4�"�$����Ȼ�����   �   �$���}>�S���j㱽���s�Žh'�`�i�{>��P���?4��n���\.��p�տa$�\��i
�j��
��#�|���׿޺��"���Gp��^5�4������Oj�����1Ľ~v�����D����#;�<���,Ež&P���+� �S��Mz��4�������Y��Y����ݤ�֕���b��j�|�<(V���-���pȾ�   �   ��ľ@�����/�L�8!������o彡.�豄�d�¾c��v�6���h��_���$��M����+ο�Nٿubݿ{�ٿ�cϿz��筨�wÏ�$Ik�E[8���	���ľ����P�/��H�| ��Ɖ��Ot�w	.�δ��|�¾"����6�L i�Zb���'������!/ο,Rٿfݿڿ^gϿ)}�������ŏ�4Mk��^8�0�	��   �   >��d����Rj�	��'3Ľtu���������;������@ž&M���+���S�Hz��1������dV��"���xڤ�֒���_��{�|��#V�a�-�	�+Ⱦ�!��Vy>�����౽�����Ž*���i��A������B4�јn���(1����տ�'�^��k
�t��
��%�����׿�����$��$Kp��a5��   �   �%�����ꕾ<�;����F���Ƅ��P������5|9��H��v���=������2��GL���`���m�Hzr��un�(�a�lN�>�4����_���gĻ�b��m*>�����᫽�G��ݜ�)���=�W����侔M%���c��]������⿆�����f"�zo+���.���+�rW#������2�1Ƽ�I���Fd��   �   .�I�����X��f�e�+�nC����P��MM�U���J��J�(�?�n��>��?2ɾ�8�n~����#�� '�z;$��7����-����̾�����t�EZ.��n�:B��V�\� �^�4����l
�:<h������w���I��≿�̳�E���m��,�2�F2D���O��^T�ʘP�`:E���3�r��p����6(�������   �   ��k�F�$��ھ;����_�?�����-�4�����b�Zd���x�zC�}�����*��%�Ⱦ�-־9۾s׾t�ʾ�ٶ�a���Zr��i�H��$��Žܸv�������&�>������O!�寉��ܾ��%���l��ߠ�:�пp"�P �f8�( R�&h��gw��}��x�i�F�R�*�8�Di�:A���п�~���   �   ���^�:�8A���Ú�`12�׺��D��HF�`�˻4������..���qս����9���\��x�ۈ�������M��Ģ{�?�`��S>�ݲ��7�?�����.�����p�4�P'��İ-�k���7��Y��N���z<��'���*�l����0��P�Vfp�����`��<ڒ���`C���q��-Q�P�0����'Z鿘,���   �   i���p?L���g�� dC��Ľ[�����UB<��0< w��8B����?�S��rnϽ�� ��g�dg!�Y&���"�j�����׽����f(T�Hۼp�׻��;�P�;@��:�&��sνG�H�*��w�	�WRN����@�Ŀ�7��ԭ��A��e�O���X���Y��{P���{������X��"�e�`�@�0��q����zÿ�   �   �`���TW�x��-����N��cͽ�*�`�i;tٵ<h��<졝<p��;�!g��?���e��i�����)H̽�Խ��ν�м�(���$v���"����� ����g<��<��< �ɺ�h$�q{ؽ��T�o������Y��ٙ���οR���&�
 L��#t��D��ڟ�&̫�B��aҫ��Ο�5���]s���J��%�\���3Ϳ�   �   ��$[�
~�9x����R�غнlw�@0�; _�<���<���<X�]< 'd��踼�!*�n�o�-ٓ��,���O��t����n����|���9���ܼx�8<`/�<���<�D�< x?9�$�ܽ�X�����D��x�]�e����pҿz��@�)���O��5y��t�������ѯ�� ��̯��q���&���<x���N��(����j�п�   �   4`���SW����A��x�N�bͽ�(���i;�ڵ<T��<���<���;h!g��?���e��i�����7H̽�Խ��ν�м�)���"v���"����� \�8�g<�<��< �ɺ�f$��yؽ��T�)n��c���Y��ؙ���οč�`�&��K�z"t�'D��(ٟ�#˫�9��`ѫ�Ο�n���\s���J�h�%�҉� 3Ϳ�   �   )ߐ��=L�Y�����aC��ĽBW�����[B<�0< f���A����?�O��{nϽ�� ��g�ng!�$Y&���"�p�����׽ꦡ�2(T�`ۼ@�׻�;�]�;P��B�&��pν��H�C(���	�pPN�f����Ŀ�5��x��0A���e��M���V���W���N���y���}��WW���e���@����d���Ryÿ�   �   ?����:��=��t���..2�������;F�0�˻�݁��� .��{qս����9�
�\��x�∅������M��̢{�?�`��S>�β��7�����ʩ.����H{4�$ ��H�-�!��|7�ZW������w<�J����'꿔��\�0��P��bp����8^���ג�����:A���p��*Q�
�0�ү�MW�U*���   �   ��k�2�$��ھT����[�R�����-�L�⼺�$�b��c���x�qC� }�����2��.�Ⱦ�-־B۾z׾{�ʾڶ�_���Tr��R�H��$�SŽ(�v�ԩ�����}>�Ȉ���K!�쬉��ܾ��%���l��ܠ���пH ���� 8�0�Q�d!h��bw�j}���w�vi�V�R���8��f�?��п2|���   �   ��I�����S��"�e�
{�>����P��IM��������(�(�n��>��@2ɾ�8�r~����#�� '�;$��7����)����̾���d�t� Z.��m��@����\���^������h
��5h�Ά��pt���I��߉��ȳ���� k����B�2��-D���O��YT��P��5E���3�������p$���퉿�   �   q�%���*敾��;��潉A��AÄ��N�������{9�mH��m���>������2��GL���`���m�Ozr��un�,�a�lN�<�4����S���TĻ�?���)>�����c߫�^D��tל����_=�_R��ь��H%�ׄc��Y��B���v��D�(���b"�k+�6�.���+�LS#���d �d,�u���i	���@d��   �   ڇ�����Ij���6+ĽNp���������2;�����u@ž#M���+���S��Hz��1������gV��%���zڤ�ؒ���_��z�|��#V�[�-���Ⱦ�!���x>�����nݱ�v��ڻŽ
$���i�n;��9��=4�Z�n�n�+��m�տ� ��Z��g
�b��
�"���򿅿׿��� ���Cp��[5��   �   ��ľ������/�DA���O����l彾.�����E�¾\��v�6���h��_���$��Q����+ο�Nٿybݿ�ٿ�cϿz��譨�wÏ�!Ik�@[8���	���ľn���V�/��E罨��o���]i�.� �����¾ߡ�8�6���h�e]���!��6���M(οKٿ�^ݿ��ٿ|`Ͽ�v�����������Dk��W8���	��   �   =���s>�����ڱ����e�Ž(&���i�I>��D���?4��n���_.��r�տe$�\��i
�l��
��#�}���׿޺��}"���Gp��^5�"��P���JNj�����-Ľ#p���������;���7<ž\J�J�+���S��Cz�8/������GS���~��Pפ�̏��&]��^�|��V���-���nȾ�   �   |$>������ګ��A��+ל���齺=�`T��ۏ�K%���c��[������+��������d"�>m+�x�.���+�fU#�����M/��ü�q���Cd���%���侅蕾ޫ;���B��~���_J�������v9��D���~���������2�CL���`�^�m��tr��pn��a��N��4����C���y�������   �   Fe��:��D�\�l�^�㛣��i
�D8h�҈���u���I�Gቿ�ʳ����Xl�P��*�2� 0D�V�O�\T�`�P�,8E���3�����P��q&��3�I�O��cV��0�e��|�?����P�tCM�Ҏ��ȥ���(�&�n�L:���,ɾr2��z���#�P'�Q7$��3����{��o�̾V~����t�;T.��   �   r�v����V��J{>�@����L!����iܾ$�%���l�ޠ�X�пJ!�����8��Q��#h�ew�}�\x��i�^�R���8�h�<@��п�}����k���$��	ھұ���]�������-��������b�\��ns��C�}�/��y��l�Ⱦ�'־۾R׾��ʾ�Զ�����.n��l�H�3��Ž�   �   ���b4����̩-����p7�FX����y<�������)�l��p�0�z�P�jdp����f_���ؒ�Ɲ��UB��� q�f,Q�D�0�ΰ��X鿙+��;��A�:��?�����/2������1F�0�˻�́�{��&���hս�|�N�9�֫\�/�x��������I����{�Ҧ`�YM>���0.�9򕽦�.��   �   �I�;�~�; ��4�&�
qν��H��(����	�,QN����E�Ŀ�6�����A���e�@N���W���X���O���z���~��X���e���@��������Fzÿ�ߐ��>L�&�����bC��	Ľ�W� ��HhB<�0< ����/����?�����fϽ� ��b�Nb!��S&�e�"�x��{�^�׽ǟ��,T���ڼ �׻�   �   �<�<@�ɺ�e$��yؽڻT�Yn�����.�Y�1ٙ���ο�����&�v�K� #t�D���ٟ��˫�����ѫ��Ο����n]s�&�J���%�,���3Ϳ�`���TW�K�����V�N�cͽb)���i;dݵ<���<Ĩ�<ൠ;�g�b9�j�e��e��4��eC̽�Խ��ν̼�����:�u��}"��욼 ����g<�   �   ���<���<�U�o6���*9g�z�ƾ-����j�����I޿}�:4�L�]�����C���E��[�����������/�����㝅���\�6J3����ݿ{���i�2��1ľ��b����VC%����: 5�<l��<0�<h`.<p��߼(�@����c��U��1��X綽+���-��l�M�����P5����;��<�   �   Pʠ< �~<�����6�X����b��þ���ۻf�ӽ��W�ڿ�"�@�0�r�Y��!�������7��r8�������<��_0�������ނ���X�E0��u�:yٿ쿡��e��[�����X^�2T�6�%� ��8V�<���<@�< ��:�Җ��1&�<��sR���bȽ7Qݽ�1�(B߽�̽�����u��d�4�������%�h�K<�   �   ��j;@{�;�c�p,9��m޽�wV�5-��.e�ɷZ�ќ���пRU�(�؜M��nv��ȏ�窡��ʭ����W���š��Ϗ��?v��;M���'����u%Ͽ˙�@JY�M$��뵾UDR��Sֽ
)�Ǽ���<`�;�$��poؼL�X��������~
�(���e-��m2��o.���!�X����h,���"i�T%���
��   �   �nǼP�e�,��R�@��TϽO�C�}���b���G�1ލ�����������4�;�3_��-���������ܞ�y7�������c��$h_��;��W����u꾿�I��;�F��_�P���G�?�Ƚ��1�����X*&�x}���0�D<�����
^��G��l����#����7��NI��4����o�LK�i"��&�NԢ�\�A��   �   nن���,����ܘR�n����,�G�����&"0�2{��T����ܿ��	��&�hD��`�5y����g0���K����y�?a���D�4�&���	���ܿ���f�z��m/���DC��ӳ)�Ӹ�P|E�r�����L�}��̽��L�Q������ť������G־�=価K�]��e�׾��¾ԧ�8㉾TqV�����Խ�   �   B���x��N�r�~�t�����b����w�ȏž�U�
CV��/���e������q���'�nP>�RQQ�P<^���b�$�^��R��?��U(����ew�4���~;���V���[�ľ@�u��Z�������i��If������l��d#6�45��Ok��H�־�1�����$�X.�w�1�Lx.� �$�v��;d��jپ�ެ�����_:��   �   �2K��A��C���ٖ�i���e���ZeJ��[��[�f�/�Y�q��e��p�ƿ���"��f���i,��6���9�4~6��-�R����y񿥓ǿ�ߞ�"r���/�E^�&��:ZI�S����������.�p�G��⏾68ž�� ����;<>��?Y���n�FT|�X��� �|�C�o��Z��?��J!������ǾM����   �   �b���K������������
ֽ\H �	z�3"��L
�h�?�uq}��'���.¿���Vk��&!����A������U �#��F<ÿ������~�S�@���
�豾� xz��) �7�ԽN���ѽ���I����>�Ҿ"#�&�6�5Ba�,�����.���$���b���~���)���fׅ��b��v8�+e�[�Ծ�   �   5{Ѿ�쎾4<�ȁ��)������{��r�:� �оޗ��IB�\�w�8)��)H��QEȿ�WڿP�忥)��s�o*ۿ�Iɿ5T�����T?y���C�f��TwѾ�鎾�0<�.~��V��m���2	���:�1�+оƚ��MB��w��+��=K���Hȿ][ڿ"濃-꿧w�	.ۿ2Mɿ)W��� ���Cy��C����   �   ��
�봾��{z�
, ���Խ>��$ν�*}��I�^���R�Ҿ��5�6��=a�z����햿���i!���_��l{��Ư��@����ԅ���b��r8�2b�԰Ծ�_����K����������`ֽ,K ��z��%���N
���?��u}�0*���1¿��o��0#�B�� D�0����lW �Z��?ÿ=���V�~�A�@��   �   ��/�za�?���\I�i��s�U|������*���G��ޏ�3žd� �����7>��:Y�4�n��N|�����n�|���o�>�Z���?�
G!����Ǿ�����-K��=�;?��!ؖ���������hJ�_^���^��/�ʞq��g���ƿ�����r���k,�!6�<�9���6�,-�H��ȋ�W��ǿ�ឿ
%r��   �   ,V���u�ľ��u��[�܉����i��Af������c��@6�:1��Wf��J�־;.�О�M$��.���1��s.���$�����`��dپڬ�^����Y:����s���r�j�t�!���4����w�l�ž�W��EV�Q1���g��9��Zs�z�'��R>��SQ�
?^�n�b�ԫ^�"R��?��W(����y�����<���   �   f�z�io/�͖�qD����)�tӸ��yE����
����}��̽����Q��������������A־=7��D����<�׾�¾ϧ��މ�XjV�~���ԽTӆ���,����R������,�꼒�l
��#0�4{�[V����ܿ6�	��&�JD�\�`��7y�0���1��M���y�<Aa�H�D���&���	�4�ܿ����   �   �J��c�F��`�C���?�?��Ƚ2�1�`���(&�Hj��8�0�4��|���W���G�+�l��������D3���D���/��ʳo��EK�Fc"���̢���A� ^Ǽ�e��&��Z�@�tVϽ�C��~���c�0�G�Bߍ�₿�č�������;��4_�/��7������sݞ��8��	Ð��d���i_�<�;��X�?���뾿�   �   �˙�KY��$�H쵾�DR�Tֽ�)� ����<`K�;�⩻�Zؼ��X�劧�8�὚����`-� h2�j.���!����w��&%���i�0������j;���;�]��,9� o޽yV�].��f��Z������п�U��(��M��ov��ɏ�㫡��˭����V���ơ�~Џ�"Av�f<M�:�'�J��*&Ͽ�   �   #����e��[�!����X^�T�L�%� ��8�Z�<$��<�
�<@A�:(Ɩ�x*&�����M���]Ƚ�KݽZ,��<߽�̽����q����4�H����V%���K< Ϡ<p�~<0����6�d����b�kþl����f�Q�����ڿ#���0��Y�"�����m8��9��¾�E=���0������ނ��X�ZE0��u��yٿ�   �   �z���i��1�C1ľU�b���㽆B%����:06�<|��< 1�<�a.<p�߼��@�����H��<���0��Q綽2���;����M����Q5���;�<��<���<�^��o6���콐9g���ƾ]���j�*���"J޿2}�V4�l�]����D���E��b�����������/�����ӝ����\�J3����ݿ�   �   r����e�5[�$����W^�wR�6�%� p�8l\�<��<�<@D�:Ɩ�j*&����M���]Ƚ�Kݽd,��<߽�̽����q��x�4������R%�X�K<Р<��~<��^�6���轃�b�jþ�����f������ڿt"���0��Y�Z!��8���h7���7�� ���0<���/��<���)ނ� �X��D0�Vu��xٿ�   �   6ʙ�IY�n#�i굾�BR��Pֽ�)� ����<�R�;�ީ�Zؼj�X�늧�;�ὢ����`-�	h2�!j.���!����u��!%���i�h������k;��;hS��(9��k޽�vV�s,���d��Z�H����п�T�l(���M�pmv��Ǐ�����ɭ����O���ġ��Ώ��>v��:M�̚'�2��t$Ͽ�   �   �H����F��^�������?�7	Ƚ��1�L����&��g��|�0��3��f���W��G�8�l��������L3���D���/��ͳo��EK�<c"���_̢�¡A�[Ǽ؃e�@����@��QϽ��C��{���a�k�G�cݍ�s����������
�;��1_��,��ʁ��J���ڞ�"6�������b��nf_���;��V�9�� 龿�   �   ��z�%l/�:��^A���)�Eθ�,sE�f�����>�}�<̽����Q��������������A־I7�E����C�׾�¾ ϧ��މ�CjV��}�+�Խw҆���,�ƿ�@�R����~�,�ɹ���꾬 0�0{�oS����ܿ�	�4~&���C���`��2y�U���.��+J����y��<a���D���&���	���ܿ���   �   TV������ľ#�u�vW�5�����i�P=f�>���c��
6�.1��Rf��K�־>.�מ�R$��.���1��s.���$�����`��dپ�٬�J����Y:����q��,�r��t�^�����w�n�žKT��@V� .���c��O��`p��'�^N>��NQ��9^���b�n�^�4R��?��S(����t�����9���   �   �/�`Z�M��VI�����禽�x��T
���)�2�G�~ޏ�3žb� �����7>��:Y�:�n��N|�����s�|���o�B�Z���?�G!������Ǿ����-K�-=��<��jԖ�8��������aJ�cY���W��/�N�q��c���ƿ���t��v���g,�L6�J�9��{6��	-�H��N��g��ǿ�ݞ��r��   �   +�
�9����rz��% �e�Խ�����ʽ�|�PI�6���=�Ҿ��4�6��=a�|����햿���k!���_��o{��ɯ��A����ԅ���b��r8�,b���Ծ}_��ܦK��~�M���O���ֽ�D �Vz�����I
�x�?��m}�`%��,¿Y���g��,����?�������S ����U9ÿk���s�~��@��   �   �rѾ�掾�+<�iv���������h����:��퍾�оח��IB�^�w�:)��-H��UEȿ�WڿT�忩)��s�s*ۿ�Iɿ6T�����S?y�~�C�Z��*wѾ�鎾�/<��z��W�����������:�-덾�о2��`FB��w��&��?E��Bȿ&Tڿ����%�p��&ۿ{Fɿ!Q��>���:y�ȊC�u���   �   �[��ΡK��{�����T���ֽ
G �Cz��!��L
�c�?�uq}��'���.¿���Xk��(!����A������U �%��G<ÿ������~�K�@���
�����*wz�|( ���Խ�����ǽ�Hy��I�ﵔ���Ҿ����6�9a����ꖿ�	��"��:\��x������E���҅���b��n8� _�ӫԾ�   �   I'K�"9��7���і��������EdJ��[���Z�^�/�X�q��e��r�ƿ���"��h���i,��6�¨9�6~6��-�T����{񿦓ǿ�ߞ��!r���/�^����YI��	��K覽�v�����M&��G��ڏ�9.ž\� �,��3>�6Y���n�(I|�������|���o�G�Z�*�?�-C!������Ǿ�����   �   ��[k��d�r�^�t����������w���ž�U�CV��/���e������q���'�rP>�TQQ�T<^���b�&�^��R��?��U(����ew�4���~;���V����ľb�u�7Y�K���v�i��6f������Z��d6�v-���a����־�*���/$��.���1��o.���$����^]��^پլ�T|���S:��   �   �ˆ���,�
��؎R�	����,�������"0�2{��T����ܿ��	��&�jD��`�5y����g0���K����y� ?a���D�4�&���	���ܿ���d�z��m/�����B����)��ϸ�<rE����p���}��	̽
�
�Q�\�������4����;־�0�i>�]���׾4|¾ʧ��ډ��bV�x��Խ�   �   (HǼxie�@��"�@��RϽ��C��|��~b���G�3ލ�����������4�;�3_��-���������ܞ�z7�������c��&h_��;��W����w꾿�I��6�F��_������?��
Ƚ��1�̌����%��V���0�C,����4R�G�G���l�\��?����.��i@���+����o��>K�4]"���;Ģ��A��   �   `kk;�ŝ;�H��'9�l޽4wV�-��(e�ȷZ�Ҝ���пTU�(�؜M��nv��ȏ�窡��ʭ����Y���š��Ϗ��?v��;M���'����w%Ͽ˙�?JY�F$��뵾�CR�@RֽL)�@����<@|�;p���,Gؼ��X�ʃ������ �����Z-�~b2��d.�u�!����́轖��
i��������   �   h֠<H�~< ����6���轨�b��þ���ۻf�Խ��Y�ڿ�"�@�0�r�Y��!�������7��r8�������<��^0�������ނ���X�E0��u�9yٿ���e��[�߄��nX^�rS���%�  �8$_�<���<��<@��:�����#&�D��`I���XȽ�Fݽ('��7߽�̽z����m��:�4������%��
L<�   �   �=�<P��<@���d�6����)Ak���ʾ�� ���o�p�Y��\��4B8�ښc������f���1�������|������-��<\�����~nc��8��S�{z⿲���o�z5 �6ɾ�Eh�q��Ե)����:�J�<�!�<���<غ0<@�X��v�D���������:���I��1����˧���|�N�������+��^�;�ީ<�   �   ���<H��<��W�67�C�"�f���ƾ\��،k�c��i(߿ �$5�t?_��������h���l�����m��������[ ���_�:�4������޿�ǥ���j�I��lžp�c���`V*� 0T��ף<�7�<��<@|�:`�����)�/ɂ�,Ы�o^̽�~�J?����LϽ�������Q5��ó�@�� -]<�   �   ��;`�;0N�,�9��Z�p2Z��Ȼ��m��V_�uޝ��oԿ6	���+���R�ª}�k����l���b������b"���m����}�z�R���+�B	��)ԿS���R�^�F������o{W��۽�g-���Ļ�\<���;�ֱ�@4޼Z^�Y|�����!�I#���0�l�5��1�q�$������(��V�j��~������   �   ��ļ@+]������nA�Xҽw�F�Ǫ��-��>L�u퐿6�ÿ����z�|�@�΄e�k3��fD��w=�� $���F��R��@����e���@��
�+���9sÿ5���$�K�¬����j�D�h�̽�:6��'��X4+�����:5�?���P�t-"�eL��;r�8'���⑾�]���?���ڈ�I9t�C�N�%�(x��y���AB��   �   L����-������S����j�/����������3��a��j�����r���*�HI�$g��t���I���s���U��R����Lg��hI�8�*����ʵ��
���D��@�3��=����-������I������!�%�ѽ����W����'٩�fvžd۾%��`����.ܾF|ƾ����p���$Z�����M׽�   �   `����`���t�nw��г�f�
�|�J�ɾ ���%[�������¿{�0����+�&wC�Z8W�b�d��^i���d��bW�6�C�f$,������^�¿0���N[�����Tɾ��{����~7��<�n��Hk�>���=��:�:��e��鳮��Uܾ�n�&P��(��*2���5�V^2��m(�������ݾ�0��S䄾�=��   �   |�N��j
�ż������Ҭ�B ��YN��̣�������3��Qw�(����˿�����R���!�T�0���:�nS>�*�:�^1�� "�*��8����˿�W���w�^�3�x���F���v�M�a0��g9��8l����H8�BYL��m���,ʾ���f�#�1C��^��\t�J$��A���v@����t��2_�z�C��$�����˾ Ĕ��   �   �Y���qO���	��ý�����ٽCf#��i�Q}¾����\D�`Ё�G���ƿ�4远��"���>���&�R����迬Gǿ�_�����E�D������¾���[#��ؽ�$��E����Z���M��N��;�׾���ߛ;�a�f�K��줚�&���3���e���S���?���������g��P<�f_��پ�   �   y�վ~֑���?������5���׽�����!�>��0���վ7-�� G��}��ꚿӥ���"Ϳ��߿�T��n￱x뿎�߿xͿ]���G��H~�͸G�`���վ�ӑ�[�?������4��iٽ�T���D�>��3��Gվ20��$G���}��횿����N&Ϳc�߿vX��r￑|�:�߿p{Ϳd��jJ����~�R�G����   �   ��
�¾����]#���ؽp#��~���~W���M�K��/�׾f��ԗ;���f�BH��ޡ������0��Ub��!P��z<���k�����g��L<�_\�@پ-V��NmO���	�H�ý������ٽ"i#�In��¾}��
`D�zҁ�����ƿg8迊��>��H�|��)�`����1�迀Jǿ3b�����D�D��   �   ��3�����p�����M��2��9��li��!븽4�@SL��i���'ʾR��t�#��C�Ԝ^�RWt�l!��Z����=��o�t��-_��C��$�Ն�˒˾=����N�>g
���������0Ӭ�� ��\N��ϣ�����6�3�2Uw�A*��b�˿�����T���!���0��:� V>���:��1��"���'"����˿�Y��1�w��   �   �[�R��Wɾ�{�����7��`�n��@k��7���4����:�ra��Ю���Oܾk�#L�*(�B&2�$�5��Y2�xi(�������ݾ,��~����y=����9[��d�t�Bw�ҳ�=�t�|���ɾ��<([�n����¿�}������+�pyC��:W�>�d��ai���d�peW�b�C�0&,�l����I�¿�����   �   �E����3��?�뿔�$�-�\��b�I�����!�6聽ѽ���lW����ө�~pž�]۾l�龐��^���ܾ�vƾ����l���Z�
��NE׽󇽈-�����S�����N�/�e���3� 4�1c��	����ῴ����*�JI�~&g�Fv��gK��Su��jW������ Og�PjI���*����������   �   ���V�K����	���l�D���̽B96����+�8����-5�����F�>'"��]L�q3r��"��%ޑ�$Y��&;��nֈ�c1t�G�N�#�$�Hn��*q���5B���ļ�]��󠼲nA��ҽ6�F��Ȫ��.��@L����ÿ�������@���e��4���E���>���%��6H���S��A����e���@�������Ptÿ�   �   ߖ���^����]���|W�j�۽df-�PqĻ�n<��; ����޼:^��t�������C#���0���5�C�1�!�$�� �뽛 ��
�j�Dk�����F�;�;�G���9�Q\��3Z��ɻ��n��W_�Gߝ��pԿ�6	���+���R�6�}��k�� �����t������Q#��Nn��У}�^�R�:�+��	��*Կ�   �   �ǥ�;�j�BI��lž��c���tU*� �M��ܣ<�>�<|�<�&�:t�����)��Ă�X˫�=Y̽}y��9���BϽl�������J5�L���@]��:]<앪<��<��W��7�R��f���ƾ�����k����)߿z ��5� @_�X��>������/m�����Wn�����w���� ��@_���4���H�޿�   �   �����o�K5 ��5ɾ�Eh�����)����:�K�<|"�<t��<��0<@	���
�D�_���a���:���I��)����˧�#����N����@�+��\�;ީ<,=�<h��<@μ�2�6�E�ｐAk��ʾ� ���o��򨿃��v��PB8���c������f���1�������|������-��-\��|��^nc��8��S�Qz��   �   ǥ�-�j��H��kžD�c�R��PS*�  H�$ޣ<�?�<�<�,�:D�����)��Ă�]˫�CY̽�y��9齉��KϽn�������J5�����W�H<]<���<̍�< �W��7�����f���ƾ*����k�-��(߿���5�?_����S������l�����;m�������������*_���4�n��\�޿�   �   �����^�`��n���yW�)�۽Lb-�p\Ļ8u<@�;����X޼^��t�������C#���0���5�O�1�)�$��#�뽑 ��ހj�|j��`��0O�;�+�;x=���9�Y�Q1Z��ǻ�nm��U_��ݝ��nԿ�5	�X�+���R���}�Sj��-��e���P������_!���l��*�}�b�R���+��	��(Կ�   �   #�����K����]����D�p�̽�36�����+������,5����{F�:'"��]L�z3r��"��,ޑ�*Y��-;��tֈ�j1t�H�N��$�-n���p���4B���ļ�]�h젼�hA�cҽ��F��Ū��,��=L��쐿 �ÿ������H�@�4�e�f2��.C��<���"��oE��3Q���>��(�e� �@��	�s����qÿ�   �   �C��`�3��:�¼����-�����I�p��x�!�p災ѽ���`W����ө��pž�]۾x�龜��g���ܾ�vƾ����l���Z�����D׽;��-�ƚ���S�(~���/�5���y��J�3��`������\����*�RFI��!g��s��jH��;r��mT������jJg��fI���*�p��ȳ�(	���   �   �[����RɾH�{�z���1�� �n��;k�=6���3����:�ca��ɮ���Oܾk�'L�/(�H&2�*�5��Y2�|i(������ݻݾ,��m����y=�����Y����t���v�F̳�����|���ɾs��A#[�-�����¿�x����+� uC��5W���d�\i��d�P`W��C�|",�^���5�¿t����   �   ��3�z���`���'�M��)��43���e���踽d3��RL��i���'ʾP��s�#��C�ڜ^�XWt�p!��]����=��u�t��-_��C��$�҆���˾ �����N��f
�@�������Lͬ�\ �VN�zʣ�<���.�3��Nw�&��I�˿����BQ���!��0��:��P>���:�1���!�T������˿�U����w��   �   Q��.�¾^��\W#��ؽ����~��fV��M��J���׾`��ԗ;���f�DH��ᡚ�����0��Yb��'P��}<���l�����g��L<�Y\�&پ�U���lO���	���ý�����ٽ�b#��d� z¾����YD�s΁����3�ƿ�1�����������$�<���{�迭DǿE]������D��   �   ��վ\Б�L�?�	����-���ҽ�Z���-�>�h0���վ/-�� G��}��ꚿ֥���"Ϳ��߿�T��n￵x뿑�߿xͿ`���G��H~�ʸG�W��V�վuӑ�\�?������/���ѽ�������>��-���
վ{*�3G���}�`蚿֢��wͿ��߿�P��j��t���߿�tͿ= ��E���z~���G�a���   �   KR��vgO�D�	��ý������ٽ�d#��h�}¾���\D�^Ё�G���ƿ�4连��&���@���&�T����迭Gǿ�_�����?�D������¾��0Z#���ؽ���'|���S�F�M��G��{�׾[���;��f��E��잚�����'-���^���L��79���욿����.�g��H<�Y�"پ�   �   ��N�db
�����B���ͬ�t ��XN��̣�������3��Qw�(����˿�����R���!�V�0���:�pS>�.�:�`1�� "�*��9����˿�W���w�U�3�M���򨣾V�M��,���3���c��^丽�/�pML��e���"ʾ6����#�>�B��^��Qt����z����:����t��(_���C�(�$����|�˾����   �   ޲��[S����t��v�z̳���2�|��ɾ���%[�������¿{�0����+�(wC�Z8W�f�d��^i���d��bW�8�C�f$,������a�¿1���J[�����Tɾ��{�J���2��ʫn�V5k��0��q+���:��]�������Iܾ�g�EH��(��!2���5�VU2�+e(�������ݾ�&��`܄�Ps=��   �   b뇽L-���z�S��~��Y�/�l���v����3��a��k�����t���*�HI�$g��t���I���s���U��R����Lg��hI�8�*����͵��
���D��7�3�}=�e���ک-�x����I����.�!�:ၽѽ+��IW������Ω��jžaW۾��ׂ�龉ܾ�pƾ���&h��1Z�����;׽�   �   ��ļ��\�L䠼\gA��ҽ��F��ƪ�u-��>L�u퐿7�ÿ����z�|�@�̄e�l3��hD��w=�� $���F���R��@����e���@��
�-���;sÿ5���!�K����Ԭ����D���̽x36�L��H�*�H骼� 5������<�O!"��VL��+r�����ّ��T���6��҈�c)t�"�N���$��c���h���'B��   �    ��;@O�;�2�b�9�_Y��1Z��Ȼ��m��V_�vޝ��oԿ6	���+���R�ª}�k����k���a������c"���m����}�z�R���+�D	��)ԿS���Q�^�@�������zW���۽�b-��PĻ��<�F�;`S���
޼ ^�=m��6��I�v>#�Z�0�
�5���1�˝$�&�K�����tj��U��@���   �   H��<���< �W��7�����f���ƾ\��׌k�d��l(߿ �$5�t?_��������h���l�����m��������\ ���_�<�4������޿�ǥ���j�I��lž7�c�W���S*� �F���<@D�<��< ��:����)������ƫ�^T̽Ttὁ4�>��2Ͻ����ã��&C5���������L]<�   �   ̡�<L��<�G8;[#�����:d�ƾT��P�k�Dt����߿p���5��Y`�������w��G���$���p������Z�� ����`�,:6����fL࿻֦�El�D���ž�c�P�ʻ��ة;�`�<,�=|��<��f<pف��%Ƽ�*5�Θ~��X����2Ե������'݁���;�(Pּ@�˻��><��<�   �   �c�<ļ�< [~:��#����_�EY¾�D�g�˫���ܿ"6���2��\����&_��b��ݤ��n9��â��Th��x��"?��\�
3������ܿA���h��!�f¾B�^��OݽS�@�X;x+�< S�<H��<���;p]{���DKu�q1��oGý��׽�_߽��ؽ��Ľ������{���"�丏��r ;d��<�   �   �T<Ȅ!<𡝻�`&��Iֽ�sS��|��r��Y�[�F�����ѿr���)�T(P�l,z��M��C�������`����>����J���Mz��fP��*������ѿAٛ�[\�Ƴ��9��pJR�g�ҽF�`)�x�H<@95<�������N�*#���޽W	�21� �+��`0� �+�<���t
��ཇɦ�D�V��qӼ����   �   Da���J�p4z��T.�Aǽ��@����W��m�H��ӎ��
�������0��H>���b�u���:������6����ݝ� ��GU����b�DP>�.N�����M�����sI�ϝ�;{��dt?��5Ľ��&���X���仌���&�k땽���c��,G�t�l���V���*���ǎ��b��@tm�gH�x��@:�����.��   �   ��{�bC��,�l�@�\��D�)��瑾�L꾭1�C}�٫�6߿�N�,�(�^	G�6pd���}��w���{���V��hP}�Nd��F�:�(�hH��߿x����A}��#1��L�+���4�(��i��$3:����V�0�s���Ƚ|$���Q��%����������+�׾�u�	C�ƃ�f�׾�6¾_��ݹ���gS�'���`̽�   �   $���>-��N\a���c����o��v��ž��O�W�����6���m��l��;*�VlA�8�T���a��Zf�$�a��iT�t�@�<�)�F3����!q��`���eX�%$���ž۫u�d������y^�:+[�ߚ��9���5����܋����ؾvo�j�˜%���/�B�2�Ă/�P�%����~�پ(��l>��!7��   �   �WH���%����P���I����HH��,��'q���$1��t��?��
dɿ�Y�"��= ��
/��8��<���8�D�.�������%���ɿ� ��� t��,1������1��|H�����n��6䌽[.����� G��r����ƾv����!���@���[�Iq���~��ˁ���~�Sq��[�S`@�%�!�����Ǿ����   �   ���`&I�NT�@ù����}�Ͻi���y�����R�>�A�H;���B��z�Ŀ�������y�&���R�����F�n忹�Ŀ&�����r�A�o]�[྾�Ty�J���IϽa���i���~��AH�S1���;Ծ���.9�/d�����w똿O������*��� ���馿䰘�%�����c��9�v����Ծ�   �   ��Ѿ�K���9��󽼩��~k��t��h9�����NѾ�����D���z�{<��Zų�3˿Y9ݿ���f��k����ܿƧʿGj������r�z�ljD����ąѾI����9�Z��ڨ��Rm��2��4l9����<SѾ�����D���z�9?��{ȳ��˿=ݿ���T��@��d�ܿ�ʿBm��w���Ōz��mD�X���   �   �_�m㾾�Xy����)KϽP��f��_{��<H��-���6ԾT��*9�U*d�ɻ��o蘿�����>'��E���x榿��������!�c�$9�w��I~Ծĕ���!I�tQ�z�������Ͻ<���!y�����U���A�^=��ME��w�Ŀ�������{�^��U�����H�Rq忇�Ŀ��� ��k�A��   �   �.1�ي���3���H�4���#n��uጽ)��{~�.G��n����ƾ2����!��@���[��Cq���~��ȁ�/�~��q�)�[��[@�f�!�����ǾW����RH�^�������펽���������KH�R/���t��'1�ct�B���fɿ�\���� ? �/�f�8�<��8���.����<����K!ɿ�"���t��   �   �X��%��žm�u��������8u^�#[��ؚ�i0���5����Ά��տؾ�k�n�}�%�9�/���2�N~/��%���@{�@پ_���:��S7��|���'���Ua���c�/����p�=v���ž����W�a���^�����m��=*��nA���T�|�a��]f��a�0lT�� A� �)��4���s��៓��   �   �C}�x%1��N�`���h�(�j���0:�$v�M�^�s��Ƚ����Q�|!��ȣ������Ќ׾6o�L<�,}�*�׾G1¾W�������`S����X̽��{�(;�(�z�@����$�)��鑾:O꾂1��}��ګ�5
߿�O���(�FG��rd�b�}�cy��}��.X��S}�~d���F���(�~I�}߿�����   �   ���� I����7|��fu?�6Ľ�&� zX���������%�㕽:{��\�c%G�m�l����Š��������B^��olm� `H����0�?����.� P��P4�)z�|T.��Bǽf�@�����t���H��Ԏ���������1�J>�b�b�+v��"<���������'ߝ�V��IV��V�b�vQ>�O����N���   �   �ٛ�#\�M���:��KR���ҽ�D���(�`�H<�R5<��������tN�u����ݽR	��+�~�+��Z0���+����p
����6¦��V��^Ӽ�R��(j<X�!<p���\a&�0Kֽ&uS�~��R����[������ѿ�r���)�j)P��-z�fN��C�������a��!��)����K���Nz�lgP�`*�0����ѿ�   �   w��h��!��¾k�^��Oݽ$R� �X;P0�<�Y�<���<0"�;�C{�����Bu��,��EBý{�׽kZ߽��ؽ��Ľ0�����{��z"�`���@� ;D �<th�<���<�w~:\�#���p�_�Z¾���g�J���~ܿ�6�~�2�� \�U���_���b��q����9��J����h��ux��n?��.�\�V3����ܿ�   �   �֦��Dl��v�ž}c������ ީ;�a�<��=L��<�f<�ց��$Ƽ�*5�z�~��X���� Ե������4݁���;��PּЁ˻�><\��<��<\��<@>8;�[#���%;d�Mƾ�����k�it����߿����5��Y`����)���w��O���%���i������J�� ����`�:6�|��<L��   �   ����h�*!��¾�^��MݽP�`�X;2�<�Z�<P��<�#�;�C{�����Bu��,��KBý��׽uZ߽��ؽ��Ľ2�����{��z"�0����� ;� �<ti�<L��< �~:2�#�d���_�Y¾����g������ܿ�5���2��\�����^���a��W����8��0����g���w���>���\��3�J���ܿ�   �   s؛� \����8���HR�z�ҽ�@���(���H<xV5<`��4����tN�r����ݽ"R	��+���+��Z0���+� ��p
����2¦���V��]Ӽ�M��@n<ؘ!<����@]&��Gֽ�rS�)|������[�����Ґѿ�q�D�)�x'P�@+z��L��Z�������_����=���	J��0Lz�teP��
*�����ѿ�   �   ����I�����y���q?��1Ľd�&��kX��p�X����%��╽{��\�c%G�r�l����ˠ��������J^��wlm�#`H����h0�
����.�`M��p+��z��N.�#>ǽ�@�۽��~��=�H��Ҏ�u	�������/��G>��b�t���9��S���к��mܝ����.T����b��N>�M����WL���   �   s?}�#"1�J�9���H�(��d���):��m�nJ���s�8Ƚb�t�Q�x!��ˣ������،׾?o�U<�6}�3�׾O1¾Y�������`S�r���W̽��{�~8��#���@�����)�\摾�J�01�=
}��׫��߿�M�κ(��G�nd��}�uv��z��?U���M}��d�$�F���(�,G��߿�����   �   �X�)"��ž��u�+�������m^�t[�@ך��/񽀔5�����Ɔ��ѿؾ�k�q���%�>�/���2�S~/��%���B{�>پY���:��7��{��2&��Qa�@�c�o���^l�t
v���ž���W�+���R����j��9*�6jA���T���a��Wf�\�a�$gT�8�@�X�)��1����n�������   �   �)1������.��8H�D���[h���݌��&���}��G��n����ƾ-����!��@���[��Cq���~��ȁ�5�~��q�.�[��[@�f�!�����Ǿ:���#RH����\����鎽�������EH�K*���m���"1��t��=���aɿ�V�l��; ��/�|�8�
<�2�8���.�������
��>ɿ���'�s��   �   �Z��ܾ�Oy� ���BϽ����b��Dz�<H�t-���6ԾM��*9�S*d�ɻ��p蘿�����A'��H���|榿��������"�c�#9�s��3~Ծ����&!I�\P�Ｙ�-�����Ͻ���
y�����ZP�C�A�`9��k@����Ŀ���2�����w�����P�����D��j�ĀĿ������&�A��   �   E�Ѿ�E����9�������f��M��)g9�Z���NѾ����D���z�{<��Zų�3˿[9ݿ���l��n����ܿ˧ʿIj������r�z�ijD������Ѿ�H����9�0��٣���e�����c9�� ���JѾE��x�D���z��9��`³��˿�5ݿ��迄�쿒���ܿ[�ʿ.g��+���փz��fD�����   �   푕�I�M�M���,���.�Ͻ���y�̻���R�7�A�F;���B��y�Ŀ�������y�*���R�����F�n忻�Ŀ&�����n�A�`]�"྾�Sy����@EϽ����_��nw�q7H� *���1ԾO��P&9��%d�*����嘿���>���#������?㦿򪘿Ѕ��f�c�)	9�<��=yԾ�   �   ELH����!���?玽���������GH�k,���p���$1��t��?��	dɿ�Y�"��
= ��
/��8��<���8�F�.�������'���ɿ� ��� t��,1�l����1��`H�w����h���ی�J"�� z�fG�k����ƾ���!��{@���[�R>q�V�~��Ł���~��q�'�[�wW@���!�����Ǿ=��   �   �r�����0Ia���c������m�v�Рž��K�W�����6���m��l��;*�VlA�8�T���a��Zf�$�a��iT�x�@�<�)�F3����#q��a���bX�$���ž��u��������k^��[��њ�;'�Î5�6��������ؾ�h���M�%�΁/�1�2��y/�؊%���w�3پV����6���7��   �   \�{�/��N�@���:�)��瑾�L꾥1�A}�٫�7߿�N�,�(�^	G�8pd���}��w���{���V��jP}�Pd��F�>�(�jH��߿{����A}��#1��L�ܨ��!�(�7f���(:��d�:B�t�s��vȽ��j�Q�2��Ȟ�� �����׾�h徢5꾚v��׾�+¾0��$���TYS����zN̽�   �   <:�����
z�8M.��>ǽ�@�־��I��i�H��ӎ��
�������0��H>���b�u���:������7����ݝ�"��GU��b�DP>�2N�����M�����nI�Ý�{���s?�3Ľ^�&�h`X�PD�0ꍼX�%�!ە�eq�W��G���l�|��O���������Y���dm�YH�w��;&����"�.��   �   ؆<@�!<�k��0\&�FHֽKsS��|��l��X�[�F�����ѿr���)�T(P�l,z��M��D�������`����>����J���Mz��fP��*������ѿBٛ�Z\�����9���IR���ҽLA� �(�8�H<�k5<������hN�-��x�ݽ_M	��&��+�^U0��+���� k
���བ���<�V�,IӼ`���   �   �o�<�ũ<�0:T�#�P��G�_�7Y¾�E�g�˫���ܿ"6���2��\����&_��b��ܤ��l9��â��Uh��x��"?��\�3������ܿ@���h��!�X¾�^��Nݽ�P���X;�4�<,_�<��<�F�;(-{�����:u�6(��o=ýZ�׽-U߽V�ؽ��Ľ����t�{�Rs"�ܠ��`!;	�<�   �   �>=�^�<;+<���3:˽ϙR�φ��X�ϒ_�,P��|;տp�	�:�,���T�)���M��@y���Q���˺�W������+������|�U�x�-�޲
���ֿtM��{�`����`���S���ʽ����@<�`=��=�t=��< 7A;0@������X�q@��[��EF���V���㈽[���LǏ��n�:@��<�=�   �   �l=P��<P<����ǽzN����>�2�[�h�����ѿ8���*�n�P��){��
�������/��荶�7+������:����{�:�Q�f�*��j�
ӿI���z�\�"�ڿ��m�N��ƽL����"< ��<x�=�<�`;<�(����P�W���|B���ȽYy��� ���ߏ��S�����h��0�$<Ԝ�<�   �   @"�<ˌ< >J;H* �,����B������@
��-P��듿�ǿ >���!�0�E���l��ԉ�~Ӛ��Y���]���<��%���Ή���l��>F��f"������ȿW���=Q���
�L��bC����(4��pF�;|�<з�< "�;,>���*����|ǽ
���:����
�!�+��L���]��ChȽ9w��~�.������c;�   �   ��5� ��� ��Z��v���0�n������`A>�
������}�\�J<5�VW�p�x�������P���l���u���x�"�V��H5�jQ���֜��oG���?������4����0���������» �h8��"����Z��n�νG�ZK8��
\��Lx��1���F��Y��<x�f�[��H8�����ϽI��h��   �   �gR����(̹�X ��(�����ۇ��Zܾ�w'��\p�㻣���Կ���!� �=���X��+p��������pc�r\o��X���<��� � ��տ���|�p�2�'��ݾ�4������w���?�������ἤ�N���LQ
�V�B�"n~�Zh��|���˾XAؾ��ܾ�ؾ1�ʾ5
��\����}���B�8�
��H���   �   �ڽ�@���}9�H<� ���Z��=(d��l�������L�n���[����@�D�D�"��p8�<xJ�<mV��tZ��U�4�I���7���!���
����Ҋ��;����M�� �r͹� �d����w��<�9���6�� �ٽ�}'�2�o�j$��t̾w���A ����Z\&���)�6!&����d��������˾@���*�o���'��   �   R18�CHｸ���/t�Io��P�ܽj�8�+���la�b�'�Lh��̘�n��`�迚��":�n,'�*30�03���/�6q&��h�"�������em���g���'�����敾��8�U�ܽ��޷r��G��1��0,8�!���-������TO���6�v
Q�.�e��r���v�~%r�u�d��1P�-6�ݛ�8���y���K↾�   �   �c��((9�E��wf������17�4�g�!!����#�7��%t��՚�>5��?ܿg������J���7����d�����U�ڿ�9��'���Qs�;\7��������g��T�޴���^��t���e#9�V���? Ⱦ�����/��"Y��h���ܑ�
v��3
���ݪ�s���;螿�1��|��/X��/�Tj��qǾ�   �   ѽľJ����*��۽~7Ӟ�n�ڽ��*�����4ž���:���n��3������;¿�ӿ~޿��޿��ҿS#��ͪ��k��y�m���9���
��ľ������*�`۽�ힽ�Ԟ���ڽ��*�����fž����:�A�n�-6�� ���� ¿��ӿ��޿�⿨޿�ҿ�&���Ϫ�wn����m��9�!�
��   �   �����~�g��V�e����]�������^9�ϓ��y�Ǿ�����/��Y�Xf���ّ��r������ڪ�;���,垿�.��v|��X���.�vg��mǾn`���#9�����c��ϛ��{����9���g�$��>��I�7��)t�Gؚ�8���ܿ �����`�� :�����f�B���q�ڿo<��S)��CUs�_7��   �   �'����镾.�8�b�ܽ�����r��B��9��~&8�5���(��^����K�R�6��Q���e���r�E�v� r�V�d�@-P�6�K��S���Ώ���ކ�*,8�2A�q��(,t��o��`�ܽr�8�����e���'��h��Θ��p��_��X��<��.'�|50�t23���/�Vs&�jj���O��f���Io����g��   �   �M�V��Ϲ�x�d� �������9���6��톽I�ٽ�w'�s�o����.n̾����p�c��	X&�/�)��&������������˾�����o�.�'��ڽQ;��4w9�.<������p+d��o������L����k���&C����"��r8��zJ��oV�fwZ���U���I���7�`�!�Z�
�ʺ忨��������   �   u�p���'��ݾ�5����bx���=����D��\�N��貽�K
�2�B��e~�\c��hv���˾�:ؾ<�ܾ��׾:�ʾ������o�}��B�ܢ
��@���[R�Ƞ�pù�r��"*������܇�G]ܾSy'�;_p�k�����Կ�l!��=���X�&.p�^������f��^o� X�x=�&� �*�1տ����   �   :H��	?�H����5����0���������» `�88h"�0 ��R����νA��D8��\�NDx�K-���B����x���[��A8�@����Ͻ����\�x�5� 퓺p��H�Vx����0�Ұ������B>�Ç�����W�`��=5��W�t�x�Ċ���������m���v���x���V��I5�HR���㝸��   �   ެ���=Q�X�
��L�� C�Y���2���[�;0
�<�Î<@b�;�)����*�!���xsǽ�����������!�֖�A���T��`Ƚ2p����.�� Nd;�,�<�ь<�VJ;�* �w���s�B�ɝ��aA
��.P�c쓿�ǿ�>�l�!�2�E�֝l�^Չ�jԚ��Z���^���=�� ����Ή���l��?F��g"�����ȿ�   �   �����\�S������N��ƽ���H�"<���<��=,�< u;< �L�P�d鎽h���S=���ȽIt��-��cۏ��R�`���(����$<���<Fo=��< <`��{�ǽ�zN���Y?��[�ߨ��6�ѿ���r*��P��*{�%�����w0��q����+�� ���e:����{���Q���*��j��
ӿ�   �   RM��C�`�n���_��JS��ʽ��򼀄@<Pa=8�=:u=���<@=A;x?��~���X�S@��>��6F���V���㈽*[�,���Ǐ� i�:Ȟ�<J=`>=^�<9+<`���:˽.�R������
�_�PP���;տ��	�V�,��T�)���M��My���Q���˺�W�������������`�U�b�-�Ȳ
���ֿ�   �   Д����\������N�N�d�ƽp���"<`��<,�=��<�u;<��,�|P�j鎽l���^=���ȽNt��5��kۏ�
�R�P���о���$<��<�o=���<`<H��ݫǽ�yN��񵾤>��[�3���W�ѿ���*��P�f){�S
�� ���m/��`����*��'����9��*�{���Q���*�.j��	ӿ�   �   �����;Q���
��J����B�<���*��Pp�;D�<�Ŏ<Pg�;�(��P�*����vsǽ�����������!�ޖ�I���T��`Ƚ2p����.�<����Vd;�.�<�Ԍ< ~J;�& �f����B�����@
�-P�듿c�ǿ�=��!�f�E�x�l��Ӊ��Қ��X���\���;��6���=͉�L�l��=F�"f"�����ȿ�   �   iF��f?�����33����0�Ҵ��
��p�» ؅8�b"�`��fR��b�νA�{D8��\�TDx�P-���B����x���[��A8�<����Ͻ����[�(�5� ����j���t��=�0�K���W���>@>�E�������i|�2;5��W���x�����v�����Rk���t���x�~�V�PG5�dP��ￅ����   �   �p�i�'�cݾ�2����Fs���6�����,����N�9貽kK
��B��e~�\c��jv���˾ ;ؾE�ܾ��׾B�ʾ������l�}��B�¢
�/@��(ZR����,������
%������ه��Xܾ(v'��Zp�����V�Կ���!���=���X�H)p����,����`��Yo��X��<�f� ��
��տ ���   �   �M�����ʹ���d���� ��x�9�n�6�n솽p�ٽ�w'�J�o����&n̾����r�f��X&�3�)��&������� ����˾����ҙo���'�3�ڽ�9���r9�<���������$d��j������L� �������f>�����"��n8��uJ��jV�$rZ���U�؟I���7���!�x�
����������   �   ?�'��|�:䕾��8�˛ܽ$���X�r�:@��ԝ�&8����(��S����K�P�6��Q��e���r�K�v� r�\�d�D-P�6�J��N���Ï���ކ��+8��?�3��%t�?j��Ǚܽ�8�й��)^�%�'�Uh��ʘ��k��������B8�R*'��00��-3�P�/�o&��f�h���翋���Nk����g��   �   �}�6��l�g��P�6���MX��x񢽄\��9�����\�Ǿ�����/��Y�Xf���ّ��r������ڪ�=���/垿�.��x|��X���.�sg�|mǾ?`��'#9����d`��}���Q����3���g�������G�7��!t��Ӛ��2��$�ۿ������@���5����b�#����ڿ�6���$���Ms�Y7��   �   ��ľz�����*��۽瞽[Ξ�Z�ڽ��*�D���ž���:���n��3������;¿�ӿ~޿�޿��ҿW#��ͪ��k��z�m���9���
��ľj�����*�V۽�螽�͞���ڽh�*�����Jž1���:���n�1�����¿��ӿ[z޿T�L޿�ҿ ��ʪ�ai���m�+�9���
��   �   �\��@9�S���\��}���ԩ���5�j�g�� ��Ҫ��7��%t��՚�=5��?ܿg������L���7�����d�ĩ��X�ڿ�9��'���Qs�7\7�������g��S�����0X���W9�p�����Ǿ��� �/��Y��c��ב��o�����oת�����➿,��Cw�R�W�,�.�ad��hǾ�   �   &&8�8�-���t��i��כܽW�8�ڻ��Ba�W�'�Gh��̘�n��_�迚��":�n,'�,30�03���/�8q&��h�"�������fm���g���'�a�澭敾��8�ܞܽ������r��;��ϖ�� 8�����#��m����G�"�6�� Q�ҁe�>�r���v��r�)�d�u(P���5�������͊���چ��   �   ��ڽ�3��k9��<��������g'd��l�������L�n���Z����@�D�D�"��p8�<xJ�>mV��tZ� �U�8�I���7���!���
����ӊ��=����M�� �9͹�,�d����%��`�9�$�6�熽q�ٽr'��o�����h̾"�����\���S&��|)��&�w���K���>�˾ݤ��*�o��'��   �   >MR�����������%������ڇ��Zܾ�w'��\p�代���Կ���!� �=���X��+p��������rc�v\o��X���<��� � ��տ���~�p�-�'��ݾw4������t��6����T����N�ಽF
�^�B�T]~��^���p���
˾�4ؾܧܾb�׾>�ʾ@���������}�ڕB��
�h7���   �   ��5� ܒ��K�^ ��t��6�0�9���ڨ��\A>�������}�\�J<5�VW�r�x�������P���l���u���x�"�V��H5�jQ���؜��pG���?������4��:�0�F�������» ��8�A"����J���νn;��=8�l�[�4<x�)��%>�������w�`�[�8;8�l���Ͻ����O��   �   T:�<݌<��J;�% �������B������@
��-P��듿�ǿ>���!�2�E���l��ԉ�Ӛ��Y���]���<��&���Ή���l��>F��f"������ȿX���=Q���
��K��� C������*��P{�;��<Ў<�;t����*�!�`kǽe�����`��B�!����6��dK���WȽ�h��|�.�p܋�@�d;�   �   �r=0��<<���ʫǽ�yN����>�0�[�f�����ѿ8���*�l�P��){��
�������/��鍶�8+������	:����{�:�Q�f�*��j��
ӿK���{�\�"�̿��2�N�f�ƽĜ���"<��<r�=H�<Ȇ;<��4���P�!厽����m8���ȽKo��c���֏���R�D���0�� �$<��<�   �   ��:=�%=재<�P���ԥ��7�&��&��jL��@��ddĿ�@��>&��`B��[h��E�����DT���Y��5Z����������Yi���C��_ �R8 ��-ƿc���r�M��P��ɧ���9�g)��@y��ث�<�%=Jj;=�s'=�L�<�xP<�뱻Hh��b-!�J�T�vcu�1��\�t�v�S� ���O��0��`�P<4z�<¸&=�   �   �('==P�<p\��Z���.4������j��^H��ʎ�5��U7��"��P?���c�Jy��㠔����a���N������ʯ�� �d�D
@�X��5����¿����=J����k���6�_Ԥ��w��lޝ<�^=.�'=��=<8�<��#;�����~Ea�\�����="��Ѧ��%Q���_�������*;�<�V=�   �   ���<���<�g<Ș��	o���&)�:��2����=�N����뷿:y��a5��mW��)y��>���A�������������y���W���5���f��t8������_?�{Z��V���h�*�Ӂ������2e<��<d�<�cm<04��(*�z�a�A���ӽB���#�<�����E���I�ҽL�js_��F�P�����m<�   �   �sk:��&<@&�;xߡ��b�����|���?�1>-�r�x��J��$
ܿ2�	�<�&�4�D���a�@�z�����ֈ�s����'z��Da��zD�x�&�j�	��ܿ#���+z��j.�1�侺ȋ��%��/������`�;�$<��@:����rJ�#��|����!��B�$$\��l�;r�>)l�)[�l�@�:��w����y����G������   �   B
�ؓ|�x*$�|>ļf�|����߳p� nƾy5�Y�[��z���aĿ�������P.�
uF�εZ�6Ah�l�l�d�g�<�Y�>|E�l�-�ZB�	�����Ŀ�ؖ�5�\���u�Ǿqtr���������Ǽ��(�L���p���4�����*��b�D��������#þ-!Ǿ]�¾t=��*����#`�(8)����򼐽�   �   ����FP�xb��rj��7f���޽��H��F��� ��;�A뀿|;���Կ6� ��� �)���9�BD�6�G�F�C���8���(��1�����Y�ӿD���t뀿�H;�4� �&�����I���ཬ�h���<�"OR��J����O�T��q��􀸾��߾� ����:t�hM�����K �O�ݾsE*���R��9��   �   ����ǽhv��/7��q[�wX��� �`i��b�Ͼy��&_T�:r���r��K׿�'��.��>=�$U"�J�$���!�$S���WG��ˬտǀ���ꋿ��S���6!о˳��<!�)`���]�
�8�V�w��dɽ.� ���p������޾p��{�&��/?��,R��*^�xb�ԕ]�n#Q��=�}�%��Y
�*�ܾ�����n��   �   �>w�0� ��ȽjG��lb�bY��ի��X:L�����-��o�'���_��j��w����?˿�@�̄���#��-�l��&��C�㿏�ɿt>��u��Ʌ^�9�&�n�����;L��
��Ж�~�b��؂��Ƚ��!�D�x�LH��p���5h ���F�A�k����鴒�ݥ���6��{6��|w����i��E��������
���   �   �����j�P��EE��b:}�P}�rz������k�}s������@e*�"�Z�h��];������EÿkͿ|�п��̿M-¿5ű�H�L���?Y��>)����������j�8���A���8}�@S}��~��s �#�k�]w������h*�G�Z��j��.>�����HIÿ�nͿ��пZ�̿�0¿0ȱ���O��wCY��A)�� ���   �   U�>����>L����~і���b��Ղ�"�Ƚ��!���x��C�������d �t�F�Y�k��������Ӣ���3��{3���쑿���7�i��E�?���������8w�� �� Ƚ�D��b��[��Ͱ��}>L�ļ�����Y�'�f�_�Dm��'����B˿D�y���x%��/�N��������u�ɿ�@��8w��2�^���&��   �   ���$о����x!!�b���]�(�8���w��]ɽ�� �p�p�3{���޾��p�&�:+?��'R�n%^�Ub�ΐ]��Q���=���%�XV
���ܾD���n�Ū���ǽh�u�B,7��r[�G[��� ��k����Ͼй�=bT�-t��u��׿�*�����8?�>W"�j�$���!�U����ZJ��c�տ񂰿r싿��S��   �   �J;��� ����9�I�����h�"��4��CR��B��Vz� �T�Xm���{��H߾0����;p�\I�����G �D�ݾP鶾	&��R�R��4������<P��V��lh��9f��޽��H�:I���� ��;��쀿h=��d�Կ�� �Z!���)���9�`DD���G�~�C���8�n�(�3�c���w�ӿ�����쀿�   �   �\�b��7�Ǿ�vr�������l�Ǽp�(������U,��u��q�*��	b�� �����'��þ7Ǿ��¾�7��"
���h`��1)����W���4��v|�0$��<ļ��|�]����p�[pƾ7���[�|��pcĿ����d��&R.��vF���Z��Ch���l���g�N�Y�~E��-��C�����+�Ŀ�ٖ��   �   H-z��k.���侚ɋ��&�r0������@&�;��$<�'C:<n���J��������	!��B�m\�ԯl��2r�B!l��![���@������*q����G��硼�^m:��&<�:�;Dߡ�6d����Ŗ��A㾙?-�V�x��K���ܿ �	�`�&���D�~�a�D�z����	؈������)z��Fa��{D�|�&�6�	�b�ܿ ���   �   5����_?�m[��귚���*��������<e<(��<�*�<��m<�瞻���a�&9��2�ӽ����"�.��̵������ҽ�壽\f_��0꼀Q����m<x��<,��<��g<����6p���')�;������=�����췿]z�l ��b5��nW��*y��?���B����� ��s��:y��W���5����D��9���   �   ���>J�G���k���6�LԤ�Xv��\�<a=*�'=`�=�A�<@S$;���
��<a�������m������L����_����p����*;D��<�Y=�*'=P=0�<�]��=��� 4�7���Pk��_H�$ˎ��5��8������?�0�c��y��X�������ۋ������u��������d��
@����t5���¿�   �   C���=�M��P�xɧ���9��(���w�����<x�%=�j;=Lt'=LM�<�zP<0鱻�g��-!��T�>cu�1��J�t�z�S�2���O��p	����P<�y�<��&=n�:=�%=��< R��ե�p�7�d��O���L��@���dĿ�@��V&��`B��[h��E�����JT���Y��0Z����������Yi�~�C�p_ �>8 ��-ƿ�   �   �� =J�����j��t6��Ҥ�hr����<�a=��'=��=(B�<`U$;� ���
��<a�������v������L����_����`�� �*;���<
Z=F+'==��<�Y�������
4�T����j��^H��ʎ��4���6�����?��c��x����������犣�ѡ������a���t�d��	@���d4��1�¿�   �   �����]?��X��4�����*�/������8Fe<`��<�,�<P�m<`䞻P�z�a�9��1�ӽ����'�6��е������ҽ�壽Zf_��0�PO���n<D��<��< �g<0���_m���%)�g9��;��?�=�՞���귿jx�2�>a5��lW�b(y�>���@������������y�ҶW���5�d��>�ￆ7���   �   �)z�*i.���<ǋ��#�j,��4��� A�;0�$<�C:xl���J����c���z	!��B�o\�دl��2r�G!l��![���@� ������q��t�G�,桼 �m:�&<�T�;ա�:`�����p����=�%=-��x��I���ܿp�	�B�&���D�2�a�\�z�|���Ո�Y����%z�$Ca�0yD�N�&�x�	���ܿ����   �   ��\�h���Ǿ�pr�>�����Ǽ��(��������+��$��V�*��	b�� �����*��"þ<Ǿ��¾�7��(
���i`��1)�y���������pl|��
$��0ļv�|����/�p�=lƾ(4���[�jy��)`Ŀ������$O.�LsF���Z��>h��l��g��Y�`zE�ؖ-�
A�۱��ӏĿ+ז��   �   fF;�q� �����.�I��ང|h�b�t0��@R��A��z���T�Hm���{��D߾0����=p�_I�����G �H�ݾO鶾&��6�R�q4�צ��B:P�XN���a�`/f��޽��H��D���~ �� ;��逿�9����Կ� �8�<�)���9��?D��G��C���8�ȭ(��/�����ӿX����逿�   �   ����о<���j!�
Z��b]�B�8�t�w�9\ɽ{� �,�p�{��Ջ޾��l�&�9+?��'R�q%^�Xb�А]��Q���=���%�YV
���ܾ:����n�h��;�ǽ0�u��%7�8h[�HS��߀ �0g��[�Ͼf��d\T�yp���p���׿�$��t��T;�S"�.�$�|�!�.Q�*��*D���տk~���苿��S��   �   ���5~��56L�Y���ɖ���b�c҂��ȽR�!�Z�x��C�������d �p�F�W�k��������Ԣ���3��|3���쑿���;�i��E�>��������f8w��� ���ǽ�A��,�a�T��Y���6L�����/��ş'�B�_��h�������<˿h=�>����!��+��������㿊�ɿ�;���r���^�K�&��   �   ������j�����:��~,}��F}��w����$�k�Ts������8e*��Z�h��\;������Eÿ
kͿ�п��̿Q-¿7ű�I�L���?Y��>)����f���Y�j�V��?���/}�\E}�>t����V�k��o��ރ�� b*�A�Z��e���8������Bÿ�gͿ�п��̿*¿%±��윿_J���;Y�6;)�����   �   �1w��� ���ǽt>��J�a�lU��J����9L�o�����e�'���_��j��u����?˿�@�̈́���#��-�n��+��G�㿒�ɿw>��u��ʅ^�4�&�T��O���X:L�\��!̖�d�b��ς��ȽH�!�{�x��?��U���Ha �g�F���k�\��#���ӟ���0��x0���鑿*��d�i��E�������o���   �   4����ǽ��u�� 7��g[�%U��� �i��8�Ͼn��_T�8r���r��J׿�'��,��>=�&U"�J�$���!�&S����ZG��άտǀ���ꋿ��S���!о����<!��\��n]���8���w��Uɽ�� ���p��v��^�޾�����&��&?�#R�m ^�=	b�Ƌ]��Q�=�=���%��R
���ܾ�����n��   �   Ǟ���.P� @��v^��/f�A�޽�H��F��� ��;�@뀿|;���Կ6� ����)���9�BD�8�G�F�C���8���(��1�����[�ӿG���t뀿�H;�(� �����$�I��཈~h�j
��*��6R�L:���t�@�T�i��Zv��7y߾�� ��Kl�ZE���H�0D ��ݾ�㶾�!��&�R��.��   �   ����J|��#�@,ļH�|�Đ�G�p��mƾp5�T�[��z���aĿ�������P.�uF�εZ�8Ah�n�l�f�g�>�Y�@|E�n�-�\B������Ŀ�ؖ�5�\�
��O�Ǿ�sr������D�Ǽh�(�P���p��=$��6���*�.b�/���������TþOǾ��¾j2��	��늾�`�\+)���Ԭ���   �   ��o:��&<�q�;Lҡ��`��ڛ�J����>�,>-�p�x��J��%
ܿ4�	�<�&�4�D���a�B�z�����ֈ�s����'z��Da��zD�x�&�j�	�"�ܿ%���+z��j.��侈ȋ�8%��-�����0U�;P�$<�mE:TW��2 J�������b!��B��\��l��*r�Ol��[���@����9���h����G�Lϡ��   �   P��<���<��g<<����m��Y&)��9��%����=�N����뷿;y��a5��mW��)y��>���A������������ y���W���5���i��u8������_?�mZ��:�����*�d���L����Ke<D��<L6�<��m<🞻��켌�a��1����ӽz���F�<���������ҽ�ݣ��X_��p�� n<�   �   .'=.=L�<PX�������
4������j��^H��ʎ�5��V7�� ��P?���c�Ky��㠔����a���N������ʯ��"�d�F
@�X��5����¿����=J���|k��H6��Ӥ��s����<c=��'=��=J�< �$;�����4a�p���)�����}���CH��ƛ_�B��T����++;��<�]=�   �   R�f=�S=ƈ= ��bn�>�mL��p꾅�2�`��������⿲��^&,�p�K�2�j�����+��x���0��M���ek�4�L�|L-�"�忛���Vみ�15�ׇ�lޏ���<gz� �G��g=̑J=�d^="HL=@ =|��<��< � ��z
���&��0���$����H����tӻx�!<���<�((=�mT=�   �   F�T=h1G=X?=�/2�]h����_����徉�/��S|�5���/+߿��LN)��'H�Sf�e9���,��]Y��s'���C���f�r�H�HJ*�z���3��~���*���1���辞،�J���Xt��N��c�<L�>=p�L=�04=rC=`Jx<��A���*���H��lh��r�&f��D���仛�@舺�o�<H�	=�p<=�   �   ��=�"=	�<�����:X�	�G���Nyؾ�-&��po�g^��D�Կ|�Z!���=��Y�dPq������������f
q��~Y��>�b�!�r���)ֿN�����q�\
(��Y۾�#�����nbc���p�0r�<"=t=l��<8�
<�-Y����*�t��6��� Ž�ٽ�O�sDؽ;a½�����l����0s5�x'.<���<�   �   ���<0 �<H�<�pL��<A������i��!ľ�e�	2[�n-��#Ŀ�������TC.���F���Z���h��lm�0Hh�6UZ��E���-�.��@-����Ŀ�����\���RgƾZm�ܦ��L#K��䬻P-�<`k�<�h^<�%��j���ɀ�b�Ľw���!��F8��F�3�K�~F���6����	�����>w���`E��   �   ,�� �P: ��;�z�2�(�C3ѽ�xI�#�����MA�'7��ž���qۿ��| ���/���@���K�R�O��<K���?��.�m��H��@ۿ�v����;B������4L���ս *1�p	��r;�r��D��B�R��	��|h���=�&n�4{��P[���
���~��f���.�����j�Nn:��-	��<��n�H��   �   �愽PJ ���_�Ppk�T:�=���.�%��捾��޾T�#�~�c��:�����Å�2�j=�
%���-�r�0��H-��$�F)���8俲¼����c��3$�`�߾tێ�^�'��-����|���H|�VP������Y���1�v�T͞�ؠ�����N���.����h���I���t޾dG������%�q�Si.�����   �   f� �ҷ���n#�P�ּb�Ý��B&�Pa�iK��j:���:�q�x�θ���ο�lL������	�*������1�޽����i`޿�M�������Uw�r5:���u��xb�S&��Ί���P�"�)�����HP���J��z�������Q�t*���'���8�E�C�`G��B��7��\&����CB��)��J[��c~G��   �   RO����\��t�1�p#�"�V�½ސ)�&4��U�ξ'���E�;*|��C����̿͘Y�޿�8꿳��[�Pݿ��ʿ�a���ј��z���C������;�ֈ�Zs)���½*�X����
a5�VЙ�
��<�Q��욾�n־6R���.��O�A!m�W�&���]���������%k�ֲM���,�:�
��Ӿ����   �   ���ĆD��|���(n,���,��Έ��ｚ�E��G��Vi۾�9���@�L�m��e���@��%߭����蹿�Z������՝�^����Dk���>�H����پ���l�D�Hw����l,�d�,��҈��x�E�[K���m۾�<���@���m�5h��UC��*⭿���>빿^��︬�I؝������Hk�:�>���ێپ�   �   \�;lو��v)�G�½°X�@��&[5�˙����h�Q��蚾�i־O��.���O�Vm��e���Z��	���@��i�j���M�d�,�>�
�Y�Ӿ9���LO�0��W����1�"#�,�V�t½��)��6��<�ξï�E�V.|�F�����ߛ̿��޿+<�*���^�4Sݿ��ʿ�d��Ԙ�fz���C�Z���   �   ���w���b�V(��Њ����༘�)�Q����K�:�J��v������cK��&���'�q�8���C��	G���B�ˬ7��X&�H��W<�%��kW��}xG�� �屖�zg#��ּ�b�H����(�%Ta�gN��<���:���x�򺝿ѿ�OO�����ʧ	� ������3����"���!c޿#P�������Xw��7:��   �   �5$���߾-ݎ�r�'�}/��d��p����-|��E�E����O�f�1�v�}Ȟ�8���\��w���~*���޴��B���n޾�A������q�Rc.�q�����(A �h�_��hk��;������%��荾��޾n�#�A�c�W<������=�忢�?��%���-�f�0��J-�B	$��*�*�V:俛ļ���h�c��   �   v=B�6������6L���ս�*1�0� �r;�z����\�R�7 ���b���=��n��v��GV��[��|y��Ia���)��'�j��g:�((	�4����H�8����VR:Pַ;�s�h�(�+6ѽ,{I� ���U���NA�o8��_���zsۿ8���!�.�/�h�@���K�L�O��>K���?���.�`n��I�QBۿm򮿒����   �   
�\����hƾ�m�����$$K�Pڬ�4�<�v�<x�^<�Ы����<�����Ľ�!��?8���F��K�X�E�:�6������Sz���w��w��hD����<�)�<�<`oL�?A�����$�i�z#ľg��3[��.��}Ŀ-�������D.���F���Z�`�h��nm��Ih��VZ�r�E���-����.����Ŀ����   �   ��q� (�vZ۾�$��<���bc��{p��v�<�=�=��<�<�Y�N��Ըt��.��1�Ľ
�ٽ�Fབྷ;ؽ�X½J���x�l�����K5�G.<��<"�=Ƒ"=��<�����<X�	�.񁾫zؾ�.&�Hro�:_��I�Կ� !���=�(�Y��Qq�@���p���ɠ���q��Y�n>��!���W*ֿ�����   �   0+���1�����،�p���Xt�@N��f�<L�>=$�L=p44=�G=P_x<�#A�@���h��VwH�"dh�V�r���e�~D����خ���4��8y�<�	=ps<=D�T=�2G=�?=�S2��^h�ο�D`�����"�/��T|������+߿l���N)�V(H��Sf��9��c-���Y���'���C��f�f���H��J*����U4�%���   �   9み\15����5ޏ�:�`fz��G�"h=6�J=Le^=~HL=� =8��<p�<�����:
�H�&��0���$����X���Puӻ�!<d��<�((=�mT=�f=DS=X�= ��> n����L���꾶�2�#`��֛��������t&,���K�F�j�����+��x���0��F���ek� �L�hL-����z����   �   *���1�����׌�\��Vt�`�M�i�<�>=��L=�44=H=`x< "A� ���X��TwH�$dh�R�r���e��D����Į��@3��py�<0�	=�s<=��T=R3G=�@=��1��[h�¾�z_��d��N�/�qS|������*߿ڍ�N)�n'H��Rf�9���,���X��'��/C��8�f���H��I*���_3�c~���   �   ��q�`	(�.X۾�"��2���]c��Cp�8{�<:=�=h��<�<hY�����t��.��/�Ľ�ٽ�Fཙ;ؽ�X½P���t�l����(K5�8H.<��<�=�"=�<�R���7X�	��rxؾ�,&�!po��]����Կ��!��=��Y�:Oq�㽀����h���	q��}Y��>���!�ν��(ֿw����   �   ��\����ueƾ�|m�����K�@���|:�<�z�<�^<�ɫ�X�����\�Ľ���!��?8���F��K�\�E�>�6������Iz��vw�Xw��^D����<D-�<��<�%L��7A�C�����i�d ľ�d��0[��,��
Ŀ*���ւ�HB.�D�F�b�Z��h�*km�hFh��SZ���E�L�-�*���+��,�Ŀ����   �   �9B��������1L��ս�!1�0�� -s;@+������R�R�����hb���=��n��v��FV��^���y��Ma���)��*�j��g:�(	��3�� �H����� �R:��;pG���(��/ѽ3vI�s~�����fKA�6��i����oۿ��@� �/��@���K�^�O��:K��?�~�.��k�bG��>ۿh﮿+����   �   �1$�7�߾(َ���'�4(������ゼx|�\C�`���WO�4�1��v�pȞ�0���X��v���~*������B���n޾�A������q�8c.���Z߄��> ���_��Pk��2�㸫�l�%��䍾�޾��#��c�9���}��������;�P%���-���0�G-��$��'�d��5俕���6.�c��   �   ���q���b��"�AɊ�^����l�)�����K��J��v��p���VK��&���'�q�8���C��	G���B�ͬ7��X&�I��U<�%��bW��OxG��� ������c#��|ּVY����R#�.La��H���8�A�:�Dx�۶��,̿��I࿷���\�	�`���� 0�&�������]޿MK��ݲ��$Rw��2:��   �   ��;Ԉ��n)��½��X����U5� ə�R���Q��蚾�i־�N�ܴ.���O�Sm��f���Z�����B��l�j���M�d�,�<�
�Q�Ӿ$��sLO���V���1��N�V�	½ �)��1����ξª��E�l&|�fA��w��ݕ̿%�޿]5�C��4X��Lݿ��ʿ-_��qϘ��z�E�C�\���   �   ��}D�6o���\a,��,�̈����E��G��<i۾�9���@�G�m��e���@��%߭����蹿�Z������՝�a����Dk���>�F����پ����D��u�o��Pd,���,�Ɉ�y����E��D�� e۾7�T�@��m�>c���=��5ܭ������乿�W������ҝ�����-@k��>�I���پ�   �   �FO����P�� �1�L�ķV��½�)��3��4�ξ���E�5*|��C����̘̿Y�޿�8꿵��[�Pݿ��ʿ�a���ј��z���C������;�ֈ��r)�d�½�X�����P5�ę������Q�!嚾�d־ L�>�.�k�O��m�큿���X��Q��������j�J�M���,��
�@�Ӿ<���   �   � �-���,[#�tּ�X�����H%��Oa�?K��\:���:�l�x�̸���ο�kL������	�,������1������m`޿�M�������Uw�p5:����t���b�d%��ˊ�L����Z�)�)����F��J��r������gE�X#���'�*�8�1�C�*G��B�y�7��T&����46����LS��rG��   �   ؄��4 � �_��Dk��2�˺��l�%�G捾��޾M�#�z�c��:������2�j=�
%���-�t�0��H-��$�H)���8俳¼����c��3$�G�߾?ێ���'�+�����T���h|�T:�����8F�4�1�P�u��Þ�ȕ��;�������&�~��T��<��ch޾y<��Cz����q��\.�C��   �   �ޕ� �T:�;`7绀�(�p1ѽxI����ڟ� MA�&7��ľ���qۿ��z ���/���@���K�T�O��<K���?��.�m��H��@ۿ	�x����;B������<4L��սH$1�(���fs;�W��맼��R������\���=���m�r��^Q��/ ��6t��\���$��x銾
�j��`:�K"	�w*��X~H��   �   p��<8�<���<�L��8A�����|�i��!ľ�e�2[�o-��$Ŀ�������VC.���F���Z���h��lm�2Hh�8UZ��E���-�.��C-����Ŀ�����\���<gƾ�~m�����4K�����>�<���<ȩ^<`}�����?�����Ľ@���!��88���F���K�:�E�r�6�H���� ��p��>�v��\＠�C��   �   �=��"=H�<�6��"8X��	�+���Ayؾ�-&��po�g^��D�Կ|�X!���=��Y�dPq������������f
q��~Y��>�`�!�r���)ֿO�����q�[
(��Y۾�#��M���_c�@Jp��}�<�=�#=H��<�:<��X�b��6�t��&����ĽS�ٽ>��2ؽtP½�����ul����h"5��i.<��<�   �   @�T=25G=B= �1��[h����_����徇�/��S|�5���/+߿��LN)��'H�Sf�e9���,��]Y��s'���C���f�r�H�HJ*�z���3��~���*���1���辑،����Wt�`�M��i�<&�>=��L=�74=�K=�qx<@�@�H驼D���oH��[h��~r�Z�e���C�L��t����x��P��<T�	=w<=�   �   ,�=�`�=FpG=��<�t���t�b�����LG��Z������]ÿ����\���-�LRF��[�v&i� (n��,i��8[���F��.��������YſwT��9]���Տž�i��u콚���
M<00=�o=�4�= �p=�J=J�=쿷<P<@!{� �[�<V�������o���y9���X�H�I<Lz�<s*=>D`=k�=�   �   �!�=�|=��A=���<�)��1OڽC�]�����Hy�<V����5�������v�*���B�R�V���d��ki���d�|W��C���+�8��c���¿���B
Y����,����jd��R�4}�x7L<F�*= �d=F�p=�[=D/=<s�<)R<�y&��@����ڼ�D�\������{ɼh�V��(�:��<�N	=j4E=��r=�   �   PX=�o[=r�/=<�<���սɽsOO��i��+R�FK�?��� �����
�Ȧ"�&�8��WK���W��\��W��K� �8�v�"�dP����+[������XM��P��ҵ��JU��Խ�C�oF<Z=tE=�WA=Z=��<`xp; ǈ�(����]���m��𝡽=��X����P�j���|F���<,��<f�1=�   �   ԉ=@�"=�=@�<���4���d9���F&���n9��,��wx��d�ӿ% ���f�)��9�<�D� XH�ZD��p9��<)�&��=0 ��YԿ�:������;�� �̯��c>��"��\�⼨2<T��<��=0��<h�-<��K�h"�(�
4Ž����8���F�� ����VE����^������p����<�   �   �o;\�<��<@�C< =��� ���7�������ܾ��"���b�����0����H��$���$��-���0�0x-��5$��N��0��X��Ѽ��f{c���#���޾�錾,!�<����=��`# < �<X�k<��'��򼼬����Խ�-�Ư>�B�c�?���Y���4��r���xq}��g_���9� ����ɽZ�q��Jȼ�   �   ���i����;p#�;�4h�~d��?��F�d�$e��/�	���@��E��{���4�ſX翔y�!�z�������*P�T��Z����Ŀ��������@���	��h���(g��I���o�X[�� ��:@I;H\�f�0��K��$�
�>�E�˵��ű��[��4GϾAxܾ�ྏp۾�[;=ʷ�r�|O}���?�G��	���   �   g󻽄I>�DÌ���0�M��
(�`ܿ�Sw2�	Ӓ�b޾�l��,S�}݆�2Ƥ�D���9ڿ���P�����������쿑gؿ(���f��/腿�R������ݾ���tu3�&�½�{/�x�q�������v�L��sĽt, ���j����B�ʾ����4�z���(%��(��y$���I��B>��ƾ����Z�d��+��   �   �>"��ܾ��A��`��8%j��V켩چ�}��=]��Ī�d���,u&�lV�aۃ�g��B��J���D�ɿͿ�1ɿ%����b��$̙��z���OT��$����	���m1\��6��z����򼈌~��c���0J�7�Ľv&�:w|�	���i��M%���/��WI�B+]� �i���m�i�h�#�[��8G���-�f����ˈ��p�w��   �   c�t��D����v(�`{��hw��&+�S����]� �w�4ŵ�B����"���I�Ivo�g;��^��3�������t��q����ㆿq�l��eG��� ���������{t��@�$���
(��x��H|���#+�㳮�2b��w�9ɵ�v���"���I��zo��=�������h���]w�����
憿��l�<iG��� �����ˉ���   �   ����5\��9�~����� �~��Y���'J�!�Ľl &�lp|��������!��/�USI��&]�0�i��m���h��}[�t4G�T�-�D���羰���%�w�+:"�W־�f A�lX���#j�t]케ކ�H��yB]�&Ȫ����x&��oV��݃��i�����.���F�ɿͿ�4ɿ񥾿le��oΙ��|��<ST�� %�֮��   �   ��ݾS���nx3���½/���q����l����L��kĽ�& �v�j�!���ލʾ����81�����$%��(��u$�,����B8�~�ƾR�����d��&��뻽?>�`���P����M��(��࿽�z2��Ւ��!޾Go��/S�]߆�gȤ��F��d<ڿ���u���K��������>jؿ����"h���酿�R�����   �   N�	��j���+g�VK�"�o�\����:�;(�[��x0�C����
�R�E�����묟��U��MAϾrܾ̠�pj۾V;�ķ�ʽ���G}��?��A��������H����;`1�;P:h�X d�kD����d��g�� �	�!�@�.G��S���_�ſ�Z��z��"���.��J��Q��������ĿY��� ���@��   �   ]�#���޾9댾�!��ᙽ`?��* <x�<`l< ['�@r�j���l�ԽV'���>�:�c��:�� U���/��򅈾�h}��__�ȼ9�@����ɽ�qq��2ȼ �;\'�<��<��C<�@��c#���9���L�ܾR�"��b�b������p��r�@�$���-��0��y-��6$�(P��1��Z俅Ӽ���T}c��   �    ;�� �鰣��>�A$��� � 2<(��<n�= 
�<P�-<��K��"��苽*Žp���:���@�@ ����x?�$���u�����v��p4�$��<�=j�"=�=��<���}���U9�8���l(��Zp9��-���y����ӿ�% �����)�P�9���D�hYH�n[D�r9��=)��� 1 �[Կ�;��J���   �   sYM�>Q�Jӵ��KU�	�Խ>D��qF<H=�E=`\A=L=��<@q;l������ȳ]�L늽Fe����������P���P�nw��SF�0�<��<Ε1=@X=xr[=��/=��<`�㼲�ɽ�PO�k���R�eK����� ��"�忨�
���"��8��XK���W��\��W�� K���8��"��P�����[��/���   �   �
Y����s����jd�S�*}�:L<p�*=��d=��p=�[=/=h|�<�>R<�&�@3��$�ڼ�<����2���mɼx�V��ߪ:���<�R	=�7E=��r=�"�=�|=:�A=���<|,��uPڽ?�]�@����y��<V���m6��3��`����*��B���V���d�pli�2�d��W��C�ޏ+�z��ǹ�)¿;����   �   ]�����ž��i�?u����(M<�0=\o=�4�=p�p=J=��=���<hQ<�{��[��U��d����o���y9� �X� �I<z�<�r*=(D`=W�=�=h`�=�oG=��<Fu����b�Ђ��vG��Z������]ÿ����n���-�\RF��[�~&i�(n��,i��8[���F� �.���n���tYſZT���   �   �	Y�!��g���~id�6Q潢z��@L<��*=x�d=.�p=t�[=b/=�|�<h?R<�&�$3����ڼ�<����.���mɼ��V���:���<�R	=�7E=ƈr=�"�=�|=4�A=���<�'���Nڽ��]�>���y��;V�����5��8��Ƶ�*�*�6�B���V�t�d�@ki�
�d��W�C��+�؄����S¿�����   �   �WM��O�Nѵ�IU�r�Խn?��~F<r=E=`]A==���<�q;����p����]�?늽Be����������P���P�fw�0SF���<���<D�1=
X=�s[=��/=��<L��:�ɽ`NO�1i���Q��K�����w���B�忆�
�*�"�f�8��VK�~�W��\�ґW��K��8���"��O����AZ������   �   s;�� �/���>�E������&2< ��<t�=��<X�-<��K�h"�[苽�)ŽV���2���@�@ ����x?�!���u�����D���1�L��<�=�"=�=h�<�	�������9��򠾟$���m9��+���w��5�ӿ`$ �(��\�)���9��D��VH��XD��o9��;)�$��`/ �LXԿ�9������   �   .�#���޾�猾v!�	ܙ��/��X? <��<�l<`A'��o������Խ4'���>�0�c��:��U���/��󅈾�h}��__�Ǽ9�:����ɽRqq�H1ȼ�;d+�<��<`�C<�1������5�l��ܾ2�"�Ƴb�ɿ������A��<����n�$���-���0��v-�(4$��M�^/��V�Hм�9yc��   �   ��	��e��%g��F�<�o��J�����:��;��[��v0�oB��Z�
�!�E�����ެ���U��HAϾrܾˠ�rj۾	V;�ķ�Ƚ���G}���?��A�s��f��@� �;�\�;@h��d�
;����d��b����	���@�RD��ո��;�ſ�U�Fx��������&��N�����թĿ��������@��   �   ��ݾY���qq3��½r/���q�P���{��X�L��jĽ�& �@�j�
���͍ʾ����31�����$%��(��u$�0����C8�y�ƾJ�����d��&�<뻽�<>�d���pڮ���M�.(�/׿��s2��В�$޾�j��)S��ۆ�&Ĥ��A���6ڿ���=����������� ��dؿ�����c��P慿�R�-���   �   ����F,\��2��t�����e~�|N���#J��Ľ &�(p|�����о��!��/�QSI��&]�0�i��m���h��}[�u4G�S�-�C���羥�����w��9"�Rվ��@��M��Hj��D�mՆ��y�"9]�����>����r&��hV�cك��d������~���S�ɿͿ�.ɿM���1`���ə��x��ZLT��$�*���   �   �ut�"<����'��d��h��+�����x]�țw�ŵ�.����"���I�Evo�f;��^��4�������t��s����ㆿt�l��eG��� ���������{t�V@���T(��i���e��
+�򧮽�Y�u�w�q���f����"�1�I�ro�9�������ߓ���q������>ᆿ�l��aG��� ���������   �   �4"�>ξ���@��C��(�i�I�u؆�c|�F=]��Ī�K���$u&��kV�^ۃ�g��C��K���F�ɿͿ�1ɿ(����b��%̙��z���OT� �$����񱩾1\�6��x�����e~��F���J���Ľ}�%��i|�q��������\�/�/OI�""]�s�i��m��h�y[�<0G���-����O��H���@�w��   �   $㻽x1>�����@�����M�
(��ڿ��v2��Ғ�G޾�l��,S�{݆�/Ƥ�D���9ڿ���R���!�������쿕gؿ*���f��/腿�R������ݾ�����t3�u�½�v/�8�q����<o��@�L�YcĽ�! ���j�������ʾ�����-����� %��(�r$�m��o��2�-�ƾ䥛���d�!��   �   ���X�P?�;@r�;�h� d�{>��Խd�e��&�	���@��E��z���3�ſX翔y�!�|�������,P�T��\�� �Ŀ��������@���	��h���(g��H�N�o��M�� ��:�);��[�Dk0��:��-�
���E�����5���JP���;Ͼ�kܾ���Rd۾2P;�������R?}�%�?�I<������   �   �;�8�<p��<��C<�2��6��"7�������ܾ��"���b�����0����H��$���$��-���0�4x-��5$��N��0��X��Ѽ��f{c���#�v�޾�錾�!��ޙ��3���A <��<�-l<�&�4X�I���h�ԽZ!���>�m�c��6���P��h+��u���j`}��W_�µ9�*����ɽ�`q��ȼ�   �   �=ԏ"=�= �<8�����9���6&���n9��,��wx��e�ӿ% ���f�)��9�<�D�XH�ZD��p9��<)�&��>0 ��YԿ�:������;�� �����>��!����⼸&2<��<j�=��<��-<�_K���!�=���� Ž����`���:�� �^���9�G��l��%��$����軀��<�   �   jX=�v[=~�/=\!�<���ɽ:OO��i��(R�BK�?��� �����
�ʦ"�(�8��WK���W��\��W��K��8�v�"�dP���+[������XM��P�ҵ��JU�]�ԽXA�0}F<t=nE=$aA=:=��< �q;�������l�]�䊽�]��M�������hI����P�@k��(F��<L��<�1=�   �   $�=< |=P�A=8��<p'���Nڽ%�]�|���Ey�<V����5�������t�*���B�R�V���d��ki���d�|W��C���+�8��d���¿���D
Y����&����jd�}R�|��>L<ʻ*=l�d=��p=Ԇ[=~/=���<@RR<@�%��&��l�ڼ�5�b������_ɼ�tV� ��:	�<2W	=�;E=��r=�   �   ��=,��=}C�=�=�������p�(��\�����p1�4v����w%̿�6������#���3�, >�@�A��>�ڣ3�>$�~�������Ϳ+����-y��=4������/��HD2�;X����~���<4�V=M˅=��=$h�=��l=
B=ڻ=h�<H�o<�; �+;@�:pG�;h3<��<d�=�7=<Yl=Z��=���=�   �   �<�=���=Ⱥ�=JQ=�ύ��Ӌ��$�)��/5��3.���q��i����ȿ[G�E��!��r0�H�:�3>��:�B{0�fE!�*��J{���Gʿ)堿гt���0�v�͘���-����0.k��^�<<�R=莁=�="{=�5V=�&=��<@y<���; ƈ�\� (�@w� C����!<���<�=��O=��=i˕=�   �   �J�=���=�q=vj=  ֺP|�:���ߊ���޾��$��he�썗�UC��G�翶��ZB���'��1��J4��0��v'�47�Я���迸>������-�g�( '�e�⾼���%!��䏽h4����<�WE=�i= |e=rE=
�=��< 8;�]�|��D-�x�:��aA���2�6�����0�̻�<<��<x�<=ށs=�   �   �fL=��e=ބU=�t=�;��R�l9� �x��rɾ�
���Q��+���"����տ����3�H"�0�"�(T%��B"�������������տ�����΋�VaS�V��g�̾����X��q��ʻ�1�<z8-=�R;=B� =��<���;$��*E&��h������q̽`཰�彊eܽn�Ľ���g�����{���<8�=�   �   DH�<�=�l*=�f=P��;�� ��r޽�aT�����BC�,�8�!�v�����c����B߿"���[	������pE��������\޿�0��̃����v��9��5��Ȱ��XY�j��x:���t����< I=� �<\n<��F��ܴ��7�׽�-�k�,��PD��S�j�W�qQ�z=@�&�&����G�ƽ�b|��~开~�:�   �   `@3�h�a<�Q�<�g�<�<lؼ�ë�Х+�Z���ܾil��R��H��,*��������ٿ6�����������!��SJؿvh��a:��������Q�=j�۸ܾ2��d�.������ �g;\�<��<��;���t=^�*�ƽFm�8�G��Qy�|��������Ѯ��(��*���;�������q��2?����r���x�:��   �   �`f�0Y�� ��;!�<P�#<pk�Z�q�*��}Wb����������+��I]�5��*F���dƿA\п!�ӿX�Ͽ��Ŀ����ޞ��ۆ�G�[��*��T��e�����b�>0�`z�d�����;��>< �~:�Ǽ}|�������2�Xx��]���þɴ�Q(���D����z��i����0߾�h��A���o���*��ٽ�   �   r���\m������A;6<����V?��,���@&�Xa��̿þdc�K�.�79X�������1�������h��������:��O]}�F�U��,����D�������$������˻����; ���Ľ��n���5�dhA����������쾠b�Ь#��Q4��>�KB���=�i�2���!�m���<϶�F���Ѳ:��   �   �8�Q�ؽN�O�X�p� U>;`� ;�z���Y��"߽v�<��Ȏ���Ǿ�e�!'$�y�C���_��Xu�cz��[���{����zs�q?]��6A�q�!�I��;ľ\��x�8��ؽ��O���p�@j>;�� ;|���@Y��)߽h�<�̎� �Ǿ�h�`*$�8�C���_�O]u��|�����������~s�wC]� :A���!��K��?ľs���   �   '
����$�u������ۻ����; �����h��c-��bA����B����i_�7�#�N4��>�2B���=���2���!�[�c��ʶ�է����:����Rm�ԛ�� GA;�7<pב��E�D2���D&�"d����þ�e�N�.��<X����_���}3������#k��5��i���<��:a}���U�ҧ,�'�������   �   ���q�b��2�4fz����0��;��><@	�:��Ǽ�u���|��2��Px�Y���{þ���!��BA����2��1���S+߾�c��� ����o��*�e�ٽ�Sf�TG���
�;8&�<��#<�,k�x�q����[b����������+��L]���OH��P����ƿ�^пϪӿ��Ͽo�Ŀ�������L݆�5�[�b�*�+X���   �   ��ܾ�����.�*���L����g;@`�<���<p[�;�x��/^��ƽ�g�H�G��Iy�󰒾�����̮�r#�������������B�q��+?�v��������:�3�h�a<Z�<k�<�<dؼ�ǫ�Ĩ+�>\���ܾon�]R�IJ��,������ڱٿ�8�5�������t�����뿏Lؿrj��<��򸅿ڞQ�l��   �   7�Zʰ��ZY�K�齈:���t���<jL=�+�<h|n<���T��<����׽(���,��ID�9S��yW���P�^6@���&�4��b�ƽ
R|��c开ȫ:pW�<(�=�o*=�g=p��;� �6v޽SdT������D��8���v�q�������D߿L
��]	�������F����%���Y^޿o2�������v���9��   �   S��ͻ̾q��Z���q��ʻ|3�<�:-=�V;=� =D&�<�(�;�����6&��`������g̽�U���![ܽ��Ľ᧠���g��������<��=\lL=��e=چU=�t= �;��R�;���x�Ktɾ;�d�Q��,���#��^�տm���4�J#�D�"�>U%��C"������������տ�����ϋ��bS��   �   � '�X��] ���!�w叽`4����<BYE=�i=�e=xE=p�=���<��8;��\� �㼠 �@�:��TA���2�ʎ�����S̻8�<<���<n�<=��s=�L�=٬�=$�q=Vj= Oֺ"S|��������!�޾��$�je�����>D��W��R��C���'��1�ZK4���0�Zw'��7�Z�����t?��H����g��   �   !�0���B͘���-����P.k��_�<&�R=���=늆=�${= 9V=�&=D�<@4y<ช;����8B� �'�pD� B���"<h�<�=��O=�=�̕=�=�=c��=���=�P=p؍��ԋ���$��)��6쾄4.�D�q��i��-�ȿ�G� F�H!� s0���:��3>�\�:��{0��E!�l���{��CHʿj堿2�t��   �   m=4�B���[/��D2��W���~���<��V=w˅=�=Jh�=�l=VB=8�=	�<x�o< �; �+;���:pH�;�3<0��<h�=Ԛ7=4Yl=V��=v��=��=��=TC�=v=p��������(��\�����p1�hv����%̿�6�����#�ȇ3�4 >�@�A��>�ң3�4$�r�o���j�Ϳ���Y-y��   �   G�0���a̘���-�G
��p%k��b�<<�R=��=9��=%{=�9V=&=��<5y< ��;���� B���'� D� >���"<��<=��O=�=�̕=�=�=���=e��=RR=0ȍ�9Ӌ���$��(���4쾰3.�/�q�Ki��X�ȿ�F�jE��!�Zr0��:��2>���:��z0�E!�Я��z��eGʿ�䠿�t��   �   1�&���⾳����	!�^⏽X�3�`��<R[E=�i=؀e=NE=�=Ժ�<`�8;�\����t �"�:��TA���2�������S̻��<<4��<��<=�s=�L�=`��=ԭq=�l=��պ@M|�N���ފ�Ң޾,�$�he�b����B��q��6���A��'�*1��I4�8�0��u'��6�2������=�����g��   �   ����̾ؑ��V��q���ɻ�;�<�=-=�X;=�� =�(�<P0�;L���6&�N`��f���g̽nU����[ܽ��Ľۧ����g������ �<&�=NmL=�e=.�U=�x= ?;D�R��7�$�x�qɾ	
�~�Q��*���!����տW���2�V!�*�"�S%��A"�����������տ]����͋��_S��   �   b4�xư�oUY�Ę�8:� 's�Ԫ�<�O=�0�<��n<@��B��ɫ����׽�'���,�tID�.S��yW���P�Z6@���&�-��I�ƽ�Q|�$c开ݫ:�Y�<��=�r*=�k=��;&� ��n޽ _T��B���8�v�����⳾��@߿"���Z	�������6D���������Z޿*/��U���S�v��9��   �   ��ܾ�|���.��������� Oh;�j�<H��<�p�;�t���-^�Q�ƽBg��G��Iy�尒������̮�n#��
�����������;�q��+?�`��m���"�:�H3�(�a<<`�<�t�<H2<��׼������+�#X��ܾ�j��R�OG��~(������P�ٿ�3����o��C������Hؿ\f���8��﵅��Q�1h��   �   N����b��,��Uz�����)�;��><���:��Ǽ�t���{齽�2�aPx��X���{þޮ��!��@A����0��2���P+߾�c��� ���o� �*��ٽ�Rf�tC���#�;�/�<$<� k�R�q�7��|Sb�������+��F]�w��&D�������ƿ�Yпz�ӿ��Ͽp�ĿH���ܞ��ن��[�o�*�vP���   �   �����$�1�����0���`/�; \�|����g��{,�lbA����'�����a_�0�#�N4��>�2B���=���2���!�Y�^��ʶ�ʧ��b�:���&Pm�ȕ�� �A;�S<����86�!'��=&��^��P�þ$a�~�.��5X����ⓑ��.��y��� f��)�����V8��9Y}���U��,�x��p����   �   F�8��ؽ��O�P�p� �>;�C!;dq����X��!߽�<��Ȏ���Ǿ�e�'$�r�C���_��Xu�dz��\���|����zs�r?]��6A�q�!�I��;ľK��;�8��ؽ<�O���p���>;�Q!;i����X�q߽��<��Ŏ���ǾTc�$$��C��_�nTu�x�����)���$vs�S;]��2A�:�!�nF�o7ľ�����   �   ���&Dm����� �A;�Y<P���>;��+��}@&�0a����þZc�B�.�09X�������1�������h��������:��P]}�E�U��,����7������÷$����f������P/�;  ޸t���|b���$�C]A�Z|�����Ĩ�Q\���#�AJ4��>�B���=�ǽ2���!�/���Vƶ�$�����:��   �   Ef��/���V�;�6�<8$<�	k��q����"Wb����������+��I]�3��(F���dƿC\п#�ӿZ�Ͽ��Ŀ����ޞ��ۆ�E�[��*�T��R���c�b��/� ]z�����#�;г><�$�:��Ǽ�n��as�8�2�jIx��T���vþ6�⾻���=�J��������%߾�^��������o��*���ٽ�   �   8�2���a<j�<Py�<2<,�׼w«�^�+��Y���ܾbl��R��H��+*��������ٿ
6�����������#��UJؿwh��b:��������Q�:j�θܾ��
�.�ܐ��|��� 8h;$m�<��<���;�a��n ^���ƽ�a���G��Ay�����񣾞Ǯ�@��𝭾������E�q��$?��}�4�����:��   �   $j�<��=Fv*=�m=��;н ��q޽.aT�����:C�(�8��v�����d����B߿%���[	������rE��������\޿�0��̓����v��9��5��Ȱ�TXY���齚:� �s����<^R=$:�<H�n<���\������ʕ׽*"�,�,�fBD��S�rW�f�P�6/@��&�O�� �ƽ�@|�tG开:�:�   �   (sL=4�e=��U=�y=@7;��R�9���x�lrɾ�
���Q��+���"����տ����3�J"�4�"�(T%��B"�������������տ�����΋�VaS�U��\�̾e���X��q� �ɻ|;�<D?-=<\;=�� =|6�<�x�;�刼�(&�gX�����]̽0Kཉ���Pܽ��Ľ�����~g�R����$4�<��=�   �   �N�=���=t�q=�m=��պ�N|� ���ߊ���޾��$��he�퍗�VC��I�翸��\B���'��1��J4��0��v'�27�ү���迷>������,�g�( '�`�⾰����
!��㏽ 4����<\E=�
i=��e=�E=��=�Ƞ<`%9;��\�X��\�nz:��GA���2�p���� ̻��<<d�<��<=��s=�   �   �>�=`��=Ề=�R=�Ǎ�iӋ�З$�)��*5��3.���q��i����ȿ\G�E��!��r0�J�:�3>���:�B{0�jE!�*��I{���Gʿ)堿ѳt���0�u��̘�n�-�[��8*k�b�<j�R=d��=㋆='{=<V=N&=��<PGy<��;pf�� *�(�'�`� R���%"<l�<V=J�O=��=�͕=�   �   ��=3��=Ꞣ=��j=�/�<^V�:\�K�\�fӶ�n�	�q�A�!���գ��_ǿ�����'��������8�&-�4�@Xȿ� ��hL��V\D�\������i�����p&F�`<b;�8=��l=6�=�֐=M��=�=>�^=H�;=PF=`<�<l��<���<��<��<hV=V(=�>R=�=~�=@0�=���=�   �   4>�=-��=/c�=j=�L�<������ٽn�W����P��8>���}�+���!Ŀ;�忊�����0���7�҄�:��v���N��Ŀ(��R����@�a�	����� d��r���=�P1�;N�=��i=�
�=2Ћ=7��=�l=f,H=�� =<F�<��<�H�<�Z<X-\<��<Hz�<��=�W2=�Gd=
�= b�=X8�=�   �   p�=Rx�=	u�=`�f=�	�<�Uм��ƽ��H�{8�����a4��p�T%��A�����ڿyN��z���=�@���&�:���=��	ۿk,���ᙿ=kr�6����O���T�w2��"�`�;��=n�`=�p|=d�x=8�^=&5=`�=HO�<�v�;�R��`TC�D�� 艼�UV��)��0_�;X4�<\�=yM=Á�=|��=�   �   V�=�G�=|(�=��_=h�<� ������\�1�C��_��!$��9\����9ɫ��ɿ���ק������,�P��%'���x㿩\ɿ�ԫ�i쌿OF]�m�%�AP�%���$;�`^���j��8J<=��O=b�Y=�C=@=�< �0;�(��,�
���J���{��/��� ����db�t�$�8'���8��L��<bP =J�c=�   �   N�:=Bj=r�t=|�R=|��<� �����;Ɓ�j�Ⱦ����B��y�բ������-˿�ݿ�h�aG���过�ܿ�bʿ�ಿ�>��1�x��aB�Y|�D�ʾ8y������W��|���ئ�<d=g4=xL%=��<Л<�g�|&����������"�b�
�����.����Z5߽�g��4r_�@ϼ�X#;\�<�   �   ��<�l=�@=:�;=��=�[;�M9�A���AS�־��,��bm$��7T�/���O9���宿K���(ɿ�u̿=�ȿ�"���⭿�G�����CS�W�#�d���o��V�8����Q�������<d�=��
=ԃ�<�N�:�1޼�|�Rͽ�_���6��Y���t�Ă��+���H����n��Q�Z�+�ְ�����*A�8H��   �   �����<(b�<��=2�=��;<`/Ѽ�?���z!�ʃ�������q�J�-�cW���~�� ��:����;��_���>���q���a叿�|�� U��,��Y�����1悾��!����ȗ�`��;�)�<p{�<�< �����9��"���]^6��/p������j`��=�̾2<о�˾�v���˨�����H�d��)�>���U��   �   �>��h���B<do�<�;�<���<�𻜵M�+���B�8Ó�Ȓξ$��a�)��J���f�K.}������߇��%��p{��d�үG�A'�����C˾K%���?�#޽�sI�P� ��-�<���<`s�<��x:� �9����	��N�kl���)��t�۾T���UY����e����`�
�������־Pϯ�,����C������   �   \���Lh��L$��X�-<���<��<h�<�T��L'��E��4S�8L��A�ɾ��������/��<A��[L���O��}K�,�?��e-���7���iAž����4TK�����b��4����-<H��<��<؄<Tc���,��5���	S��O���ʾ�������q�/��@A��_L���O���K�¡?��h-����/����Ež����:YK��   �   �?� )޽�{I�@� ��)�<Ć�<�y�< z:�������=�	�
�N��h��m%��H�۾����.V�����a�o��L�
������־˯��򇾈�C�R����8��4��HZ<�u�<=�<H��<���M�b1�X�B�9Ɠ���ξ���O�)�1J�u�f�Z2}�����⇿�'�� t{���d�
�G��C'�>��YG˾(���   �   _肾��!�Tũ�@�� ��;�)�<��<x��<�+��������w��nX6��(p�����묾K[��߅̾�6оa˾�q��QǨ�����]�d�_�)���~G�����(�<�k�<�=�=��;<�:ѼqD��/~!�.���� ¾�s���-�yW�t�~����U����=��� ��h���}���C珿h�|�p#U�,��[�����   �   r��+V�g��0R����L�<��=* =���< `�:�޼�|�ͽfZ�&�6�đY�կt�ￂ�c'���D���n�zQ��+�n���򰽮�@� �G��,�<�r=�@=��;=�=@*;�S9����:ES�B���n��yo$�k:T�����;��z箿^���*ɿ�w̿[�ȿ�$��l䭿AI�����BFS�;�#�P���   �   >�ʾ�z������Y�������<�d=�i4=�P%=@�<x�< og�4n&�/~��6������
��	������,���*߽6^���a_��μ�	$;�-�<��:=�Fj=�t=>�R=h��<�� �������ǁ���ȾB���B�Vy�>�������}/˿�ݿ�j�aI����`�ܿ:dʿ$ⲿ@��V�x�HcB��}��   �   �Q�-&��J&;�f`��do���J<|=l�O=l�Y=C=,F=�+�<�1;8����
���J���{�^'��������<�a���$�����ǡ����<LX =��c=��=,I�=V)�=,�_=���<x&��4���U�1��D��]�9#$�s;\����hʫ�<�ɿs��r���f���-�"���(��(z��]ɿ�ի�K팿�G]���%��   �   E�����T��3ཪ�"���;��=��`=�r|=b�x=>�^=\5=�=T^�<���;`���*C�d.��҉��*V� ح����;<E�<��=:M=N��=y��=�q�=Iy�=�u�=\�f=��<�Zм��ƽS I��9������a4�_�p�&��!�����ڿ�O����*>����'�����>���ۿ'-��+♿6lr��6��   �   ��	������ d�s��v=��/�;��=L�i=&�=�Ћ=:��=��l=�/H=r� =�N�<���<0S�<X�Z<�B\<���<P��<F�=�[2=lKd=��=6c�=H9�=�>�=���=\c�=�j=�J�<؊���ٽf�W������49>�e�}����7"Ŀ�����������
8�"��������IO�m�ĿK(������@��   �   �[�ҙ��n�i�+����%F��Bb;9=�l=56�=�֐=k��=	=��^=��;=�F= =�<��<,��<h��< �<�V=l(=�>R=�=��=:0�=���=��=$��=̞�=L�j=�.�<W��\ར�\��Ӷ���	���A�8���գ��_ǿ�����'��������8� -��3�+Xȿ� ��TL��1\D��   �   �	���c�q��� =��?�;��=Z�i=��=Oы=���=0�l=0H=�� =�O�< ��<�S�<��Z<hC\<���<x��<Z�=�[2=�Kd=��=Ic�=l9�=?�=޼�=�c�=
j=DN�<����A�ٽ�W�����Q8>�C�}����f!Ŀڿ�N��z����b7�~�����(��MN濓�Ŀ�'������@��   �   ��'����S�0�N�"��7�;t�=��`=Xt|=��x=N�^=B5=�=�_�<��;����)C��-���щ�(*V��֭����;�E�<��=zM=q��=���=�q�=�y�=Bv�=��f=�<�Pм�ƽ��H��7�������4�4�p��$������	�ڿ�M������<����X&����{<��ۿ�+�������ir� 6��   �   3N꾃#���";�![���`���'J<N!=R�O=��Y=� C=�G=x.�< /1;\����
���J�*�{�1'������칅��a�j�$�8������<��<�X =�c=�=�I�=Z*�=4�_=$	�<���3�����1��A����� $�n8\�,���7ȫ���ɿ���U�������+�z���%��Dw�M[ɿ{ӫ�b댿�D]�%��   �   ��ʾvw��$���S��������<vi=�l4=tS%=��<x�<8ig��l&��}��Ǖ��b�c�
��	������ ���*߽^���a_�\�μ�$;�.�<��:=Hj=z�t=�R=l��< � ��섽����ā�u�Ⱦl��KB��y���������,˿9�ݿ�f�gE���迣�ܿ�`ʿ߲�d=����x��_B��z��   �   ^m��XV����X�Q�����<�<�=�=@��< ��:�޼~�|�XͽZ���6���Y���t�⿂�Z'���D����n�nQ���+�Z��v�*�@�@�G�/�<6t=F@=� <=*�=`�;�F9���轐>S�����K��k$��5T�ˮ���7���㮿P����&ɿ�s̿�ȿ� ���୿�E��(�MAS�:�#����   �   �ゾӯ!�v���,��p �;�7�<(��<��<�ξ�¿�����v��X6�p(p�����묾<[��ԅ̾�6оZ˾�q��KǨ�����L�d�I�)�����F�x���0�<4q�<�=2�=��;<�Ѽ�:��xw!����������o��-��W���~����1����9��-������Z���o㏿��|�wU�	,��W������   �   �?��޽�hI�8� �=�<���<���< �z:���{���̔	��N��h��L%��-�۾p���(V�����a�m��J�
������־	˯���n�C����8��� ���d<�}�<I�<�<П𻸫M��$㽒�B�a����ξ�����)��J��f�\*}������݇��#��l{�.�d�w�G�&>'�����?˾/"���   �   `���m\�����H�-<d��<0#�<��<(N��&������S�L���ɾl�������/��<A��[L���O��}K�+�?��e-���1���`Až����TK�t���Ab�������-<L��<<$�<8�<�A��;!��J���R��H���ɾ���������/�G9A��WL��O��yK���?�Bb-��|�����=ž)򒾨NK��   �   1�����`<`��<�K�<��<p��ȲM�*㽀�B�Ó���ξ��V�)��J���f�J.}������߇��%��p{��d�ӯG�A'�����C˾;%���?��"޽�qI��� �|7�<��<<��<�8|:���|�����	�FzN�,e��!��A�۾����S�b��c^�)��,�
�#�����־�Ư����C������   �   �p��x�<�{�<�=Է=��;<�(Ѽ�>��^z!�����l����q�@�-�]W���~�� ��:����;��_���@���s���a叿�|�� U��,��Y����悾V�!�O�����켠��;6�<$��<�<�������C��n���R6��!p����C笾@V����̾W1о˾�l���¨�e�(�d�X�)�<���7��   �   �@�<�z=v@=�<=B�= �;K9�S��oAS�������Zm$��7T�-���O9���宿M���(ɿ�u̿=�ȿ�"���⭿�G�����CS�V�#�]���o���V������Q��޹�x�<�=�=d��<���:�޼ġ|��ͽ�T���6���Y���t�ѻ��1#���@��)�n�6Q���+�ͥ�,鰽�@�дG��   �   ��:=�Lj=��t=`�R=���<0� ��B��Ɓ�S�Ⱦ����B��y�բ������-˿	�ݿ�h�dG���迉�ܿ�bʿ�ಿ�>��1�x��aB�X|�<�ʾ(y������V������|��<�i=�n4=2W%=�!�<��< @g�`&��u������
��
���������\���߽�T��Q_�h�μ��$;�@�<�   �   ��=�K�=t+�=*�_=��<@��脩��1��B��N��!$��9\����:ɫ��ɿ���ڧ������,�P��)'���x㿩\ɿ�ԫ�i쌿NF]�l�%�:P��$���$;��]��Pg�� !J<!=l�O=,�Y=�$C=,M=�<�<��1;����"�
���J�~�{����f������a���$����J�� ��<�` =��c=�   �   rs�=�z�=�v�=,�f=��<Sм3�ƽ��H�l8������]4��p�T%��B�����ڿzN��z���=�B���&�:���=��	ۿl,���ᙿ=kr�6����I��zT�&2� �"� ,�;�=&�`=�u|=�x=��^=� 5=(=Xm�<���;p���pC�D������@ V�p������;tV�<H�=��M=��=Đ�=�   �   �?�=r��="d�=zj=hN�<H�����ٽV�W����N��8>���}�+���!Ŀ<�忊�����0���7�Ԅ�<��v���N��Ŀ(��R����@�a�	����� d�sr��\=��7�;��=|�i=��=�ы=H��=D�l=�2H=�� =�V�<p��<�\�<@�Z<HW\<���<��<Կ=�_2=Od=0�=�d�=p:�=�   �   b��=F�=��=G��=J�==�>8;v%p����Ѫ���ɾ��}D���{�J]��2���^�Ϳ��{I�[��XJ���-ο0��b	���f}��(F����!о,��|J$������㿼T'�<�(=�e=vف=<��=!>�=��t=��`=v�K=2Q9=�
+=��"=t�"=2�*=�;=N$U=��u=ۍ=��=|��=z��=�o�=�   �   Z��=���=5$�=�v�=��?=�7�;�7f�h����}��ž�S�o@��Gw�����趲�	�ʿ3Uݿ�_�W��MX�7Yݿ�ʿ���wV����x��wB������˾�������ួ�ï�,��<�>*=زd=.�=RN�=:fz=Zg=�fO=&7=n!="�=�G= ==*�
=0�=f�6=�ZY=���=v��=���=�ܾ=���=�   �   ���=�w�=}�=���=��E=��<wI�v��2�l��#��4^��56�݆j�D$��-쩿������ҿ_޿t��1�ݿpҿŢ������}����k�a�7��]��=����y�B���6��܈��,�<��.=R�`=��s=�Yo=�c[=*�==��=4�<\̭<��p<�](< <�i!< Hj<�D�<\B=V3=
h=�_�=gY�=�l�=�   �   �b�=N��=�M�=a �=<�L=�Ae<��#�2�R����J��@&�9�V��,�����y0������>̿��ϿU̿�c��ిd뛿�3��`�V�'�����W����p]����$�c�������<,4=z�X=@]=��I=�7%=���<�~< ;��(������.�������ݼ q���
����+<��<�/7=*�x=.��=�   �   ���=�[�=!�=^�=<�S= 2�<|s˼�Ƶ�`�1��r��!DԾ���<��i��Z���R��*��W���ӯ���C��#����Ĝ�Iቿ�i���<����X�վ*𒾮9��4˽�����];0A�<�_7=�PI=�5:=�*=H�<�%;d������Hj��,��ǰ��I�����xk������s�V{�x^x�X5<p��<�O=�   �   p2*=4�k=}O�=��=��V=�<�Z%�nf��%�8�l�ߺ������u��J�F�Z4l�����r���E����d��\���풿2ⅿ��j�T�E��:��f����?n�&�$F��`k���:r<�{=�R5=��/=�9=4��<��ֻx��ɘ��`���r�����^*��96�*�8���1���!�	���׽@ڕ� %�8����<�   �   Ȉ0<��=��P=(h=�CS=��=��;HW$��Dν��6�����ľ[��;@"�)�A��]�uFs�́�����������q���[���?�Ol � ��"¾� ��n�4��fν/�@Ӊ�d��<�O"=j�*=�	=�Ȃ<ț�H>-�r����P���R)�)�S�Qgy��H���B�������L���e���n��EE���5�ӽ��v������   �   `�ܼHx<�B=(k==�OG=b!=Lΐ<����OÅ����^gQ�|_���ȾQ��\�ɟ.��G@��iK��N�w�J�a�>��,�3��A����$ľa����I��_���z�Ȍu�<ي<,�=l�+=�=��<�ɻft-��β� ����I��u��[���3��ܮϾ�yܾxJ���ھ:4̾�1�������lx�6:�x��'葽�   �   �,��P�Ǽ�i*<~�=��1=a+=���<��c;2��6᧽|��+X��J��(�����~V��ù�l�����}� ��3޾������K�*)��&��ܚǼh�*<�= �1=^`+=��<@.c;���1秽��1X�N��4��`��(Y���ʼ�o���������n8޾v��N��
�K�(-��   �   �f��z�P�u��Њ<*�=j�+=�=4�<pyɻRj-��ǲ����H�I�&r��[���n/����Ͼttܾ?E�ޭھh/̾�-�����;fx��:��	��Dᑽ�oܼ@�<�G=n==�PG=!=ǐ<x��ȅ�;���kQ�}b����Ⱦ�U�����.��J@�-mK���N�ɡJ���>�Т,��������r(ľ>����I��   �   �4��kν
/��d��p��<O"=��*=�	=�ӂ<x{�43-�.����G��7M)���S�`y��D��x>��r���H��b����m�[?E�K�$�ӽH�v�������0<�=��P=0*h=�CS=��=`�;B^$��Iν@�6�k��M�ľ^���B"���A�%�]��Is�����[���p!��/�q���[�A�?��n �� ��%¾�"���   �   ;Cn����I���t��80r<�z=4S5=�/=�==̩�<�ֻ"������wW���h�����W*�Z36���8�T�1�l�!�&�	���׽�ѕ��%�h��,��<d9*=4�k=	Q�=˹�=X�V=��<pl%�j�����l�a�������z����F�$7l�>������ ���Lf���]��}�ㅿ��j���E���6�󾲎���   �   ���9��7˽�����];�>�<`7= RI=z8:=4/=8�<��%;⎼���Jj��$��཰��?�������a���
���s�Dl��*x�Pa<P��<�O=6��=j]�=F	�=t^�=��S=L-�<0|˼mʵ���1��t���FԾ����<�A�i�\��XT���+���m���eE������Ɯ�}≿�i�[�<�4��v�վ�   �   ����nr]�������c���뻜��<4=h�X=B]=,�I=`<%=��<x�~< �; �(�����Lv鼪�� ����ݼ0W��૤�P%,<p��<�77=��x=���=~d�=���=�N�=� �=f�L=9e<��	&�d�R�����W��&�ւV��-�����1��P���C@̿I�Ͽ�̿e��;᰿c웿�4��� W�7'�K����   �   h>��.�y�% ��7��������<z�.=��`= �s=�[o=zf[=$�==n�=�$�<ڭ<8�p<�~(<�><��!<�jj<8U�<�I=<&3=
h=�b�=|[�=,n�=���=�x�=��=Ƴ�=�E=��<zI������l�)%���^��66��j��$���쩿����~�ҿW޿m��!�ݿ�pҿ�������1~����k�%�7��^��   �   E�˾�����8➽ů�h��<�>*=$�d=��=�N�=�gz=dg=fiO=)7=�"!=�=�K=xA=��
=v�=|�6=�^Y=P��=���=���=�ݾ=���=���=F��=h$�=�v�=X�?=�-�;�9f�%����}���žhT��@�tHw����[�����ʿ�UݿL`�ڂ��X鿨YݿW�ʿH���V���x�BxB�=���   �   ~!о�+��LJ$�z���L㿼�'�<&�(=2�e=�ف=P��=:>�=Ҙt=�`=��K=�Q9=B+=�"=Ɣ"=p�*=N�;=�$U=�u=ۍ=��=���=���=�o�=`��=
F�=��=(��=��==�58;<&p��������V�ɾ��D�Ө{�\]��E���n�Ϳ
῁I�]��UJ���-ο�/��S	���f}��(F�ɜ��   �   +�˾���������������<�?*=N�d=��=LO�=�hz=g=jO=�)7=d#!=f�=�K=�A=ĳ
=��=��6=�^Y=Z��=��=���=�ݾ=���=��=���=�$�=w�=��?=P>�;�6f���2�}���ž�S� @�WGw�s���������ʿ�TݿO_�ׁ��W鿵Xݿw�ʿ���V����x�RwB�����   �   O<���y�����4�������
�<B�.= �`=ܒs=�]o=�g[=f�==��='�<�ۭ< �p<��(<�@<8�!< lj<�U�<:J=j&3=Fh=�b�=�[�=`n�=��=2y�=��=���=��E=X�<^tI������l�%#���]��46��j��#���멿�����ҿv޿���<�ݿ'oҿ���1���|����k�^�7�']��   �   ����.n]�����ғc����h��<�!4=��X=�D]=x�I=`>%=���<��~<��; �(�󪼨t������Ȍݼ�V��p���p&,<���<�77=�x=��=�d�=5��=�O�=��=*�L=HOe<� �J �X�R�ż�����+&��V��+�����d/��ָ���=̿��Ͽ̿�b���ް�N꛿�2����V��'�v����   �   M�|9�u0˽���^;�J�<�d7=�UI=�;:=�1= �<@�%;<ގ�����	j��#��g����?�������a���
��ºs��k�0)x��b<,��<2 O=���=^�=T
�=�_�=$�S=�:�<�h˼�õ��1�Lq��BԾ���u�<���i��Y���Q���(��͏��@���BB������<Ü��߉��i���<�H���վ�   �   �;n�)��A��<]���Rr<x�=DX5=�/=XA=���<��ֻж������V��,h������W*�*36�s�8�8�1�R�!��	�Ӷ׽~ѕ�%�X�����<l:*=��k=2R�=}��=`�V=8#�<8B%��b�������l�������������F��1l�<���ۊ�������b��UZ��8쒿����-�j��E�����ɉ���   �   t�4��`ν��.� 爺��<�U"=��*=	=�ڂ<`o��0-�����F���L)�V�S��_y��D��b>��`���qH��b��m�m�G?E�2��ӽƭv�H�����0<��=�P=�-h=�HS=2�=�C�; O$�/?ν �6��
���ľy���="���A��]�4Cs����ѹ�������q���[���?��i � �r¾	���   �   \X����y��hu���<��=��+=�=@��< _ɻxg-��Ʋ������I��q��1���L/��۩Ͼbtܾ2E�ӭھ_/̾�-��	���$fx��:�\	�������mܼ8�<"J=Vq==�UG=X!=ܐ<押轅�V���bQ��\����Ⱦ�L�����.��D@��fK���N�!�J�0�>���,��������!ľD ����I��   �   �����Ǽx�*<.�=x�1=�f+=��<@�c;D���ߧ���B+X�xJ��������rV������k�����}����3޾���
��ȽK�)�L&��P�Ǽx�*<"�=��1=g+=l��<`d;����ڧ�K�n&X�eG��5�����S�9�ȶ��h�����z�X� /޾v�����V�K��$��   �   �Wܼ`�<�O=�t==WG=�!=\֐<����
�O���fQ�K_����Ⱦ�P��N���.��G@��iK��N�v�J�_�>��,�0��:����$ľT��m�I��_��b z�ȅu�xފ<4�=^�+=��=h��<�.ɻ�^-����������I��n��h����*���ϾWoܾ
@ྻ�ھ�*̾
)�����D_x��:� ���ّ��   �    �0<*�=��P=40h=�IS=�=�)�;�T$��Cν(�6������ľK��/@"�"�A���]�sFs�΁�����������q���[���?�Kl �
 ��"¾� ��J�4�'fν�/�@�����<�T"=��*=�	=<�<�R��&-�d���>���G)�9�S��Xy��@��P:��4���RD��^��,�m��8E������ӽ��v�L����   �   �A*=��k=�S�=j��=��V=X �<�O%�ce�����l�����|���j��C�F�X4l�����s���E����d��\���풿2ⅿ��j�S�E��4��[����?n����E���g���Er<�=rX5=ڼ/=�D=к�<`Sֻ|������N���^��4���Q*��,6��8���1�9�!�o�	�ì׽�ȕ�p�$� ���Ț<�   �   t��=!`�=��=�`�=�S=�7�<<o˼1Ƶ��1��r��	DԾ���<���i��Z���R��*��X���֯���C��#����Ĝ�Iቿ�i���<����T�վ 𒾍9�;4˽<��@�];`G�<�d7=�VI=>:=�5=�+�<�-&;�ʎ�����i��������R6�����4X�������s��\���w���<��<�'O=�   �   �f�=���=�P�=F�=�L=Je<6�h"���R�𽧾:��8&�6�V��,�����{0������>̿��ϿU̿�c��ిf뛿�3��_�V�'�����O���}p]�����F�c�`��H��<x!4=�X=JF]=2�I=^B%=p��<( <�@;@�(��ܪ�`\�"��l���rݼT=��0K���P,<���<�?7=��x=��=�   �   l��= z�=#�=���=��E=�<vI�F���l��#��.^��56�݆j�C$��-쩿������ҿa޿u��1�ݿpҿŢ������}����k�^�7��]��=����y�,��o6�� ����<��.=N�`=ғs=>_o=lj[=��==��=H1�<��<��p<P�(<�`< �!<Ȍj<�e�<�Q=&-3=8h=%e�=�]�=p�=�   �   ���=���=%�=Kw�=��?=�<�;7f�P����}��ž�S�m@��Gw�����趲�	�ʿ4Uݿ�_�X��OX�8Yݿ��ʿ���wV����x��wB������˾}������ួ�¯����<�?*=N�d=6�=�O�=�iz=�g=�kO=�+7=(&!=��=tO=lE=��
=|�=^�6=(bY=���=n��="��=�޾=� �=�   �   `@�=���=�D�=A�=�7�=�z=�~d�+���
'��K����̾�=���7�U�c�8��T���ߨ�c[������2[��[먿$5��ŉ����d��a9��h��Ӿ����=��Tڽ�I�`���g�<�o=�]3=rD=YH=�E=0�>=�J9=λ5=�]5=`�8=B;A=v�N=�a=�y=��=���=~��=ի�=s��=�}�=B��=�   �   H6�=��=��=ğ�=GȌ=xE=xJH��S����"��I����ȾW�
�W~4�/�_�sބ�]i��G ���S������oN�����s���Z ����`���5���f�ξ%7���)8��(ӽ<Q?�0|黰�<��=~�4=wC=�E=6?=\6=H�-=& '=��#=��$=@�*=j�6=T�H=��`=�f~==�^�=F��=��=t �=��=�   �   ���=6�=��=���="1�=
�=����Ő�"}����������*��T� |�5������<���4���p����������b<|�k�T�O�+��i�����B���v�)�T��`!���캐ں<�y=S7=�?=�:=��,=X�=��	=�c�<��<�9�<x{�<��<�B�<F�=l6=,]=4t�=�I�=\|�=�N�=z��=�   �   \�=8�=�y�=�]�=���=��)= 4�9>=c����	b��z���I�Ny��A��f�먃����ճ��Tv������CG��Em��EPf�[�A�#���V���"m��� ŝ����p,�;���<2�%=x�9=L�7=8�&=Z=}�<�U�<�.<Я�;@ �����ः�@��� 
�;�d<HF�<��=�X=�5�=$��=/˹=�   �   W�=��=l�=�Y�=DP�=��;=`�<��#�%p׽<�?�w ����ξ���8*�P:K���h�������}���ֆ���~��g�UjJ���)�����Ͼ�锾�G����h��5X�X��<�r= �2=X,9=Rm(=�=0[�<@2<���Y��X$���$�΀@��8L���E�8�+����������C:��<��=L�f=s̒=�   �   ���=�s�=��=5��=�َ=�M=��<����|�����Ar��9�����y���;,���E�`eY���e��#j�qe��cX�J=D�v�*��k��|� ���?q��(�{����;� �M;(��<h�)=�-== 2=�(=�U�<���;HF�����~l�^`������ڽ���0�罭lٽd载	��4�O��5м �9�z�<��==�   �   6i=�Tk=��=i�=�@�=�HZ=���<��ɻ0�Y�<Q潆�<��舾Vٷ�v�辫�Z!�<�1��<�:q?��d;�XV0��W�A�	��[������t�6��߽6�X���'���<��=�;B=.�A=8t!=���<p�;x����F��ġ�eR�)���,)��-=�l�H���J���B��\1�u��DH�����B�F���|���h<�   �    �<=D[Y=6F�=���=��`=:�=�`<|������I�	�w$N������ȳ��پ�W����
�/����	\�OH	�^���1"Ծ���z����@�����j���h���(S<B=��G=V�T=,�===0�6<�����R�N%��f���4���_�F���.Q��:=��z���pȗ��t��lw�D/M�x����޽h>��,�˼�   �   ��ټK<J=VXN=�i=
D_=��/=�η<�ܻLE5�w��� �<K�6���.ؠ�u���m�ξ1X۾3 ߾UپI�ʾ�鴾/���|�v���8�N���\�����ټ�g<@O=�[N=�i=:D_=�/=�Ƿ<�?ܻ�M5��|�����@K�2����۠�n�����ξ�\۾�߾�Yپ��ʾ������l�v���8�>�����   �   �������x�R< >=<�G=��T=�==�= �6<����.R����N���4��_���M��^9���|���ė��p���w�Y)M�d���޽�7��p�˼p�<F%=�_Y=�G�=N��=N�`=�=�O<���Ж����	��(N�t���̳��پ�[��(�
��1�����^��J	�����&Ծ\���4����@�د���   �   8߽^�X��(�$�< �=::B=H�A=�u!=`��<0A�;,�����F�b���TJ�h��H')��'=�.�H�R�J���B��V1� ���>𽊃��.�F���|��"i<@p=6Zk=��=j�=�@�=�GZ=���<��ɻ��Y��V��<�9눾Uܷ����	��!�ҟ1��<��s?��g;��X0� Z�L
� _�𙳾b���6��   �   �+�}���vA��VM;���<��)=6-==2=+=�]�<͂;d6��l���l��X��z���t�ٽ�{�K~��bٽ߽�k ��֮O��м ��98��< �==ԧ�=�u�=V!�=���=�َ=xM=(��<���U���x���r�<�����L���=,���E��gY�pf��&j��se�fX��?D�|�*�lm���f����Bq��   �   FG�h����h�(EX�ܟ�<q=r�2=�,9=�n(=Գ=�c�<�I<����(G��(��Ju$�s@�*L��uE���+����������F:�0�<|�=��f=Sϒ=��=��=}�= Z�=-P�=�;=`t<�$��s׽��?�8"���ξ!��:*�L<K�Ԃh�N��������׆�E�~�5�g�2lJ�Q�)�����ϾR딾�   �   $m����Vǝ��㼀�;���<`�%=v�9=�7=�&=H=H��<�`�<��.<��;�������0R������p]�;�.d<�X�<"�=`�X=�8�=¿�=F͹=��=` �=[z�=,^�=l��=�)= ֶ9�Ac�,��Sb�.|���K�z���A���f�۩�����ݴ��_w������8H��$n���Qf���A�8��\X�a���   �   򕅾�)��U���	!�@�<غ<Dy=�R7=��?=@�:=��,=�=j�	=�l�<$'�<8E�<��<\�<8P�< �=�6=2]=�v�=L�=k~�=�P�=���=���=�6�=N�=��=�0�=��=p��X������#}����������*��T�`|�幏�ң����������9q��A���J���x=|�X�T��+�~j������   �   t7��*8��)ӽLR?�0��l�<B�=h�4=DwC=�E=7?=~]6= �-=t"'=��#=��$=� +=��6=ئH=
�`=�i~=v��=`�=~��=��=R�=���=�6�=(�=��=ğ�=Ȍ=�D=8PH��T����"�J��K�Ⱦɏ
��~4���_��ބ��i��� ��`T��񆲿�N���������� ���`���5�f��Тξ�   �   ��=��Tڽ�I����g�<�o=�]3=(rD=6YH=�E=|�>=K9=F�5=V^5=��8=�;A=�N=0a=$	y=�=���=���=櫿=���=�}�=J��=h@�=���=�D�=�@�=�7�=�z=��d�����^
'��K��(�̾	>���7�t�c�8��a���ߨ�k[������2[��V먿5��������d��a9��h��Ӿ�   �   �6���(8��'ӽlO?� q���<ȣ=΄4=�xC=�E= 8?=�^6=�-=L#'=4�#=6�$=+=N�6=0�H=R�`=
j~=���="`�=���=�=j�=���=�6�=T�=��='��=�Ȍ=BF=�FH�S��v�"�FI��:�Ⱦ�
�~4���_�6ބ�i�������S��*���N��>����� ���`��5������ξ�   �   V����)��Q��$!�@��@ߺ<L|=�U7=��?=~�:=��,=��=4�	=�o�<�)�<�G�<��<��<�Q�<��=R6=l2]=w�=*L�=�~�=�P�=��=��=7�=��=܆�=�1�=��=p��$�̏�� }�����V���*��T�|�����o�������y����o��و������$;|�T�T�^�+�"i�x����   �   �m�<��O�܆��I�;x��<��%=8�9=��7=<�&=4=Ċ�<xe�<x�.<���;����@���I�������b�;�0d<�Y�<~�=��X=�8�=���=�͹=R�=� �={�=3_�=ﶏ=j�)= ��9�8c���b�[y��H�Dx�̫A�u�f����(���ײ��Ou������FF��Wl���Nf��A�����T�t	���   �   �G�g��Ҽh�H X�t��<�v=~�2=019=�r(=��=�j�<�V< ����A���	��ps$�|q@��(L��tE�ʍ+�l���t����%F:�1�<�=��f=�ϒ=��=,�=V�=^[�=�Q�=h�;=��<@�#�gl׽��?������ξO�c7*�8K��~h��}�_���|��Ն���~��g�YhJ���)�(��JϾ�甾�   �   �%���44�`�M;���<b�)=�2==�2=�/=f�<��;h/��8��$l��W��y�����ٽN{��}�~bٽ�޽�( ��T�O��м �9`��<��==L��=mv�=J"�=^��=�ێ=R M=̒�<����Fx������r�U7��˶�½��9,�W�E��bY�$�e�!j�fne�aX��:D�R�*��i��y⾙���;q��   �   � ߽��X���'�%�<:�=�@B=�A=�z!=��<�b�;x줼�F�Ǽ���H�����&)�E'=���H��J���B��V1���P>�L�����F���|��%i<4q=�[k=��=vk�=�B�=�MZ=���<�hɻ2}Y�pK�Ҩ<��戾pַ���辢�!���1�=<��n?�Nb;��S0�mU��	��W�󓳾�
��x�6��   �   ���Ĕ�� 2S<RH=B�G=�T=v�==p=��6<����R�6�����4���_�����YM��:9��q|���ė��p���w�>)M�F��ޯ޽B7��˼�<�&=�aY=�H�=N��= �`=`�=~<<��;�����	��N�䰌�Kų��پS��U�
��,�`��|Y��E	�����)Ծ���������@�r����   �   �ټX�<ZV=�aN=��i=J_=��/=p׷<0�ۻ�A5�ou�� �l;K�ﺃ��נ�G���J�ξX۾ ߾�Tپ;�ʾ�鴾$���f�v���8�������<�ټhl<�P=4^N=��i=�I_=��/=ݷ<P�ۻ`:5�Gp������6K�+����Ԡ������ξ�S۾��޾oPپ��ʾ�崾����F|v�j�8����������   �   �<-=*fY=sJ�=��=�`=��=(p<���o�����	��#N�h���iȳ���پ_W����
�/����\�IH	�R���("Ծ���n��t�@��������p��� S<.D=ơG=�T=�==v!=8�6<옋���Q�j����G�4���_������I��}5���x������4m���
w�8#M����޽$0���h˼�   �   |x=�`k=��=�l�=eC�=:MZ=���<@�ɻX�Y��O���<��舾 ٷ�K�辛�N!�4�1��<�7q?��d;�VV0��W�>�	��[����	��R�6�w߽j�X� �'�$�<`�=�?B=�A=2|!=8�<P��;�ޤ��F�ɶ��yA�]���!)��!=���H���J�b�B��P1�l���4��z��H�F��s|�0Ki<�   �   8��=�x�=�#�=:��=(܎=�M=P��<���a{��C���r�l9��y��i���;,���E�^eY���e��#j�qe��cX�J=D�t�*��k��|����?q��(�(����:� �M;|��<��)=82==�2=|1=�l�<��;L!������k��P��������ٽ�q�1t��Xٽ�ս������O�,�ϼ ��9 ��<:�==�   �   7�=��=v�=\�=R�=��;= �<��#�Io׽��?�O ��w�ξ���8*�K:K���h�������}���ֆ���~��g�UjJ���)�����Ͼ�锾�G�����h�81X����<.u=��2=Z19=t(=�=�q�<0k<`f��$1�������g$��d@�"L��fE��+����j���I:8F�<��=2�f=�Ғ=�   �   ��="�=�{�=�_�=���=��)= �9�;c�@���b��z���I�Fy�
�A��f�먃����ճ��Tv������DG��Em��EPf�Z�A�!���V��� "m�����ĝ��㼐5�;8��<��%=�9=$�7=��&=�	=���<�n�<p�.<P5�; �����~������L�� ��;8Wd<�k�<��=�X=<�=�£=�Ϲ=�   �   "��=�7�=S�=��=2�=l�=���(􊽒���!}����������*��T� |�5������>���5����p����������c<|�k�T�L�+��i�����<���f�)��S���!�@���ܺ<�{=dU7=2�?=P�:=$�,=�=��	=�v�<H2�<HQ�<��<�*�<�]�<��=L"6=8]=�y�=xN�=���=]R�=d��=�   �   p7�=��=T��=P��=�Ȍ=&F=`HH�lS����"�~I����ȾT�
�U~4�.�_�sބ�_i��G ���S������rN�����s���Z ����`���5���d�ξ#7���)8��(ӽ�P?� y黰�<b�=��4=�xC=�E=�8?=V_6=0�-=�$'= �#=N�$=|+=��6=��H=(�`=�l~=ބ�=Ta�=���=��=.�=���=�   �   � >���=`��=���=�-�=8�v=�п<��мIE��6[+�|�����!���V���>��[�~Lq�_��87��3��[q�[O[�|?�cc �� �&�ľ����5D��������M�X��@ܻ;xyY<ܨ�<XÊ<艉<���<�e�<l9�<���<, =�=:�8="�X=��z=���=�;�=R˳=��=�r�=���=j��=Z��=�   �   ���=�=�D�=.+�=�4�=��x=ܘ�<D����z��d)'�����C��ɹ��d[��o;��W���l���z�8����z���l��FW���;�WJ����]���ы�<&?�
"�Y��4l�� �0*�;��n<�ݍ<�<�_�<��<ذ�<\��<��<,�<�}=�T)=f�G=0�h=9��=o�=l�=_�=Z��=���=���=jh�=�   �   p��=(��=�,�=T~�=��=�$~=�k�<ז��מ�N�&hv��$������KK1���K��q`��m�
Ir���m�H`���K�As1�M�M�?����P��=t0�@�۽��n�Ԓü@���x.C<h�<�Ǥ<�>�<G�<HX�<�ju<P�|<���<�<0��<�J�<�`=(�2=~ U=� {=/�=Hڦ=:s�=���=��=���=�   �   ԓ�=l��=�6�=�l�=B�=4��=�=��+�d��w���\�}�Ծ�I�xz!�P�9�i�L�hY�,]���X��nL��E9�{)!�I���վ-�����f��~������7��)X����;d��<T>�<H��<���<`m�<�H\<�| <���;P%�;���;���;P�<�!j<P_�<PI�<`=�L=d}=z�=2Z�=p��=��=�   �   8��=2��=j��=�H�=B^�='�=�_=�A[�l�K���b9<�V]�����O��Bw�K�"���3�5�>�TB�Y>��83�{"���j龆0��[ቾgA������抽��� x�94�<��<��<,O�<��<hV�<��< �:  Ļ�F��+���衼lۦ�\敼�(Z��y����;u�<(�=&�F=T�=T͞=6�=�   �   $	�=nu�=Yf�=�g�=�=���=""-= �<��W���ƕ���b��L��s�ľ�g	�����!��$��y �"��Z�����$��N�F^�J���o��V/�X�0,�<���<��=��=�#=���<X�V< �O:(�G�<Uμ����E�6�h�d�}��u���u��_U��5#���ü�����m<~�=�Y=*=�   �   <q}=^m�=?��=�?�=�e�=,A�=H�==�'�<| ��r�z�g��m2���u������꿾�޾���kU�&��΂�H���پ�U��������h�B(&�3Nս&Ob��}����J<��=�.=�;=�:/=|�=�4�<��; �?��� �tT�D;���/����ؽ����|�����n��~�ɽ�4��v�`������7���<��3=�   �   �=^[e=�n�=	��=�Ɠ=��=<�G=X�<�j'��9�jg��f��k�:���q������l���佾\Vɾ�̾NǾ����)�������_���%�8߽��|��T���D<�H=#A=(]=��[=�a@=2�=D��<�#���$񼮍j�7���Wz����{�,��P?���I�{�J��8B��:0�Dk�q��ը�BEE������[<�   �   @X<Ti=�KR=��z=��=��t=&�H=�=�G<Þ�h�W�S���Y��D�/���W�,<{��8��kg���>���q��P_���j�:�A�&:�|�Ͻ��s� ���w<po=JPR=j�z=�=�t=R�H=�=<<�̞���W�d������d�/���W��A{��;���j��DB��u��qb���j�T�A��>���Ͻ�s��ϴ��   �   �e��p*<�C=A=F
]=��[=�`@=��=��<��`�h�j�����}s����Ĳ,��K?�N�I���J�13B�o50�^f����&Ψ�t8E�@��Ȳ[<��=�`e=�p�=��=�Ǔ=E�=��G=X�<�'��?��k��\��>�:��r�a�p��Z轾Zɾ̍̾�Ǿ���`��z����_���%��>߽��|��   �   �Wb�@���H�J<��=��-=��;=b9/=4�=�6�< -�;Ц?�X� ��T��5��9)����ؽ����s������O����ɽ�,����`�|���!7��,�<.�3=w}=�o�=���=�@�=3f�=EA�=8�==�"�<x)��P{��k�8q2���u�'�����޾����eW�*��Ƅ���h�پ�X������$�h��+&��Sս�   �   t��/��&��#�<��<n�=2�=#=d��<h�V< �P:��G�PHμ�����E�lxh�B�}��n����u�bQU��'#���ü�P��@Gm<.�=&	Y=#ō=��=Pw�=�g�=�h�=p�=���=� -=�<�����K��B�b��N���ľ�Hi	�����!��$��{ ��������꾳��k򖾲^�����   �   �����銽(�� �9���< ��<H��<M�<�<�W�<x�< |�:��û(�F�����֡��Ǧ�4ѕ��Y��"���p�;Ј�< �=�F=�W�=0О=��=��=���=n��=�I�=t^�=��=�]=�\�>L�����;<��^���	��˭꾵x���"���3��>��UB��Z>�h:3�"�{����x2���≾�iA��   �   6������7��6X� ��;���<�:�<���<���<�m�<�M\<�� <���;`H�; )�;`��;��<0@j<o�<Y�<�g=�L=� }=�|�=�\�=���=v�=4��=x��=�7�=�l�=I�=ܭ�=H=��+�Hf���x��\���D�Ծ�J��{!���9���L��Y��-]�T�X�^pL��F9��*!��I�D�վx���� g��   �   ^u0��۽z�n�ėü�䬺�'C<x�<�Ť<�=�<G�<�Y�<�pu<�|<`��<D�<���<�S�<�e=R�2=�%U=�%{=��=oܦ= u�=���=Z�=��=X��=ֈ�=4-�=�~�=��=�#~=�h�<�ۖ��ٞ����iv��%��_�꾲��8L1���K��r`�@�m�.Jr���m�I`��K�t1��M�p�)���AQ���   �   �&?��"����n��� Ỡ!�;(�n<h܍<p�<�_�<̍�<���<؅�<d��< 0�< �=zW)=�G=��h=���=ip�=Zm�=-`�=\��=���=���=i�=��=j�=E�=B+�=�4�=Z�x=��<D����{��(*'�x���%D�������[�vp;�l W���l���z����Z�z�{�l�0GW��;��J�D��ʢ��wы��   �   l5D��������M�0��`ڻ;�xY<���<@Ê< ��<@��<�f�<\:�<л�<� =��=ȭ8=��X=>�z=1��=�;�=�˳=��=s�=��=���=l��=� >���=Z��=~��=�-�=��v=�Ͽ<�м�E��r[+�6|�����S���'V���>��[��Lq�i��:7��0��x[q�NO[�	|?�Uc �� ��ľ����   �   z%?�� ����i�����1�;��n<��<	�<0c�< ��<���<���<���<@2�<�=BX)=��G=p�h=���=�p�=~m�=K`�=r��=���=ĝ�="i�=*��=��=DE�=�+�=J5�=��x=���<8��� z���('�����"C��S���[��o;�jW�r�l�i�z����3�z�`�l�+FW��;��I���������Ћ��   �   �r0�4۽X�n���ü�Z��H7C<��<�̤<|D�<�M�<�_�<X|u<�|<D�<l�<(��<�V�<�f=R�2=r&U=X&{=��=�ܦ=Nu�=˗�=��=��=���=$��=�-�="�=��=j&~=�o�<Җ�K֞�J��fv��#�����=���J1���K��p`��m��Gr�l�m��F`���K�Wr1�8L���#����O���   �   �|����(�7��X���;��<�D�<Ș�<$��<w�<(_\<� <���;`c�;�@�;P��;��<�Fj<�q�< [�<~h=HL=t!}="}�=�\�=ȶ�=��=���=��=N8�=�m�=��=���==��+��a���u���\��ힾ�Ծ�H�Zy!��9��L��Y��*]�F�X�tmL�,D9�<(!��G�Ӹվ����O�f��   �   b����㊽��� ��9l�<8��<���<�X�<p�<�b�<��<��:P�ûvF�����С��¦�P͕���Y����`x�;T��<��=��F=�W�=rО=��=x��=%��='��=�J�=�_�=��=�c=�Z�(�K����6<��[���������u���"�O�3�k�>�<RB�DW>��63��"������`.���߉�BdA��   �   .k���/����6�<D��<��=��=�)=��<��V< �Q:�G�d>μF����E�Duh���}��m���u�PU��&#�8�ü�K���Im<ҽ=�	Y=zō=��=�w�=|h�=�i�=�=��='-=��<����������g�b��J����ľ���e	�����!��$��w �>�����i�j����]�P���   �   �Eb�Hn��0�J<n�=�.=:�;=V@/=܊=�C�<@^�;��?��} ��T��3��\'��T�ؽK���r���������C�ɽ',��<�`�4��`7��-�<��3=�w}=8p�=���=B�=�g�=�C�=��==�4�<�����z�$a�Rj2� �u������翾=޾I���rS�%��Ҁ�y��~�پ�R��=���J�h��$&�-Hս�   �   ,B���b<4O=�(A=r]=&�[=�g@=�=d��<�֌�H�L�j�f���iq�����,�K?���I�q�J��2B�550�*f�\���ͨ��7E���p�[<��=�ae=Uq�=���=qɓ=��=�G=��<��&�0�}a��Ѹ��:���q������i��J὾�Rɾ9�̾�Ǿ�}���
�������
_�F�%��0߽r�|��   �   ��<vv=XVR=��z=��=��t=j�H=�=`^<\���b�W����N��Y�/���W��;{��8��9g���>���q��8_���j��A�:�4�ϽV�s�����Hz<vp=�QR=h�z=��=N�t=*�H=�=�g< ���
�W�����X����/�K�W�C6{��5��d���;��jn��\���j��A��5���Ͻ��s�Ԧ���   �   ��="ge=Ts�=��=^ʓ=��=��G=��<�'�85�?e��l����:�1�q�@����l���佾4Vɾ�̾4Ǿ{����������_�z�%��7߽b�|�XS��PH< J=�$A=�]=d�[=�f@=V�=���< ���T�yj�����:k�����,�,F?���I���J�n-B��/0�Ha����/ƨ��*E�j��[<�   �   �}}=pr�=l��=DC�=�h�=�C�=�==�0�< ����z�He�*m2���u�H����꿾u޾����]U���Ƃ�;����پ�U��걗���h�((&��Mս�Nb�$|����J<l�=�.=&�;="?/=��=�D�<�n�;H�?�|x �dT��.��e!��Z�ؽl��Dj�����Ԁ罻�ɽ7$����`��h�k6��?�<*�3=�   �   B�=�y�=�i�=�j�=��=��=&-=x�<p �������F�b��L��:�ľ��{g	�����!��$��y ���V�������D�.^�2���o���/��x.�<��<r�=r�=�(=��<��V< �R:تG��3μ&y���E��jh���}�Cg��t�u�`BU��#�T�ü��qm<j�=�Y=hȍ=�   �   @��=���=$��=BK�=0`�=��=�b=��Z���K����8<�]�����*��4w�A�"���3�1�>�TB�Y>��83�w"���c�~0��Tቾ�fA������抽8�� ��9��<܍�<p��<�V�<��<�c�<�<�g�:��û�aF�	������`���<�����Y�pǮ��Ǳ; ��<H�=>�F=[�=:Ӟ="��=�   �   ̖�=؜�=�8�==n�=��=o��="=`�+�1c���v���\��]�Ծ�I�oz!�K�9�e�L�gY�,]���X��nL��E9�y)!��H���վ%�����f��~�Y��0�7��&X���;��<8B�<Ė�<즰< w�<�a\<�� < ��;@}�;pb�;`��;��< aj<��<(i�<bo=�L=�'}=��=D_�=���=\�=�   �   d��=���=
.�=j�=��=8&~=�n�<�Ԗ�Oמ���gv��$����޸�EK1���K��q`��m�	Ir���m�H`���K�@s1�M�K�<����P��1t0�"�۽4�n��ü����2C<��<�ʤ<pC�<@M�<D`�<�~u<��|<��<D�<��<�]�<�j=��2=�*U=�*{=��=�ަ=w�=F��=��=��=�   �   ���=��=tE�=�+�=X5�=��x=,��< ���\z��H)'�蔃�uC��¹��a[��o;��W���l���z�:����z���l��FW���;�VJ����Y���ы�8&?��!�C���k����0-�;�n<Tߍ<x�<�b�<��<ص�<4��<��<�3�<�=�Y)=V�G=@�h=� �=�q�=en�=!a�=;��=B��=Z��=�i�=�   �   ��>qA>5" >�E�=��=��=Y= �<���ڰ�����m�j�����о���� ��Ŵ"���,�oe0���,�1�"�|���'�Ӿ�7���/�ې8�߃����>,Y��0��\޼��ѼQ��.����X�$��K��,ᵼ��4�@j;d�<]�<Zn7=�Co=��=T��=f_�=���=���=��=�i>xH>�   �   |\>�&>ܚ�=��=e"�=G��=x�Z=h��< �伺���.0���h������̾�����ȡ���)�7-���)�Р��7�R����]Ͼ'���Q"y���3���������N��J���˼�տ��$ռ�����)�� �(������h=���m:��l<̤�<L�,=Įc=��=ly�=�^�=�H�=^��=Ԅ�=Z��=I�>�   �   �&>W� >(o�=(x�=�=3s�=H1_=H/�<P~��=ڜ��x��1Z�*,�������꾌��	���0 ��h#�� �������뾹�¾�˙���g��y%�:�߽���>�-���Լ�c��<��� Σ��ɼ@�����f�6�<ݴ���Y�`�-�x�<�z�<,�="@=�dr=6��=��=��=�!�=���=���=���=�   �   ���=���=�Q�=p��=v��=d^�= �d=l��<���\t��/C����C��������Ծ�������<}�9\��6�Ve�2���=�Ӿ"���5��;0L�fJ�-�����a�Բ����t��#� >�� �0��P���]����м��߼��ؼ��� ��P�� �йP�<X�<Z�=�a1=�.b=���=��=fa�=h��=�M�=̭�=�   �   @H�=���=V��=���=�(�=�{�= �h=���<����
W��Uֽ8(�l�j�Kؗ�c��!L׾.�����W���������ԾĎ���U����g��i)���[���t�8�f���S�@v�;���;��:P��� �L��z��Ha��0AѼ��Ӽ\�żɨ� 	}��t��!�Z<\L�<��=�f7="�m=P��=�٪=$��=��=�   �   ���=/S�=d�=)�=4ݷ=�Ǜ=jNh=^ = ݹ�������
��B��X}����a3��`�Ǿ�ZԾؾC�Ҿ��ľ:���쟕���q��8�����H2��Uy����;�Gz<���< �<pT<-�;��k�ؙK��Y�� ,޼ K� ��,�������t����Q��p@K� �8��l<`;�<�]<=�J{=�$�=S�=�   �   z�=#ʱ=��=$H�=�}�=(V�=�7a=�#=05�;�y׼6Ⴝ�/ٽ��ϱJ��~x�ht�� (���ȩ��I���T��K\������ g���6�6[�S챽$E�Xc����;L�<��=v�=�h=�)�<hZ|<��;H-�h̨�2_�� 3�V�[�vc}��y��&ޏ�=�������[_��(��Qɼ0ּ�@�e<�:	=�R=��=�   �   4�p=Ê�=�r�=�͞=嶖=���=�(Q=8�=
)<�����"?�E/����>s�̌>��#]�xt����NJ��l>{�>�f��<I��%�=	���}���B��J���(<���<�j-=�7G=�?I=��6=��=h'�<�R<�s껀�ʼ�/�>�z��Q��
���<�۽m��$��s���ܽᲽ��U����K�D�̼ 4n�@�<$S/=�   �   �N= QP=B�v='�=�,=%d=�7=��<5;<�c �����	q� ����你b�z� ��y0���8���8��/���֫���н��"�0*��ew<bU=�VP=��v=0�=�/=�'d=7=T��<�4;<�i � ��q����G���e�;� ��}0�)�8�L�8���/����ݲн^����"�X>*��Fw<�   �   ��(<��<�e-=3G=�;I=b�6=�=�#�<O<�o�X�ʼ�/�0�z�fM��ԝ���۽f�b���z�
ܽU����N����K��p̼ �d���<�Y/=��p=5��=�t�=<Ϟ=N��=���=�)Q=��=H)<���v'?��2��9�Hv�~�>�*(]��|t����L���C{�,�f�RAI��%�K��ރ��
B�l��   �   �q��P��;�׾< �=<�=e=#�< P|<@�;`/��ʨ��\��3��[�\[}��t���؏��������.N_���(�t:ɼ@�����e<�B	=�R=��=�|�=A̱=A�=�I�=�~�=�V�=�8a=|#=@'�;��׼�ソ|3ٽ<�+�J���x��v���*���˩��L���W���^��v����$g���6�X^��񱽴,E��   �   �O2��my��l�;�4z<��<8�<`�S<��;`l�ȞK��Y��P)޼H������ �D��\����=���K� �8 "m<�L�<be<=LQ{=�'�=��=���=�T�=je�=$*�=	޷=ț=�Nh=] = J޹������
���B�G\}�����5���Ǿ�]Ծ�ؾ
�Ҿ*�ľ�������a�q��8��W����   �   �����y���f� U�PU�; |�; �:�˹���L�~���b��@Ѽ؛Ӽ�ż@�����|��Z��2��x<�[�<�=�m7=��m=P=�ܪ=n��=��=�I�=���=n��=R��=D)�=|�=��h=X��<ؚ��W��XֽO(�"�j��ٗ� e��fN׾���R���>Y�F���;��C�Ծ����:W����g�l)�w��   �   ݖ��4�a�������t�82��X����0�tV��hb���м��߼p�ؼ伻������ �ι<��<�=�g1=4b=j��=���=�c�=Z��=|O�=@��=���=���=LR�=���=���=q^�=��d=���<���Fv���E����C�I���c���}�Ծ�������Y~�Y]�8�^f������Ӿ����c��02L�L��   �   ,�߽����V�-���Լ�i��t���ӣ�0�ɼ��ι�Hg�06��۴��Y�`�-���<P��<��=�@=�hr=��=��=��=\#�=��=���=���=F'>�� >�o�=|x�=F�=.s�=�0_=�,�<p����ۜ��y�03Z�-������V��H��Ӻ��1 �Ui#�� �ʌ����	뾽�¾�̙���g��z%��   �   '��������N��L���˼ٿ��'ռx��0���)�� �����P���<��Kn:��l<���<p�,=��c=��=zz�=�_�=xI�=0��=���=���=��>�\>-'>��=��=z"�=:��=�Z=���<��伷����0�h�h�����\�̾�����9��-�)��-�(�)�2���7�����^Ͼ����#y�9�3��   �   ���*���,Y�r1�0^޼��ѼR�8/���fX�μ�J���ߵ���4� x;$�<�^�<&o7=�Do=X��=���=�_�=���=���=��=�i>�H>��>|A>;" >�E�=��=��=�Y=P�<���Vڰ�@����m�������о���2��Ӵ"���,�te0���,�/�"�v����Ӿ�7���/�א8��   �   �������N��I���˼Կ��"ռH�����0'�B��������H�<���n:P�l<��<l�,=��c=�=�z�=`�=�I�=P��=���=��=��>�\>@'>L��=  �=�"�=���=\�Z=d��<�������/���h�İ��F�̾����N�p��Z�)��-�R�)�f��D7������\Ͼ����v!y���3��   �   G�߽�����-�X�Լ�_��ď��Lɣ�,�ɼ���ش�xb�-�pӴ� �Y���-���<̅�<��=`@=�ir=���=��=��=�#�=��=��=���=b'>�� >p�=�x�=��=t�=T3_=�3�<�x���؜�{w�t0Z�_+�����������R���/ ��g#�� �F��,���뾚�¾�ʙ���g�qx%��   �   r���2�a�T���@�t��#��Xw0��H���T��@�м$�߼ԍؼT���L���� �̹�<�<�=:i1=V5b=⢉=䪡=�c�=���=�O�=���=*��=H��=�R�=���=���=�_�=8�d=���<L���q��@���C�샇�����#�Ծ�������*|� [��5�Hd�<���y�Ӿ������� .L��H��   �   ����n�p�f���R�p��;p��;��:���X�L�xm���R���0Ѽ��Ӽ��żp�����|��K� s�H�<�_�<��=�n7=��m=�=�ܪ=���=N��=6J�=h��=��=��=[*�=�}�=�h=T��<pz��W��Qֽ�(���j��֗�a���I׾���$����V����F�쾳�Ծ�����S����g�6g)����   �   �A2��=y� ��;�Zz<0��<%�<hT<p^�;@�k��zK�lH���޼�@�ҽ�>��(��8��̦��p8���K� �8('m<�N�<<f<=R{=(�=	�= ��=hU�=f�=+�=>߷=�ɛ=DSh=�c = �ٹ�����<
���B��T}�P���0����Ǿ'XԾ)ؾo�Ҿ��ľ����������q�L8����륽�   �   TT��R�;x�<�=��=@n=|5�<Hu|<�,�;�
�����^T��3�>�[�vU}�er���֏����G�&L_��(��7ɼ@y��X�e<�C	=��R=��=�|�=�̱=��=tJ�=��=�X�=�=a=@*=�o�;�h׼4܂��)ٽ#�ԭJ�.zx��q��R%��Ʃ��F��R���Y������g���6��W��汽�E��   �    )<|��<:p-=�<G=�DI=^�6=�=�5�<�r<`)�xzʼ$�/��z�*J��
�����۽+d����ay�ܽ����N�� �K�8o̼ �c��<�Z/=��p=���=mu�=О=���=a��=�.Q=�=0))<����?�S)����Xo�l�>�	]��rt�����G��	9{��f�8I�`%�����w��^B�h'��   �   P\=z\P=`�v=��="5=~-d=B
7=���<�U;<�C ���jq�ֳ��5��aa�r� ��x0���8�!�8��/�F���� �н��R"��*�(hw<V=hWP=$�v=��=22=
+d=j7=L��<�T;<�? �����p�������佌^�� ��t0���8���8�{/������٣н<쐽h"��)�p�w<�   �   8�p=���=Kw�=�ў=ĺ�=T��=�/Q=��=�&)<܆��>?�*,����r���>��"]�Owt�F��J��>{���f��<I�m%�����}��jB�@H�P�(<���<�k-=�8G=�AI=x�6=��=�1�<�n<)��wʼ,�/��z��F������/�۽�]����rܽX���>G����K�XY̼ fZ���<Za/=�   �   J�=�α=y�=�K�=��=_Y�=H>a=(*= f�;,n׼iނ��,ٽh�ʰJ��}x�t���'���ȩ��I���T��2\������^ g���6�[�챽�#E�8b���$�;��<܏=�=k=�/�<l|< �;(������R��3�N�[��N}�2n���я�����d,@_�,�(��!ɼ�'���f<tK	=x�R=��=�   �   ���=�V�=Ug�=,�=�߷=Pʛ=�Sh=*c = �ڹ4�b����
��B�X}�-�� 3��/�Ǿ�ZԾ�ؾ-�Ҿx�ľ,���ݟ����q�~8�h��諒XH2��Sy�`��;0Kz<,��<��<�T<�I�;@�k���K��I��޼�>�������"�����H����&����J� 0�8�Im<�^�<vm<=fX{=�*�=b�=�   �   �K�=� �=���=܋�=�*�=�}�=
�h=���<����W�GTֽx(�¡j�ؗ��b���K׾�����W����������Ծ����|U����g��i)�f�*����s��f� �S��}�;���;�
:Н��x�L�(q���T���1Ѽ��ӼL�ż������|��7�����<4m�<J�=pu7=��m=rő=>ߪ=���=��=�   �   0��=��=vS�=&��=��=�_�=�d=(��<h��s��B��T�C�܄��������Ծ�������6}�5\��6�Se�*���6�Ӿ���,��*0L�VJ����@�a������t�H!�`6��x�0� M���X����м�߼��ؼ�������� �˹X*<�#�<4�=�m1=�9b=!��=��=�e�=Y��=4Q�=���=�   �   �'>� >hp�=>y�=�=0t�=63_=�2�<�z��mٜ�)x�p1Z�,�������꾃�����0 ��h#�� �������뾵�¾�˙���g��y%� �߽硎���-��Լ c������`̣�l�ɼ��T���c��.輌Դ�`�Y�`�-���<(��<��=�@=�lr=ꦑ=T�=�=�$�=,��= ��=���=�   �   �\>Y'>x��=$ �=�"�=å�=h�Z=4��<@��W���0�]�h������̾�����š���)�6-���)�Ϡ��7�P����]Ͼ%���L"y���3���������N��J��˼,տ��#ռ���L�� (������L	��`�<���n:X�l<���<��,=��c=��=;{�=�`�=J�=���= ��=x��=>�   �   }�
>��	>#i>���=Q�=���=��=$GD=�o<��Ѽw1����v�=���{��)���>����̾{�ھ�G߾ƅھ��̾�	���K��n^���M��y����UU��L�����p�D�w�ލ������tƽXA���i������ ߽��u���pH���Ƽ �>9�P�<�6=���=��=@��=���=XF�=6 > >+�	>�   �   ��	>s�>Yw>2��=���=P��=j�=�zD=Rx<�fȼhM��k[��(�9�.�v�u��5���СȾ�%־W�ھ[־S�Ⱦ'���Ś���~���H�0
��N�ⵥ�B}���/e�DKl��ׇ��U��翿��Qڽ5�6�����"�ٽ�2��a����E�8�Ƽ k��W�<��0=��}=A�=
��=���=.��=\�=9�>�L>�   �   �>zS>�>:��=d�=�[�=x_�=6yD=�C�<̪��zE��J��^3.���g��������ϼ��xɾ�;!ɾ�E��3�������l�2h9�*&��Iʽ�o��4�_���C�~�J�ʣl�d܏��V���Vƽ(ٽ�Lὣ�ܽ�˽�J��{S��d�?�Pʼ`�%���<N�=��g=e'�=�=��=�\�=���=ع�= (>�   �   4��=\S�=���=vx�=�i�=x�=�+�=iB=X��<�����(l��Խ���bmQ������������ݵ��y�����E��얾ߦ���Q�`�!����ʧ��_h�ƚ(��������5�pf��?�������Ⱥ���Ľe(ý#d��L���:Ҁ��o9���ּ`��G<��<�
A=�r�=ċ�=���=^7�=& �=���=D3�=�   �   �H�=V��=���=���=�J�=r��=/��= {;=���<HK�\�G� ̶�2���5���a�(����̓��P��s��&����ΐ��z���	Y�	�-�Dy������_w�h��xü�����V����߼x#���P�]^��c��1���|����ĝ�(_����o��9� ����l�@�:|�<�8=HC=tw}=(�=�|�=M��=�*�=���=�   �   �=���=|��=�B�=`�=��=~�}=��,=X��<����s%�	T���s�Fa�T�<���\�qeu����6҃�.��gk�x�N�\�+��/���½ �����4��`	�� �9: ֈ�H:������@���.�.�Y�;y�����ԅ�tF���f��4E�0�\kۼ�Fl� ���N<ty�<`�)=t�c=�i�=�-�=��=|��=�   �   �=�_�=�>�=vs�=x.�=�ɋ=�_[=�=0kw<���F��Ɛ��ڻ�����l:���0��B�DM�N�|dE�ӹ3�������[���J%v�P-�� � 8�;�m�<�I�<W�<1H<�T;�B�$����
���2��@Q���d��1n���m�N�d���R�~9���eټ8�i� ���<s<���<R�<=^�w=�@�=�S�=�   �   g�=Ȍ�=~��=�k�=؆�=�c=�i,=X��<h(	<�5��o�f.[�����_Xƽwc�,��T�����Z��9��n��I4ѽ������Q�,�Ҽ�4����< ��<$�=F'=(�=�=���<�#<@pO�L����z�;%�ҵM�B�o�������O���Ȑ�����+s���F��r�p�� �Ľ�<�_=�P=�=�=�   �   (T=rn=��t=,i=�MM=�$=� �<h�W<����	���Z
��J�Rw���x��������ɽ�Խ9�ս��̽)ٸ�m��B�j����x�m�0��;��<��&=T=� n=(�t=1i=�RM=n$=�)�<0�W<@��H���Y
��J��x��4{�� ���C�ɽJ�Խ��ս��̽R߸�p����j�6����m�p�;x��<,�&=�   �   ���<:�=�'=��=f�=���<З#<@�O�������l=%�.�M�ƅo�5��u��}L��gĐ�9���� s���F��h���� �ٸΔ<4g=XP=�@�=�=7��=͡�=!n�=�=�c=.m,=X��<�0	<8�5�^p��0[������[ƽ�g����Y����1^�I=�Eu���:ѽ^�����Q��Ҽ��4���<�   �   ��;�a�<�=�<TK�<�H<��;�Y������
���2�nCQ�L�d��1n��m���d�r�R��9�d��Uټ�i� Ӧ��]s<��<@�<=��w=�C�=V�=N�=�a�=x@�=Mu�=00�=Sˋ=�b[=
�=�ow<����:���ݻ������<��0�^�B��M��N�4hE�d�3��������Ĺ��.v�x5��� ��   �   ���@9�� ;8: ���R������L����.�v�Y��?y����օ�<G�8�f��2E�`,�|aۼP/l� I��8�N<,��<�)=��c=�l�=@0�=��=���=��=Z��=��=[D�=la�=���=f�}=4�,=���<P��,v%� V���v�Wc���<���\��hu�� ��ԃ���kk�ͣN�[�+�"2�4�½������   �   D��(�üh����a��ܦ߼<)��Q�&a���e��}���P���Ɲ��_����o�F9�������l�@��:\��<,>=fMC=�|}=��=�=Y��=�,�=^��=<J�=���=��=���=�K�=C��=ƿ�=�{;=��< NK�:�G�>ζ�����5��a�����qΓ��R��=��鿛�SА�R|���Y�z�-�^{�J���Dfw��   �   �dh���(�^��؉���5��f�4B��(����ʺ��Ľ*ýQe��쏟�OҀ�o9���ּp�߻�*G<4��<tA=�t�=���=���=9�=�!�=��=�4�=H��=ZT�=���=By�=�j�=�=�+�=iB=��<P���h+l�Խ<��5oQ� ��澘�����Wߵ�;{��
������햾
����Q�"�!����=ͧ��   �   �q����_�>�C�N�J���l�\ޏ��X��rXƽ�)ٽ'N���ܽ��˽GK��yS����?�`ʼ��%����<��=v�g=�(�=x��=e��=^�=���=κ�=�(>I>�S>=�> �=�d�=�[�=�_�=yD=HB�<̭���F����콂4.�S�g���������м��yɾ'�;:ɾ�F��#���䏐���l�xi9�I'��Kʽ�   �   ���h~��2e��Ml�ه��V��.����Rڽ;	�7����g�ٽ�2���`����E���Ƽ ��d[�<��0=��}=�=ܟ�=���=���=�=��>�L>ѽ	>��>�w>v��=���=s��=j�=pzD=�Ox<�hȼ1N���\��ޕ9��v����Ĕ��i�Ⱦ�&־��ھ�־�Ⱦ���+ƚ�X�~�^�H��
��O��   �   �U������p�p�D�w��ލ�7���uƽ�A�?��d���i��? ߽�������2H��Ƽ @9�R�<�6=$��=��=���=���=�F�=,6 >8><�	>��
>��	>,i>���=Q�=���=��=�FD=��o<��Ѽ�1������=���{��)���>����̾��ھ�G߾ͅھ��̾�	���K��n^���M��y�����   �   K����|��/e��Jl�zׇ�(U��Z����Pڽ=�5��&���ٽ$1��F_��
�E�8�Ƽ ��T^�<��0=��}=w�=$��=���=��=$�=��>M>۽	>��>�w>���=��=���=�j�=�{D=�Vx<�cȼ�L���Z����9���v���ɓ��W�Ⱦt%־��ھ�־ǡȾ���DŚ�ř~��H��	��M��   �   �n����_�r�C�l�J���l�ۏ�gU���Tƽ&ٽUJ��ܽ1�˽H���P���{?�ʼ��%�8��<,�=.�g=s)�=���=���=\^�=ή�= ��=�(>d>�S>`�>$��=e�=�\�=�`�=�{D=8I�<�����C��8��(2.�z�g�E�������μ��wɾ�;
ɾ�D��9���/�����l��f9�%�Hʽ�   �   �[h�2�(�H������5�nf�\=������ź���Ľ�$ýp`��v���T΀�0h9�l�ּp�߻0:G<@��<�A=�u�=f��=��=t9�="�=P��=�4�=���=�T�=��=�y�=\k�=��=1-�=�lB=���<����$#l��Խ���JkQ����O������[ܵ�.x�����
��)떾�����Q���!����ȧ��   �   6���nüȃ���M��T�߼R��P�[��v_��0���.���:���sZ��H�o�9�t����l�@1�:��<A=�OC=N~}=;�=��=���=�,�=���=�J�=��=���=h��=�L�=l®=^��= �;=���<X/K�VyG��Ƕ���6�5���a�����˓�O�����U����̐�,y�� Y���-�w�
����Yw��   �   ���P߃���::�3���$�����<3����.���Y��1y������υ��;���f��)E��$�0Uۼhl��ˠ�x�N<؋�<ԋ)=�c=2m�=�0�=5�=���=V�=���=���=E�=Wb�=>��=��}=�,=��<�p�jk%�[O��Rn�P^��<�1�\��au����6Ѓ�@��ck��N�B�+��,��½#������   �   �i�;�x�<dT�<�a�< HH< �;@&�${��.y
���2�6Q���d��%n���m��yd���R��9�d��4Mټ`�i� ���(es<���<j�<=��w=,D�=tV�=��=Sb�=�@�=�u�=1�=�̋=f[=��=��w<����v��Bջ������6�F�0�$�B�;M��N��`E��3�*��ȱ��͹���v�&%�v ��   �   X��<��=�#'=��=��=���<��#<@�N�0����f�0%��M��zo�C���,���H��s���ֱ��s���F�`f�@ �� 8׸XД<h=	P=A�=k�=���=S��=�n�=ۉ�=��c=�p,=���<�I	<xz5��e��#[������Qƽ�\��������V��5�Hg���-ѽ����
�Q��rҼ��3��	�<�   �   �T=J&n=p�t=p6i=FXM=�$=�7�<X<�	�|�O
���I�Ir��8t��������ɽx�Խ�ս��̽�׸�m����j������m����;���<T�&=�T=�!n=$�t=J2i=:TM=�$=�/�<P�W<@=�t���lP
���I�q��{r��򆷽��ɽ��Խ��սq�̽Ҹ������j�����m� ��;���<,�&=�   �   ��=���=>��=�p�=���=��c=�s,=`��<�R	<�t5��e��$[�'���Tƽ`����4����Z�@9��m���3ѽ�����Q���Ҽ�4���<d��<��='=2�=V�=���<��#< 4O�`����m�23%�r�M��zo�X���Z��0F������ĭ��s��F��\�@ \Ƹ�ߔ<�n=P=�C�=�   �   ���=d�=�B�=�w�=�2�=�͋=�h[=��=8�w<0��Ε�؈�T׻�����9�ԓ0�"�B��M�pN�
dE�~�3�e�����������$v��,��� ��<�;�n�<K�<�X�<�5H<�n;�9�䄵��}
�F�2��9Q�.�d�D'n�T�m��wd�j�R���8�V��h?ټ��i� ᡹X�s<|��<��<=F�w=�F�=�X�=�   �   � �=,��=��=BF�=zc�=J��=��}=J�,=��<(r��l%��P���p�`�D�<���\��du�����у���Bgk�E�N�0�+�Z/�`�½���.��T��`�� �9:�����6����=����.���Y��6y���mх� >���f�H)E� #�Oۼ�
l�@.��0�N<4��<r�)=z�c=�o�=�2�=7
�=���=�   �   �K�=(��=���=R��=\M�=,î=���=��;=쟜<X2K�4{G��ɶ����5���a�օ���̓��P��M������ΐ��z���	Y���-�*y�r���p_w�
��<wü�����U��$�߼�"���P�t]���a������`�����[��"�o��9�4s����l����:�<�D=�SC=\�}==�=��=x��=�.�=��=�   �   l��=lU�=���=fz�=�k�=|�=�-�=$mB=h��<$����$l�HԽ	���lQ����d���]����ݵ��y��w��6��r얾Ԧ���Q�L�!����aʧ��_h�z�(�Z������5��f�-?������Ǻ�ԑĽ�&ýAb������xπ��i9�L�ּ �߻�>G<��<A=�v�=ď�=c��=�:�=6#�=d��=�5�=�   �   �>)T>��>���=`e�=�\�=�`�=�{D=I�<̥��MD��8���2.�|�g��������ϼ��xɾ��;ɾ�E��,���	�����l�&h9�&��Iʽ�o���_�P�C�B�J�l�l�*܏��V��(Vƽ�'ٽ�Kὰ�ܽ��˽iI���Q��>}?�ʼ��%����<��=F�g=*�=���=���=_�=���=���=�(>�   �   ��	>ė>�w>���=D��=���=�j�=�{D=8Wx<4dȼ�L���Z���9���v�a��$���ġȾ�%־P�ھW־P�Ⱦ#���Ś���~���H�'
��N�ٵ��6}���/e�$Kl��ׇ�tU��ƿ��vQڽ��d6�����ٽ2��(`����E���Ƽ /�<]�<��0=��}=��=R��=���=H��=`�=��>!M>�   �   �>�]>��>�1>ސ�=�9�=��=�q�=��9=�m�<�iu��P�Μ��Gv��+��N��2j�R�{�􀾪�{���j�=Q��u2�a��齥8������Ӑ�����
�����5��1� �O���h�U�y�8���y�Lh�D�L�~'*�\$�-p��fEM���j�B�<>�:=�ߍ= ��=�Z�= ��=�1>�>\>�   �   �p>v7
>�s>���=D�=4��=���=s��=�.7=��<�bo�^�L��������J3(��OJ�e8e��ev�T*|��v��Ee��	L�h�-��!�F�oc���7���������R9��=R�����N,�{eJ��sc�*t�}-z��ot�6[c��H�L�&�p� �߱�H2I��7e�t��<�q8=��=�ȳ=L��=�"�=t��=q>n5
>�   �   ��>��>J�>��=T��=���="Ҭ=��=�\/=�:�<�{a�xFA�ک�K���J1��=���V��f��k��ue��(U��<���I��̽~������q�J ���`���`ʽ� �E���c;�,mS�P�c���i���d��&U��]<���g0�䧽4>��JX�|�<�p0=WV�=��=���="��=&z�=��>w�>�   �   L�>�� >^I�=���=t��=�Ϳ=�=lww=h" =Pn<`�W���2��X��vU޽�!�z:+��
A�9{N�5*R���K�`,<�"{%���
�)ݽ ����C���%K�|e8�VJ�Ru~����'۽\D	�0
$���:��J�rP���L��s?�t�)����5ܽ����V�/��$P�h1s<(� =8�w=��=�ÿ=l��=ش�=l4�=�� >�   �    l�=|��=JG�=tD�="��=��=ʎ=�W=�\=hw-<@�d��%�ˋ�!�Ľq��2���:&�^�0��|2�<�+�������޽� ��{���0��| ��-߼����.�THx��,��Rhܽ���a��*���0�"/�O�$� G��M����½5i����#�Hv_�X�0<��=j'W=���=)��=��=��=@%�=<��=�   �   W�=�V�=K�=�j�=�=��=(�j= (=P��<@j`;,���"�@'~�O<����ս�3���m	���^��H�P��mͽLd��D�h����蕪�X�+��G�0a(�$P���u�d�e��u��k6˽�W�J��Bl�F��0L��3���CԽ�媽,|�� �lE��@9d;�6�<��'=$)j=ϔ�=O˫=�$�=n�=@<�=�   �   ���=14�=�0�=c��=vT�=�`b=�C'=p��< <h��tJμ�S-���q��&������|N̽۽��߽�ٽȽ�r��=:���C�P�鼸G6� 4; �?<�$s<�sB<`NJ;�.������@��b���t��WƽΓ׽z�ݽJٽ^�ʽ(p���H����p���,��Vμg��<���<�4&=�Sa=[ڊ=^��=��=��=�   �   rU�=��=�'�=.	v=ցF=^�=�ͣ<�C�;Hc(��qɼ�<�P�L�x�x�~����y���ʦ��é�N��|����&��^�P���X����K���j<���<L�
=d�=|d=03�<8fq< �|��ŋ��-�j�M�͏���8��0棽>����ե��Μ������x�&:M�d���˼HS.�0i�;�<�,=p/E=p�t=�ʌ=vT�=�   �   ��j=X�a=�G=�=��<��,<��0p����D�>�(Rf�_���Y<������:#��r����e��h��A����X��������$<h��<��=��F=�za=t�j=P�a=:�G=H="�<@�,< ���8a�������>��Lf�����e;������*$��J���Ph��z"h��A�D���黻`�$<ę�<4�=��F=�ta=�   �   $�=�]=|%�<�Hq< D���֋�R6��M�񓂽P<��k飽����Mץ�EϜ�Q���ʖx�b6M�V���˼H9.�О�;8��<03=x5E=&u=>͌=W�=X�=ņ�=�*�=v=�F=��=�ڣ< u�;�L(��gɼ9�$�L�
�x�9����{��.ͦ��Ʃ��Q���Ř��*��(�P�6'�`�� �M�|j<���<�
=�   �   �
s<�XB<��I;�%.�P�伴�@��g���y���ƽ�׽3�ݽMٽ��ʽeq��I����p��,�`OμHT�x<���<|:&=PYa=�܊=ԙ�=\�= �=0��=�6�=�2�=���=�V�=fb=�H'=��<0)<؋��Eμ�R-���q�!(��7����Q̽�
۽�߽��ٽ�Ƚ>w���>����C����Pd6� �3;�?<�   �   p{�0|(�t^��n}���e�9z��/;˽�\���yn�@���M�B6��xEԽt檽�+|�V� �$@���qd;?�<�'=�-j=��=lͫ=�&�=b�= >�=�X�=�X�=M�=�l�=�=��=�j=�(=<��<@�`;(���p"�,)~�>��R�ս 7���o	���³�����rͽ~h����h����$����+��   �   �9߼�&��`�.��Ox��0���lܽV��Fd��!*���0�$/���$�VH�uO����½Xi����#��n_���0<�=�*W=|��=﷬=���=B�=�&�=���=�m�=���=�H�=�E�=���=�=�ˎ="W=�^= |-<��d�F�%�H̋�$�Ľ�s�����<&���0�(2���+�8��:��ʦ޽K���{�Ġ0�Ă ��   �   �j8��!J�D{~�����۽BF	�1$���:��J��sP�n�L�u?�t�)����q6ܽ㢙���/� P��9s<�� =��w=��=ſ=���=��=�5�=6� >��>� >�J�=��=���=�ο=
�= yw=�# =�n<8�W��2��Y��eW޽�"� <+��A� }N�.,R���K�F.<��|%���
�1ݽŏ��BF�� +K��   �   �#q�}"�� c��bcʽN� �ğ�xe;��nS�ʟc��i���d��'U�v^<�p���0�䧽D3>��EX���<rr0=[W�=	��=���=��={�=��>�>�>]�>��>Ѕ�=��=���=�Ҭ=�=`]/=�:�<H~a��GA�A۩�ۘ��F2�1�=���V���f�b�k�qwe�$*U�Y�<�R��e��̽�������   �   u�������:��T�����O,�{fJ�ptc��*t�2.z�kpt��[c�I�H�O�&�P� ��ޱ�1I��1e����<�s8=u�=�ɳ=���=*#�=��=\q>�5
>�p>�7
>t>��=��=���=��=���=�.7=��<8eo�r�L�}������3(�XPJ�.9e��fv�)+|��v��Fe�R
L��-�N"�{⽩d���8���   �   KԐ������
�����=6��1�\�O���h�v�y�7����y��Kh���L�'*��#�Eo���CM���j��D�<��:=S��=���=�Z�=L��=�1>�>3\>�>�]>ˣ>�1>��=�9�=��=�q�=r�9=m�<Pku���P� ���vv�8�+��N��2j�u�{�(􀾺�{���j�=Q��u2�:a� ���8�������   �   ޞ��o���29��R�����N,�"eJ� sc�l)t��,z��nt�*Zc���H�*�&�V� ��ܱ�\.I��)e��Ï<�t8=��=ʳ=D��=`#�=4��=qq>�5
>�p>�7
>*t>@��=��=���=Z��=��=�/7=T�<�\o���L��������2(�OJ��7e�ev��)|�v�&Ee��L�ٷ-�2!����b��@7���   �   �q�Z���_���_ʽ8� �p���b;��kS��c�2�i���d��$U��[<�=���,��৽*.>�H5X�䅉<�t0=PX�=���=8��=x��=V{�= �>��>,�>y�>��>��=l��=%��=bӬ=��=�_/=�@�<�ma��BA�ة����0���=�H�V���f�s�k��te�\'U���<����K��S	̽�|��㭂��   �   b8�J��q~������ ۽
C	��$�Ò:��J��oP�~�L�Uq?��)����:1ܽ������/�pP�8Ks<�� =v�w=���=�ſ=D��=���=�5�=[� >��><� >�J�=|��=��=FϿ=��=�{w=�& =�"n<��W��2��U��!R޽���8+��A�&yN�(R�۾K�m*<�Vy%�`�
�Q	ݽ�����A��2"K��   �   %߼\����.�>Cx�*���dܽ���_�.*���0�U/�t�$�FD�EH��p�½'d��z�#��S_��0<<�=�-W=���=θ�=4��=��=8'�=��=�m�=T��=2I�=rF�=Q��=��=�̎=%W=�b=P�-<��d���%�ǋ��Ľ�l��ʁ�(8&�Η0�Vz2���+���������޽@����	{�R�0�x ��   �   �M(�lE���o���e��q��2˽�R���Qi�6��I�-���=Խ�ߪ�� |�$� �T1��`�d;H�<r�'=80j=���=*Ϋ=d'�=��=�>�=HY�=�X�=tM�=,m�=��=��=��j=
	(= ��< �`;`���8"��~�S7��v�ս*.���j	��������#���hͽ�_����h����􉪼��+��   �   h:s<��B<��J;x�-�Tw伔�@�H^���o���ƽ��׽�ݽ}Cٽ��ʽ�i��GB��R�p���,��@μ�<��.<���<=&=B[a=�݊=m��=��=��=���=�6�=Y3�=Z��=�W�=�gb=rK'=���< ;<Ht�7μzI-� �q�O!��P����H̽"۽��߽(�ٽpȽ)m��M5��6�C�P�鼈+6� f4;�?<�   �   ��=�i=�>�<�q< �u������$�"�M�)���s2���ߣ������Υ��ǜ�ߘ���x�~-M�2�d�˼�'.�`��;T��<5=�6E=>u=�͌={W�=lX�=&��='+�=�v=:�F=v�=Tߣ<���;h;(��\ɼ�1�8�L��x�����t���Ħ�����H������!����P�*���  J���j<|��<�
=�   �   ��j=��a=�G=f=�/�<H-< q���M��4��X�>��@f�����4������`�������a���h�z A����L��@���h�$<��<��=��F=B{a= �j=�a=�G=,=t$�<��,<����`[������>�~Ff����s6������U�������_���h���@��������c����$<��<0�=��F=�a=�   �   {Z�=4��=P-�=�v=8�F=ʽ=��<���;%(�hRɼ�-��L�F�x������t��eƦ�#���5K��F����$����P���L����K�p�j<���<��
=�= e=�4�<Xiq< �{�,Ë��+��M�#���T6��f㣽����dѥ�vɜ�����x��+M�����˼�.�p�;H��<r:=
<E=u=�ό=�Y�=�   �   U��=�8�=65�=U �=�Y�=Xlb=P'= ��<hL<e� 1μ�G-���q��!��ě���J̽/۽m�߽3�ٽ�Ƚxq��l9����C�P��xD6� 4;h�?<�&s<vB<�WJ;�.���伦�@�,b���s���ƽ��׽-�ݽ+Gٽ��ʽ�k���C����p���,�=μ�1�=<���<`A&=�_a=�ߊ=k��=��=R�=�   �   �Z�=jZ�=�N�=�n�=o!�=~�= �j=�(=l��<�a;䧏��"�x~�j8��_�ս�0���l	������������lͽ�c����h���������+�@Dເ_(�O��u���e�Bu���5˽�V�����k�`��K��0��}@Խ�᪽<#|�$� ��0��@�d;dL�<4�'=J3j=���=�ϫ=�(�=\�=�?�=�   �   o�=n��=XJ�=�G�=���=8�=�͎=�'W=�d=��-<P�d���%��ǋ�4�Ľ�n��"���9&���0�^|2�֜+���������޽k ���{�2�0�r| �,-߼H��2�.��Gx��,��hܽٓ��a�@*��0�p!/�r�$�F�EK����½�e��j�#��V_�8�0<J�=�/W=���=깬=d��=��=X(�=.��=�   �   `�>�� >�K�=V��=���=0п=��=D}w=N( =�&n<H�W�l�2�4V��`S޽� ��9+�P
A��zN��)R���K�.,<��z%���
��ݽҌ��}C���%K�4e8�J�u~�����۽>D	�

$�Z�:�vJ��qP�Z�L�s?���)�5���3ܽW����/�0P�(Is<*� =0�w=|��=wƿ=��=D��=�6�=�� >�   �   d�>��>�>���=���=���=�Ӭ=��=�`/=B�<`ma�CA��ة������0���=�N�V�Ҥf���k��ue��(U���<���7���
̽�}�������q�5 ���`���`ʽҲ �0���c;�mS�$�c���i�P�d�`&U�V]<�t��/�⧽�0>�@<X�ă�<zt0=KX�=���=~��=Й�=�{�=N�>,�>�   �   �p>�7
>Dt>t��=�=��=���=f��=~07=8�<�[o���L�����4��3(�jOJ�68e��ev�:*|��v��Ee��	L�\�-��!�7�ec���7���������C9��0R�����N,�peJ�rsc�*t�b-z��ot�[c�ݙH��&�� �Lޱ��0I�h0e�4��<�s8=��=�ɳ=,��=d#�=>��=zq>�5
>�   �   ��>`
>��>2� >b��=���= ��=��=��=� 7=��< �/��˼�/K��镽�\��w��e���f���T��������Ƚ�g��!"��Nsy�*>q�i8���t���c�8h��qL����{C��Zݶ�g�˾y)پ��ݾ�+پAm˾�
��\����y�|�;��0 �Mڒ�0�ɼh�}<�dG=
t�=�O�=N��=��=�>,X
>�   �   q
>e	>8>\�=���=v��=e��=D��=f�~=�1=4C�< �G��:˼h�H�G��ml��moܽ�|����0�ｻ�ܽ������n����m�6�e�4.��Ԥ���޽~���8G���|�
������]Ǿ��Ծgپ4�Ծ�ZǾ2f��������t���7�����X��̓�����<r�G=6ә=B0�=�2�=D*�=$$>�G	>�   �   �>��>p� >��=��=]�=��=��=��h=XR=�՘<��7�4μ�AB����[���ͽoF߽����۽��ȽSC��rk����n���K�d�C��'_������Ƚ
�68�7%k�D�����������Ǿj̾�2Ⱦ����}姾����0f�8�,�aM�j!��\����<BTG=!��=��=L��=2��=�2> >�   �   yq >Z��= U�=���=��=�и=��=SV�=\PB=�<HG<0#��
ڼ�;��T���_���o��9XŽ��ƽ��ޔ�����:�h�¸7�~�������'���f��V��E���] ��|O��v�j㕾}짾�س��H������Fw��º��F8����O� ���ѽ�Xh�����.�<�D=W\�=��=R��=��=��= P >�   �   ���=�<�=���=�B�=X�=�:�=z�=\E=^�=�<@��:��m�d���@�:��Yr��ۏ��y���\�����m9�������S�>o�x�⼌椼(k��<�����t�𠸽RB��j,�`YW����ʏ������NI��Ւ�����m`��4�����ⴽNND��x@��F�<��==���=���=�P�=��=,�=��=�   �   Db�=,O�=\x�=���=p�=z�f=�E,=l�<X�V< �^�0Ch��ڼ
��p6F�؝h�l����#��}v��j9|���\��|1���������� ����O:��u��+��L���|��S��X��G;*���L�>�i��B}�^肾�=��4�s�J[���;��H�?���ӗ�j�"��[�,�<�!.=�p=���=�:�=t3�=ؿ�=$	�=�   �   <(�=���=޻�=��z=�@=ܓ = �< ,�9�+_� �Լ�O���7��kR���d��n��o�Ʃf�BS�^�4�Ν�,f���%����:X�E<�P�<ؒ�<(�<�y�;@��<��^�q��S�����E�102�w�C��L��K�@�A��i/��:�cH������w}���
����h�{<:�=�e\=�Z�=�֣=x:�=�)�=�q�=�   �   �-�=ė�=DS=n�=�ܛ< �N:쭌���	�lYC�^(p��s���ʏ�"������� ��o�~~N��P&�<�������a�� <�x�<b�=�=t(=b=d��<8k�<����T�ʼ@qM��*���ν���������m��p��n�����m;Ž����Z���H�3��
<Xn�<��,=�7d=���=��=�f�=���=�   �   >JV=Fu)=p�<P�;�^�d���if�8񘽋Ķ�K�ʽ�,Խdӽ5�Ƚ�����䞽�'����I���
�X������XXV<���<�$=(�M=��i=^v=��o=�PV=r|)=��<PP�;x�]�\��^f�,똽������ʽ�'Խ�ӽ��Ƚw���_㞽2'��V�I�̂
�8Ó�`��hEV<���<n$=��M=��i=�v=��o=�   �   p��<�[�< ���|�ʼ||M��0����νj���B��9 �r���������콊=Ž&��Z�ԫ�`�3�(�
<8v�<�,=<d=���=7�=qi�=;��=�0�=�=hS=\�=�<��P:������	�lOC��p��o��vǏ�����ṍ�?��o�r�N�$T&�� ��%���.b�h�<dm�<��=�=�(=y=�   �   �?�;�����r��Y��(	���H��32�0�C���L�:�K�&�A��k/�c<��J�������x}���
��h�{<`�=|i\=i\�=�أ=�<�=�+�=�s�=�*�=B��=㾖=j�z=@=�� =��< K�9�_�\�Լ$I���7�*hR���d�ʑn���o���f�PFS�n�4�b���q����%� ��:��E<E�<l��<��<�   �   L:�����v�|�`Y��e���>*�{�L��i��F}�3ꂾ�?��)�s�wL[��;�GJ���⽴ԗ���"��W�܂�<$.=�s=���=]<�="5�=���= �=Nd�=pQ�=�z�=���=]�=��f=L,=�x�<��V< D]��0h�$�ڼ���5F�ڞh�����[%���x���>|���\���1�8������H�������
N: `v��   �   �����t�v����D��m,��\W�v��̏�ѱ������J��v֒������n`�4�4�����㴽�ND��u@��I�<��==���=���= R�=h��=��=V�=H��=l>�=��=�D�=��=K=�=T�=�`E=��=��<@C�:��m�������:�P[r�ݏ��{��G_������A<�����T�S��t���⼤񤼜v�������   �   ��f�]Z��O��?` �jO��y��䕾�ڳ�J��Դ��lx������ 9����O������ѽ�Xh�����0�<��D=H]�=��=P��=���=�=�P >r >���=zV�=6��=���=>Ҹ=Ф�=�W�=^SB= �<�G<滜
ڼ�;��U��Fa���q��eZŽ �ƽS�`�������"�h���7�D�����V�'��   �   z�����Ƚ�
�8�Q'k�g���O��������Ǿ!k̾�3Ⱦ����槾X����0f���,��M�4!��4Z�����<�UG=곗=̢�=��=���=�2>x >s�>q�>� >��= ��=~�=��=��=j�h=�S=�ט<��7��μ�BB�����\����ͽ"H߽���ސ۽|�Ƚ1E��Nm��t�n���K�^�C�,_��   �   �դ���޽���:G�^�|�������~^ǾK�Ծ�gپ��Ծ�ZǾcf��������t���7�2������������<�G=�ә=�0�=3�=�*�=g$>H	>Dq
>�	>S8>�\�=D��=��=�=���=2�~="1=�C�< H��;˼H�H��G��=m��`pܽ�}����N��ݬܽ����������m��e��/���   �   �u���d��h�RrL�����C���ݶ���˾�)پ��ݾ�+پm˾�
��
���y���;��/ �(ْ�$�ɼP�}<NfG=�t�=kP�=���=f��=�>MX
>ǥ>4`
>��>F� >|��=���=(��=��=��=� 7=��< 20� ˼*0K�ꕽ�\����Ὠ�������������'�Ƚ�g���"��Bty�d?q�/9���   �    Ԥ��޽����8G���|�������h]Ǿ'�Ծ�fپ��Ծ�YǾje������~�t�|�7�;���%�� ������<B�G=eԙ=G1�=`3�=+�=}$>H	>Rq
>�	>_8>�\�=f��=4��=)��=��=�~=H1=�F�<��G�D7˼��H�=F���k���nܽ�{����L���ܽG���� �������m��e�,.���   �   5�����Ƚ�
��8�Y$k�����i��������Ǿ�h̾�1Ⱦ����?䧾�����-f�,�,��I�:��Q�����<PXG=ഗ=���=���=`��=3>� >��>��>� >��=@��=��=���=|�=�h=�U=4ݘ<`�7���ͼ�=B����Y���ͽ\D߽���۽��Ƚ�A���i��>�n���K���C�&_��   �   ��f�.U��K�뽼\ �R{O��t�R╾4맾�׳�G��߱���u��!����6���O�i��y�ѽ�Ph� ���:�<P�D=�^�=��=��=|��=��=�P >7r >��=�V�=~��=��=�Ҹ=r��=�X�=�UB= �<�#G<����ټ�;��Q���\���l��,UŽ��ƽ��;���������h��7��������'��   �   ���(�t�7����@�i,�WW�>�Hɏ�H���: ��^G��"Ӓ�����~i`���4����^ݴ��DD�xW@�XU�<�==�Ë= ¯=�R�=
��=�=��=���=�>�=>��="E�=�=�=�=��=�bE=~�=�&�<@��:�m��v��d�:��Qr��׏��u��Y��N����5��x����S��i���⼤ݤ��b��X����   �   �!������||�/P�����8*���L���i� ?}�U悾�;�� �s��E[��;�ME�����͗���"�h6����<�(.=Tw=� =R=�=�5�=(��=l�=�d�=�Q�=0{�=��=��=�f=�M,=\}�<�W<�L\�0h�آڼ~z��,F�p�h�̶�����r�� 1|��\��u1�|���L��h��@_�� �P:��u��   �   ���;�y�h��Z�q�O�������A��,2���C�ɆL���K���A�\e/��6��@��1��&k}���
�P]�p�{<B�=m\=�]�=�٣=:=�=D,�=0t�=+�=���==��=2�z=@=� =4�< j�9��^���Լ4D�h�7��`R���d�X�n��vo���f��8S�f�4�V��|V��`�%�@[�: �E<�[�<��<\�<�   �   8��<(w�< ���X�ʼ�gM�%��ԥν��������P��O��Z�����4Ž*�����Y�j���w3�X�
<��<��,=�>d=���=��=�i�=���=1�=H��=S=�=��< @Q:������	��LC�>p�`m��ď�♑�����E鄽��o�6tN�G&�����
���[a�H) <���<F�="=�(=��=�   �   �UV=>�)=�!�< ��;(�]�,��vRf��䘽����(�ʽ Խ3ӽ�Ƚ����6ܞ�n ����I�w
�|���`/��iV<(��<�$=�M=:j=Xv=R�o=RQV=})=��<�U�;0�]�X���\f�@꘽I�����ʽ�%ԽNӽv�Ƚ�����ޞ�"��2�I��v
����� �vV<D��<�"$=ʽM=*j=Zv=��o=�   �   3�=���=hS=:�=���<�=S:D���D�	��BC��p��h��p���x���貍��焽��o�,tN��H&�H�Ｔ����a�( <�|�<�=�=R(=�=���<Pl�<@���,�ʼ�pM�*��v�ν����O��=����N����A�콄7Ž������Y���� w3���
<؃�<@�,=�Ad=v��=�	�=�k�=���=�   �   �,�=���=���=|�z=@=�� =��< E�9p�^�L�Լ =�H�7��[R�2�d�x�n��vo�*�f�6;S���4�����_��x�%�@��:��E<�R�<T��<\�<�}�;H��³���q�tS��.���D��/2��C�`�L�8�K�V�A�dh/�'9�"E��`���po}�:�
�@a�0�{<d�=�n\=�^�=�ڣ=�>�=�-�=�u�=�   �   f�=`S�=}�=,��=A�=J�f=�S,=X��<�#W<��Z�Ph��ڼ4w��*F��h�;��� ���s��5|���\�pz1�T������x���镺��O: �u��*�������|��S��:��';*���L��i��B}�*肾�=��~�s�I[��;��G�U�⽝З�z�"�P>���<).=8x=�à=:>�=�6�=P��=��=�   �   ���=�?�=���=�F�=��=�?�=<�=HgE=��=@/�< I�:P�m��r����:�Rr�e؏�Dw���Z��a���,8�����0�S�Hn����T夼,j���������x�t�Š��@B��j,�HYW����ʏ�믚����I���Ԓ�.���Hl`��4����Aഽ ID�b@�hR�<x�==�Ë=W¯=�S�=���=��=��=�   �   �r >Ě�=�W�=���=4��=*Ը= ��=oZ�=�XB=��<�-G<��廴�ټ��;�R���]��n���VŽy�ƽ�］>���������h�.�7���d����'�J�f��V��)���] ��|O��v�^㕾o짾�س��H��_���w�������7��@�O�9��O�ѽ�Th�����6�<F�D=n^�=��=T��=��=�=+Q >�   �   ��>��>S� >��=��=��=~��=z�=�h=�W=h��<@�7��ͼ�=B�J��>Z����ͽ�E߽Y��k�۽0�Ƚ
C��;k��`�n���K�*�C�r'_�ꊑ���Ƚ
�08�.%k�@������}����Ǿj̾�2Ⱦڙ��\姾�����/f���,�KL�5 ���V��|��<�VG=~��=X��=���=z��=*3>� >�   �   Zq
>�	>|8>]�=���=���=���=���=�~=D1=XH�< _G�,6˼j�H�DF���k���nܽM|�;����ｏ�ܽ����g��V��~�m��e�*.��Ԥ���޽z���8G���|�	������]Ǿ��Ծgپ-�ԾwZǾ!f��������t���7�-������@������<ƈG=�ә=�0�=,3�=�*�=w$>"H	>�   �   H5> �>��>v��=¤�=�e�=���=.��=���=ڤq=��8=���<XÃ<���:`H;�<1��*4 ���~%���,s�h�鼤�Ӽ\߼�����W�3ަ������S7���}�O9��}�ҾY���'Q��!���+��{/���+���!�x��9����Ͼ�ࡾ��k�.�"����F��<r�^=�T�=�{�=B�=ڌ>�>�   �   R�>�
>�� >�N�=�{�=���=:��=\h�=>}�=:f=�.=�-�<@{l<�}8:�C�t3��,���������H� p����ؼ�����̼6��ԒL��V������fo2���w������.ξ�����q������(��+,��(�����E��]��ݍ˾򘞾�f�{�_����ټ���<4#`=TR�=��=$��=u� >��>�   �   �>���=x��=^�=���=��=�V�=���=ʱu=t�B=�\=^�<� <��7�x_����� �� ��6.�t8��xͼh���tA��T���`Ӽ�,�/R��׽ݽ�<$�� f��Ԙ�6g��ʳ龭����9���"�{Z�h��i:��R龗ȿ�y#���_X�>��1꙽$������<�Yd=	�=3��=�'�=�/�=�0>�   �   (��= ��=%�=��=
�=B3�=��=XPf=��4=�s=(�<H�"< F��8��Xꍼ䡾��<ܼ��㼄�Լ�-��d}����4�p_��e���p�4��^�Ϋ������J��%��O~���Ҿ�G��9���n��������(�����ӾF���x����B�kN��j���w�|~�<$ki=�Φ=z�=�^�=���=���=�   �   ��=���=.��=��=T|�=�s=\C<=l�=L�<@�< �߷��� py�e��twƼ(yռ��Ӽ�W�����8ER�`b» I�9�;@�;  ��5^�^w�@��������'�f�fK���b��rӾϝ뾬q��|� ������q־aT��閾��h�?�&���ӽ�GR�p&���<��l=Z��=�z�=���=�M�=ԟ�=�   �   �y�=6´=��=�x�=��A=�� =�ƀ<�ˠ:0h:�� ��|�Ｎ�����x.���d���n߼\����O�`�w� U�;��S<\��<(á<,��< *�;�fl�R6.��t��ޘ ��T6���o�����V�����þ�wѾ�־�,Ӿm�ƾ�2�������{��fA����������=:�(=�(l=�ǝ=���=2e�=D��=V��=�   �   ��=��=bX= �=��|<���TE���r#�̘Z��ွ@ދ�Qn���b��6�{�,�Z�ک2�@?��������;�'}<pD�<8k=�B=�= ��<h<(�}�z%@��	�����5�n(e� ~���H��t@��x<���ɨ�(=��h����
w�JnI�����B׽p&���Ѽ��;�D=xd=	�=�[�=�N�=p�=(�=�   �   4�u=��4=��< +�:�y��.�E��Q���ɺ��Zٽ��T��%�뽔Uڽ4q���j���uy���.�dɼ����J<��<x-="K8=dYK=b�I="�0= ��<Ȣ:< k��e<��]��r����E#��_G���d�~cy�g��T@���r�B�[�j=�^{�Un뽑¢�̘<�׀�P_2<,	=��S=!�=�Q�=q��=~s�=���=�   �   0�=��<x��x��ˍ��gͽ���o���-��7�rw7�M/�y���
�Z,�ޗ��
,o�0/�pQ�^A<��<��8=�if=��=6��=�qz=�tT=��= ��<������č�`ͽ� �k�+�-�%7�<s7�TI/�>����
�c(�$����(o��-�PR��XA<8�<��8=�ef=��=Ӑ�=
lz=:nT=�   �   H�:<�@k��q<��d��l���J#��dG���d��hy��i���B��o�r���[�m=��}��q뽻Ģ��<�,؀�(b2<�	=T�S=��=�S�=���=�u�=�đ=��u=��4=��< ��:La����E�dJ��º�+SٽJ��O����KPڽm���g���qy���.��ɼP�xB<��<�)=G8=�TK=(�I=�0=�|�<�   �   ��}�0@�L������5�@-e������K��BC��6?��ų�z?��i���9w��pI�|�� E׽�'��Ѽ �;�E=�yd=Q�=]�=TP�=�!�=�*�=��=k��=�iX= �=p}< Ǝ�\-��Hf#�8�Z��ۀ��؋�bi���^����{���Z�<�2�^>�����0��;}<�<�<�f=�==��=`v�<��<�   �   @?.�
z��� ��X6��o�o��������þ�zѾ��־L/Ӿ��ƾ�4���!��s�{��hA��������|��6:�)=N*l=	ɝ=��=�f�=��=\��=�{�=�Ĵ=��=G|�=�A=ؔ =�ـ<@�:@A:� �����N�����*�0����$o߼��(O��x� 8�;8�S<T�<@��< ��<���;��l��   �   ��������'��f��M��e���tӾx��[t��Ȥ �c���2��G ־�U��8ꖾ��h�b�&��ӽIR�p'���<D�l=4��=�{�=��=�N�=v��=��=Ħ�=���=窭=}�=ps=�J<=��=���<��< p������_y�`_��DtƼ�xռ��Ӽ<[��<����QR�0» K�9�ƙ;`�; [��M^��~��   �   ������U�J�L'��0���-�ҾJ��a��p�ғ�����)�-����Ӿ+�������B�MO������w���<Vli=<Ϧ=�z�=�_�=���=��=���=���=�&�=!��=U�=�5�=n��=�Uf=��4=Px=�#�<(�"< ������鍼�����>ܼ��㼈�Լ�3��胆��
5�P~���u�Xq��*�^��   �   �ݽ�>$��f��՘��h��p�龍����:�Ď"�1[����:�>S�ɿ��#��U`X�X��꙽����ȯ�<�Zd=�	�=��=j(�=�0�='1>��>���=���=�_�=`��=���=�X�=6��=��u=`�B=x_=b�<0&< �7�x_����X�����@0�H=�~ͼ¦��G�� �����Ӽ6,��T���   �   �����p2�X�w������/ξ����{r�S��6�(��+,�[�(����E��]���˾ᘞ���f��z�����|	ټ���<�$`= S�=���=���=�� >ו>��>$>N� >�O�=r|�=���=��=,i�=~�=�f=�.=8/�<�|l<�8:�C��4�������0���I��s��(�ؼ8���l�̼���L��X���   �   ���ZT7���}��9����ҾΤ��ZQ�,�!��+��{/���+���!�F�J9�� �Ͼlࡾ�k�0-����� B��<�^=�U�=T|�=��=�>;�>e5>#�>��>���=��= f�=���=;��=���=��q=V�8=��<`<���:�J;�|2���4 ����(&�����s���鼈�Ӽ�߼���ԼW�Yߦ��   �   �����o2�Ίw������.ξo����q����a�(�'+,���(�H��!E��\��Ҍ˾����q�f��y�쒨�xټp��<�%`=zS�=��=���=׵ >�>��>0>[� >�O�=�|�=���==��=bi�=L~�=Ff=��.=�1�<x�l<��8:�C�X0��8����������F�8n��ؼ���P�̼<�� �L��V���   �   *�ݽ=<$� f�Ԙ��f�����,�s��G9�+�"��Y�����9��P�ǿ�"���]X�:���晽���춯<�]d=�
�=���=�(�=1�=F1>��>���=��=�_�=���=��=�X�=���=�u=țB=<a=�f�<81<��7�`�^���������B+�3��sͼ,����=��@����|Ӽ�,��Q���   �   F�����H�J��$��D}��ʙҾ=F��O���m����m���'�l}��ʒӾU��������B�qI��G�����w����<�oi=�Ц=�{�=d`�=4��=P��=���=��="'�=Z��=��=6�=���=�Vf="�4=8z=�(�<�#< ������ލ�Ж��$2ܼ�㼈�ԼT%���u��@�4��G��Z�h�p�<��^��   �   �������'�� f�J��a��'pӾ���1o��*� �?}��R���־�Q���斾�h��&��ӽl>R���� ��<��l=ƻ�=�|�=���=�O�=ޡ�=�=��=���='��=��=4s=�K<=�=D��< < ��� ���My��T���gƼxjռ<�Ӽ�J��pv���/R�P;» {�9��;@(�; T���'^��s��   �   �0.�dq��֖ �\R6���o����&���f�þ�tѾ.�־�)Ӿ��ƾ*0��c��4�{��bA����脩�����m	:0=*/l=�ʝ=_��=�g�=���=���=H|�=LŴ=i��=�|�=��A=�� =�ۀ< 2�:�9:�,	�� ��P�����2$�d��|��x^߼L�h�N���w�`��; �S<� �<�ˡ<���<�K�;`Tl��   �   ��}�n@����\��R5��$e��{��8F���=���9���ƨ�?:�������w��iI�q��C;׽* ��D�м�`�;~L=�~d=�=p^�=@Q�=:"�=
+�=�=���=tjX=��=�}<����<+���d#�Z�Z��ڀ�׋�`g��L\����{���Z���2��5��ߨ���� �;@}<dO�<4p=@G=��=P��<�-<�   �   ��:<X�j�"]<��X������A#�h[G���d�F^y�Vd���=����r���[�e=��v�2f�p���F�<�P���(�2<h	=�S=l��=�T�=r��=�v�=ő=��u=N�4=��<���:(`����E��I��`���MRٽ#��������Mڽ7j��`d��vjy���.�\�ȼ@�� g<x�<3=8P8=*^K=�I=ޣ0=\��<�   �   ��=��<����ྍ�Yͽ����f�i�-�&7�'n7�JD/�`���
���}���o��!��'� ~A<�#�<\�8=�lf=��=��=�rz=�uT=~�=<��<������č��_ͽV ��j���-��7��r7��H/�8��A�
�{%�Б��r!o��%�81�hzA<D$�<p�8=�nf=��=|��=.vz=�yT=�   �   D�u=�4=x%�<���:dL��`�E�sC��U����Jٽ���j���뽭Gڽ�d���_���cy�6�.���ȼ`��g<d�<X1=�M8=n[K=��I=$�0=���<�:<�k�Ze<��]��4���E#��_G���d�4cy��f��@��n�r�d�[�i=�z�tk�k����<��Ȁ�@}2<�	=t�S=���=�U�=���=x�=�Ƒ=�   �   �=!��=XpX=�=0&}<@s�����NY#�B~Z��Ԁ�ы��a��YW����{�R�Z�̚2��2��ܨ���0�;P9}<�J�<�m=LD=T�=���<�<0�}�
%@��	����x5�V(e��}���H��X@��Q<���ɨ��<�����
w�FmI�t���?׽�#����м0I�; K=�~d=Z�=_�=2R�=v#�=�,�=�   �   �}�=8Ǵ=���=k�=pB=R� =��<�V�:�:�0��������0}��ʈ�L��([߼d屮��N�@�w��q�;(�S<��<�š<��<�/�;�dl��5.�xt��Ș ��T6���o�򋔾L���ӑþ�wѾ��־�,Ӿ:�ƾ�2������{�fA��������4���:�-=.l=�ʝ=���=@h�=���=��=�   �   N�=���=���=\��=V��=%s=R<=��=��<@$< �A�`��@8y�L���aƼ�fռ��ӼlK���x���6R�0L» G�9���;p�; ���h3^� w���������'��f�_K���b��rӾȝ뾢q��u� ������C־$T���薾O�h�x�&��ӽ*DR���Ў�<2�l=~��=�|�=H��=$P�=΢�=�   �   ���=��=x(�=��=n�=(8�=+��=�[f=0�4=@= 2�<�#< @�����ڍ������1ܼ�㼴�Լ�(��xy�� �4�@W���a�p�p�T�j�^������~�J��%��J~���Ҿ�G��7���n��������(����ŔӾ���<���8B�4M�����0�w�d��<4ni=Ц=�{�=�`�=���=��=�   �   �>���=���=�`�=���=6��=bZ�=.��=P�u=�B=Hd=(l�<�:< }7�H�^�L~��؞�R��,�85�`vͼ����@@��`����~Ӽ|,�R��ýݽ�<$�� f��Ԙ�4g��Ƴ龬����9��"�wZ�b��a:�nR�zȿ�U#���_X����Z陽����p��<�[d=
�=>��=�(�= 1�=h1>�   �   ��>F>~� >*P�=}�=p��=욽=#j�=�=�f=��.=�4�<��l<�59:�C�0/������|�����\G�o���ؼl���0�̼
����L��V������co2���w������.ξ�����q������(��+,��(�����E��]��Ѝ˾☞���f��z������
ټ���<&$`=�R�=���=���=ŵ >�>�   �   �^>_� >�E�=Bd�=���=%�=�y�=��=�ޑ=<�=L�\=L�;=.=��=���<��<h��<\��<�c�<l�<`x�<0�\<��;�����I�����B��/����þQ��������>��LZ�Cp��a~�ɡ���c~�V4p��Z��>�ǂ�m$���ʽ�fH��0)��������L��<6= {�=�b�=Bg�=Î >�   �   y� >8��=�#�=�W�=���=h]�=P�= Û=u�=�m=VL=��,=��=Hi�<���<D��<$�<(��<<]�<\W�<�Ύ<X�r<P��;@:л����U6���･�=��芾������������:�MGV�o�k���y�:�~�,�y���k�� V�D�:����G��9���f��a�$��A��,@��!�<���=�y�=���=ܹ�=6��=�   �   �=�=/�=���=���=ϯ�=�۪=s��=��=�[=>�7=T�=���<,��<�n�<�H�<��<��v<л�<���<P��<\�<��<0�I< �F������k�rٽ��.�ig��-t��P��A��8�0���J��>_�z�l� 1q�׭l��l_�	�J�p0�k���5龬设�%t����&ǚ��׆�4v�<)%�=�7�=���=���=,��=�   �   ��=0z�=)�=���=���=D��=@�S=`9%=Pv�<$�<��{<��,<Њ�;`;�;p��;�f�;�##<�V^<x�<���<���<$�<�<@8<�J��3�����Y��r)e�����btԾ&���U ��\8�evK�<�W�O)\�3X���K���8�G� �����`Ӿ�˝�qZ��}�⒁�xU�*�
=.��=��=���=*w�=���=�   �   B/�=hQ�=�3�=+��=�GO=��=tʦ<p��;��y���C�dy��T��Զ��(a�� _?��
�����: Q<�A�<�$�<t'�< �<�D�<,ܚ<@{�:p�ټa=��Ms����?��͈��󶾣������7!��T2�So=�:kA���=��3��5"�]���m�@귾�Y��tW:�F߽LE���c:�z=���=�(�=�8�=��=d��=�   �   ^6�=N
�=8�a=nd=x��< t\�@*�����ȫN��o���}�y���d���B�:=�0�ʼ tA��^�:��\<�N�<�=��=��=l��<Dj�<�S��q)��,��[�\�[������¿�n龃�b�����y9#�5K �*�d��Z��׵þ�V���&a����OԬ�"��0�1<:�3=�_�=���=D�=�F�=�=�   �   ޽�=�C<=\<�<�D3�=ܼ�cX����ƽ���G�������S��ֽ�m����Q�h����17��W�;dչ<�=�52=p?=�2=��=�`<p�t�؅[���ѽ�$�V�f�.o��8����)ؾ�&�E� ����ͬ����c�ܾ�쾾����Zt���0�Ϛ�ʌu��<��(M�<гC=�P�=Q��=Q��=�F�=�D�=�   �   p�!=�|<��]���<�d��}�;�&.�_<@�uI��,H���=��u+�	��ٛ�r��:�g��b�@l�`��<8=&	D=�_=��a=PF=�=X�6<�-��u��۽��#���\��e���ţ�+8����ž,V˾U7Ⱦ�޼�����9�p��99����X����  ��(��< �L=Ԧ�=���=���=!Ԏ=��l=�   �   �7<����8�k�X�˽���jg?�Ŷg�E:���X��`7��v��`���y��V�rv.������AT�f��@|#<�=01M=0�y=箅=B[�=��X=F=(8<h⤼�~k�ҁ˽����a?���g�7��AU��4���r��;]���y�ґV�s.�x|�[����<T��`��P�#<l=�/M=��y=��=�X�=��X=d>=�   �   �B��2u��۽ˠ#�H�\�i��ɣ��;����ž�Y˾�:Ⱦ⼾y�����Ƌp��<9����/��x�� 3�����<�L=ާ�=��=���=�֎=<�l=��!=h7|<p�]�dz<��[���s��5��.��6@��I��'H��=��q+����3��4���<�g�`[�@�k���<B=D=
�_=��a=�JF=
=��6<�   �   �[���ѽ8$���f�1r��� ��F-ؾ�*�H� �����������d�ܾﾾ����]t�*�0��潐�u��@��4L�<~�C=�Q�=���=��=�H�=�G�=c��=~L<=�P�<�?0�X!ܼ�SX����ƽ���V����������ֽ1h��������Q�����x'7�`_�;�Թ< =l32=�?=& 2=�{=�_<Xu��   �   O2������[�.����ſ���h!�b�����u;#�M ��+�������ַþtX��)a���,֬�����1<��3=�`�=���=��=�H�=k��=B9�=��=~�a= n=�Ǉ<�[���� ����N�&�o���}��~y���d�D�B��6���ʼhA� ��:`�\<M�<�=��=�=D��<�^�<����z)��   �   �x��(�?�Ј�A�����羦��i9!��V2�9q=�mA���=�V3�E7"�{��fo龗뷾�Z���X:��߽�E� �c:{=��=�)�=�9�=���=B��=�1�=)T�=37�=�=<PO==�ަ<���;��x�H�C��e����������T��@L?�`��۷:�S<A�<"�<T#�<Ty�<�=�<,Ӛ< ȩ:x�ټ�A���   �   ����,e������vԾz��8W �u^8�xK���W��*\��X���K���8�%� �����aӾ�̝��qZ�n~�G���@U�ı
=���=k�=���=Zx�= ��=��=<|�=�+�=~��=���=���=��S=�@%=T��<��<�{<��,< ��;0\�;���;`v�;h'#<�V^<�v�<���<���<��<`۞<�'<hK���3�����   �   %�.��h���u��7��S��c�0�͚J��?_���l�2q�خl��m_���J��p0����Q6��设�%t�����ƚ�ֆ�Dx�<�%�=\8�=N��=r��=< �=0?�=�0�=\��=d��=ڱ�=ު=ˠ�=E�=�[=��7=��=��<H��<�s�<HL�<P�<��v< ��<ԩ�<��<��<<�<�I<��G�p���,k��ٽ�   �   C�=��銾�������Ń���:�HV�,�k���y�ң~���y�"�k�� V�d�:�����G������e����$��@���<��$$�<y��=Nz�=,��=���=��=ڱ >��=�$�=�X�=��=�^�=��=5ě=��=D�m=BL=��,=��=k�<���<���<��<��<|[�<(U�<�ˎ<h�r<P��;�Oл,���f8������   �   �B�T0��h�þ���ښ�J�>�MZ�QCp�b~�ʡ��rc~�$4p�zZ�K>�n���#��>ʽ��G��5)����������<�7=�{�=Hc�=�g�=�� >�^>�� >�E�=�d�=��=P�=�y�=��=�ޑ=&�=�\=��;=�-=4�=h��<\�<��<��<xb�<��<�v�<��\<��;������NJ��a����   �   ��=�銾�������������:�GV��k�z�y���~���y��k��V���:�2��NF�����e����$�'?���7���'�<��=�z�=|��=º�=��=� >,��=�$�=�X�=(��=�^�=��=Xě=��=��m=�L=X�,=��=<m�< ��<\��<��<d��<_�<�X�<�ώ<8�r< ��;P=лܸ���6������   �   ��.�&g���s�����׉���0���J��=_�~�l��/q���l��k_�ԱJ��n0�[���3�箾�"t�l���Ú�l̆�(�<'�=69�=���=��=� �=b?�=�0�=~��=���=���=7ު=���=��=8[=��7=��=���<ؒ�<�w�<Q�<`�<��v<���<���<���<��<�!�<��I<��F�L����k�ٽ�   �   v��@(e�ۢ��FsԾn���T ��[8� uK���W��'\��X���K���8�Ͱ ����4^Ӿʝ��mZ�V{�����`:���
=q��=��=p��=�x�=���=��=x|�=�+�=���=Ѻ�=ݘ�= �S=�A%=��<��<8�{<� -<@��;Ps�;p��;���;8#<�h^<��<��<���<�<|�<H@<��J��3������   �   �p���?��̈�0򶾽��Ѻ�<6!�>S2��m=�biA��=��3�4"�����j龥緾ZW���S:�i߽��D���e:�='��=	+�=�:�=T��=���=�1�=jT�=o7�=!��=�PO=�=�ߦ<��;��x���C�Pb��8�����N��P<?� ͸��z�:@i<\L�<�-�<h/�<��<K�<�< ܪ:��ټ];���   �   \)��I���[�ͻ��t�������������|7#�/I �(�{����쾲�þ3T��9"a����ά� ��(2<�3=�b�=R��=��=VI�=�=�9�=�= �a=�n=dȇ<`�[�d��6��|�N���o�µ}�h|y���d���B�@2��}ʼPRA� J�:�\<�Y�<�=��=j�=���<�q�< 2��l)��   �   �~[�#}ѽ	$���f��l������j&ؾ_#�\� ����Ū������ܾ
龾���JUt�T�0�0��8�u�(��P^�<�C=�S�=;��=>��=�I�=&H�=���=M<=�Q�< '0�| ܼ�SX�W���ƽ�㽙���*���_�\�ֽVf��w�����Q�����7����;��<�!=�:2=�
?=�2=��=(`<8�t��   �   `��$�t���ڽs�#�Z�\�Pc���£��4��H�ž^R˾3Ⱦۼ�~���꒾�p��49�@�����Ο�����l��<v�L=&��=���=ڼ�=�׎=B�l=p�!=�9|<��]�z<�q[��Vs��5�{.��6@��I�'H���=��p+����(�������g��O뼠�k��Ó<�=D=��_=��a=~TF=�=@7<�   �   x"8<tѤ�Ftk�?{˽���]?�3�g��3���Q���0��oo���Y��w�y��V��m.��w�L����.T�PI����#<�=7M=^�y=e��=H\�=�X=�F=�	8<l᤼�~k���˽����a?���g��6��*U���3���r���\��L�y��V�(r.�l{�����7T��U����#<�=6M=��y=��=m]�=|�X=�K=�   �   �!=8V|<��]��n<��T��Uk�21�n.�"1@�I��!H�F�=��k+�Z��ٌ������vg�PB뼠9k��ɓ<R=TD=��_=V�a=�QF==��6<p,���u��۽�#���\��e���ţ�8����žV˾37Ⱦ�޼�d����풾,�p�99������8���[�����<��L=���=��=���=�؎=\�l=�   �   Ă=S<=8a�<��-��	ܼ:FX����V�ŽB�㽢���G������ֽ{_������2�Q�Hq�� �6�0��;��<�"=P:2=�	?=�2= �=x`<��t�\�[�j�ѽ�$�J�f�(o��4����)ؾ�&�@� ����¬�����3�ܾJ쾾^���Yt��0���潾�u�4��TV�<��C=lS�=Y��=⴮=�J�=�I�=�   �   �;�=��=<�a=&v=�ڇ<��Z�����4��ƎN���o���}�Poy���d��B�|)��oʼP=A� ��:��\<\�<�=L�=$�=���<�l�<0M�Bq)�_,��I�J�[������¿�l龂�b�����v9#�/K ��)�T��+�쾝�þ�V��.&a�����Ҭ����2<L�3=b�=.��=9�=.J�=N��=�   �   J3�=HV�=�9�=��=�WO=�=��<p3�;�1x�ТC��M���ힼ@����>���"?�������:0s<4O�<�.�<�.�<d��<�H�<�ޚ<@��:,�ټ-=��*s����?��͈��󶾠������7!��T2�To=�8kA���=��3��5"�P��ym�귾OY���V:�߽��D���d:�}=C��=�*�=�:�=���=���=�   �   ��=�}�=f-�=���=G��=���=r�S=�H%=���<��<8�{<H-<P��;��;0��;��;PB#<@o^<���<�<��<��<��<�;<��J���3�Ս��L��g)e�����_tԾ&���U ��\8�evK�=�W�P)\�2X���K���8�<� ���d`Ӿ�˝��pZ��}�쑁�M�v�
=p��=#�=T��=0y�=��=�   �   �?�=l1�=���=���=���=�=��=��=�[=r�7=X�=��<��<�~�<W�<��<H�v<�Á<б�<���<��<@!�<��I<��F� ���pk�Yٽ��.�dg��*t��O��@��8�0���J��>_�|�l��0q�׭l��l_��J�p0�d���5龔设a%t�T���ƚ��Ԇ�(y�<�%�=�8�=���=؎�=� �=�   �   � >b��=$%�=RY�=���=x_�=��=aś=��=�m=DL=��,=��=0q�<���<��<�<��<D`�<�Y�<dЎ<��r<���;08лD���@6���｢�=��芾������������:�MGV�n�k���y�:�~�,�y���k�� V�B�:����G��-����e��@�$�|A���>���"�<$��=z�=��=���=��=�   �   d��=���=$��=� �=���=�K�=�=���=�=�"i=U=�QG=8>=h�9=��9=��<=� B=�
H=�XK=��G=�6=�@=���<� ���<D�b.׽
A;�Ry��n�Ѿ^����8���c�v���k����;�������ⴿ����t0��j�����\�b�(�6��`�e˾�ƈ��$�9 ��(M5�8|=�Z�=J��=Ԫ�=�d�=�   �   ��=FF�=s�=�[�=࿼={&�=�=�.�=�i=��P=��==R1=�!*=P_(=�
+=�*1=��9=@B=�H=��F=� 8=`�=,��<`4»޾9�D�Ͻ$T6��%��,b;���F5���_�[����▿T��阮��α�E����S��ɖ�+L����^���3���	�LPǾ_Ʌ�T��؆���~��/=n��=b��=��=�x�=�   �   �d�=�P�=8��=�·=bZ�=�;�=h=@=�= �=R�<��<l��<�W�<�p�<>�=��=z0=>�==HC=��:=��=���< ���C�$��	(����G�����E�*��S��!{�����✿�¥��ڨ�zإ�����Y!����z�� S�c�)�����z��2=z�ʼ�Q��0���ң%=*�=F��=,R�=Ȗ�=�   �   bb�=k(�=��=�p�=��d=�$*=x�<�0�< ��;�Dk:������ 3�9���;�Y?<�<��<,q=�7*=;=:�==l6*=pA�<�l�; i׼�W��n���j�2Ŭ�	���:�@�@Ae�ق�C����뗿�Ӛ�������ٚe���@����J�뾟���N_�l� ��xX��'F;�5=�|�=�P�=,��=N\�=�   �   �=�	�=Hs=l*=>�<��j;=c�b꼀9"�V=���D���9�>��t	�^���_n��!<\�<�
=�u,=<�==��7=,�=�L�<`?>��a�;��r�D�@���<�;v
�}�(�NiI�֌f�+�}��B���ꈿ����t~��g� XJ�"k)�<c��<;�ԑ��j=�pҽ�����G<��F=�Օ=~�=���=^&�=�   �   x��=��I=��<�X; ��ZD��o��⥸�|�Խ���㽐�ֽ����娛��9g��u�hmo�`c�;�<j�=�6=BqB=ʌ/=�r�<�Ğ;@��>������מn��A����� ��l�)��=C��[W�
gd��i��e�T{X��D�w+����n�U���o�.���睽�W��\γ<W=k�=6�=Ĭ=�G�=�   �   ��*=�:�<�vL��:�z��eR���T�.��c@���H���F�,K;�>�'��b���޽RA��8�A�|t�� �;�+�<��&=�G=R�H=V�%=D?�<P����O��ڽ��3�}���j����⾾	��k��f/��w:�h�>�\9;�?�0�D[ ��^��y�����ه���:�1<�0?Q� t��8��< �c=Z!�=M��=�o�=x{v=�   �   �1;<h��ē|���ؽg���J�`t�4��ij���;�����<F��
���]�,3���7d����L�������M<9=.9D=��[=(:O=
x=�~v<ܖ������-����=������竾�tҾ� ���n��������q��1
�����ؾ����޽��#OL�=������ ڼ�"8<��=lpi=y=�=Q�=sc=��=�   �   ��ļh$���$��%�5�ds�����V��;NɾG�׾L�ݾ�ھt�;)���U䟾�ۂ���I�>n�Z����.�����\��<
7=�g=�r=�=W=�=Я4<�jļ�����h�5�c]s������R���Iɾ��׾��ݾ]ھj�;����F៾;ق���I�Hk��U��(�.�������<�
7=�
g=Fr=�8W=��=h�4<�   �   p���6���>�ȋ���뫾EyҾ�%��cq����1��ct�	4
����q�ؾ�ò����lRL���� ����
ڼ�8<�=�qi=�>�=��=,yc=��=h[;<e����|�ݘؽ����J�?t�h����f���7��E���B�����y�]��'3����?_����L�����P�M<�9=08D=`�[=$6O=Dr=�_v<�����   �   �"ڽ@�3�c���������	�|n��i/�Xz:��>��;;���0�^] ��`��|�Y����ۇ��:�s?�.CQ��������<�c=�"�=$��=r�=@�v=6�*=�P�<0AL���:��p���G�O��2�.�F]@�t�H�ӾF��E;�U{'��^�Ӗ޽�;��8�A�li�� :�;/�<z�&=n~G=`�H=�}%=�2�<8	��O��   �   �����n��D��'������)�$@C�3^W��id�i!i�`e��}X��D��x+�G��p����`�o�����靽�[��xͳ<�W=\�=��=$Ƭ=fJ�=��=��I=�$�<��X;����C��f��R�����Խ��ъ� ~ֽꤽ�i����.g��m�HUo� ��;���<6�=��6=RoB=��/=i�< ��;��� ����   �   "�D�����(�;5���(��kI�F�f���}�D��숿����$v~���g��YJ�al)�1d�>;�Ց��k=��qҽ:��(�G<p�F=�֕=��=x��=�(�=��=>�=�s=,*=PT�<�Tk;�c�pE��*"���<�&�D���9����P�� O��@ n���!<��<\�
=v,=4�==|�7=ή=C�<�X>���a�����   �   r�j�XǬ����5��@�<Ce��ڂ�X����엿�Ԛ��������
�e���@�K��K��I���O_��� �hyX��+F;�5=w}�=�Q�=���= ^�=zd�=�*�=��=,t�=��d=�-*=�!�<�D�<���; �m: J��� �9�2�;(o?<��<���<�r=N8*=X�;=��==64*=;�<0I�;�t׼�[�����   �   X������*����*���S�|#{����h㜿xå��ۨ�"٥�0 ���!����z�C!S���)����z��c=z�ļ��P�������%=�*�=��=6S�=��=bf�=�R�=F��=�ķ=]�=t>�=\	h=�@=��=d�=8^�<��<��<�_�<8w�<��=@�=20=@�==jGC=��:=��=���< ��H����T(��   �   '���c;���.5���_�����㖿�T��\����α�����&T��:ɖ�@L����^���3���	�
PǾɅ����څ���w�,1=6�= ��=���=dy�=��=\G�=8t�=�\�=H��=(�=��=D0�=H�i=��P=��==�1=�#*=�`(=&+=L+1=ԉ9=@B=BH=�F=��7=��=x��<0M»��9���Ͻ�U6��   �   �y��;�ѾӬ���8�p�c����������;������ⴿ����T0���i��ޢ����b���6�p`�Dd˾Bƈ�j$�w��PB5�Z~=�[�=���=\��=Fe�=���=��=r��=!�=��=�K�=8�= �=�=�"i=��U=:QG=�7>=��9=�9=̷<=& B=�	H=XK=�G=��6=F?=h��<`2��^?D�0׽$B;��   �   8&��eb;��L5���_�D���d▿�S������5α�Ԟ��nS���Ȗ��K����^�Î3��	��NǾLȅ����-���n��2=��=���=&��=�y�=��=pG�=Ft�=�\�=V��=(�=��=T0�=|�i=�P=��==@1=F$*=�a(=�+=6,1=Ҋ9=0AB=|H=8�F=8=B�=@��<�:»�9��Ͻ�T6��   �   �������έ���*���S�,!{����✿¥�	ڨ��ץ������ ��Z�z�OS��)�����x��Z:z�����M���w��4�%=�+�=ާ�=�S�=`��=�f�=�R�=h��=ŷ=$]�=�>�=�	h=�@=��=��=|_�<���<8��<tb�<Dz�<T�=2�=R0=��==�IC=H�:=��= ��<�h�C�����(��   �   ��j�lĬ������C�@�@e��؂�j����ꗿ�Қ�~���쏿����e���@�
�����{��YK_��� ��pX�`�F;�
5=�~�=�R�=4��=|^�=�d�=1+�=�=It�=*�d=�-*=\"�<�E�<���;��m:�;�@�� ؉9�@�;�w?<���<(��<�u=�;*=��;=��==~8*=E�<Pz�;`e׼�V������   �   ��D������;t	�8�(��gI���f��}��A���鈿I���q~���g��UJ� i)�~a��9;5ґ��f=�1jҽ���X�G<��F=}ؕ=��=H��= )�=L�=��=�s=f*=�T�<`Xk;�c��D�\*"��<��D�z�9�4�����I����m��!<���<4�
=Bz,=̇==��7=�=�Q�<�3>�za�����   �   ���"�n��?��6�ྉ����)��;C�,YW��dd�i�e��xX�w�D��t+��	�k�Q ��%�o�F���᝽\D��޳<�%W=c�=�=Ǭ=K�=i��=N�I=�%�<��X;h󷼤�C��f��$���h�Խg�D��H}ֽ����C���6,g��j�@Go����;$��<Ȳ=��6=uB=>�/=Ty�<0�;�|�A����   �   'ڽ��3������������	��i��d/�u:���>��6;���0��X ��\��u羀����և�ڙ:�v4��2Q��$�����<�c=�$�=���=	s�=~�v=
�*=�Q�<�?L���:��p���G�B���.�(]@�F�H���F�OE;��z'�!^�v�޽a:����A��a��`\�;d8�<��&=H�G=<�H=H�%=�G�<���L�O��   �   L����'����=�*���嫾nqҾ����l������Zo�?/
������ؾ��������IL�����8�ټ�I8<.�=�wi=�@�=��=�zc=��=X^;<d��F�|�Øؽ���xJ�7t�a���vf���7��+���B��̾����]�1'3�ԙ��]���L�p���h�M<�>=�=D=�[=L>O=�|=`�v<X����   �   �Yļ^������5�Xs������N���Eɾ?�׾�ݾ�ھߗ;J���[ݟ��Ղ�ďI�Df��M��z�.�`I��t��<�7=g=zr=^@W=��=�4<Tiļ���[��_�5�^]s������R���Iɾ��׾��ݾIھM�;j���៾�؂��I��j�6T��l�.� �����<�7=�g=�r=bBW=H�=��4<�   �   �y;<�Q��bw|�<�ؽ��J��	t������b���3��N���>��V�����]��!3�b��pV���L�y��HN<^B=�?D=��[=n=O=>z=��v<���i���N-����=������竾�tҾ� ���n��������q��1
����ݍؾ���������NL����F�����ټ�28<��= vi=�@�=��=~c=��=�   �   �+=a�<�L�(�:�i���>���n�.�W@��H�Z�F�R?;�Tu'�&Y��޽A3��R�A�P��@��;lA�<l�&=��G=N�H=�%=�B�<���(�O�Iڽ��3�v���h����⾿	��k��f/��w:�g�>�Z9;�9�0�;[ ��^��y�ۺ���ه��:��:�(<Q��X��@��<җc=J$�=��==t�=z�v=�   �   ���=� J=�5�<�vY;8۷�n�C��^��B����}Խ�㽗���sֽa��������g��_�0$o��ؤ;��<"�=��6=�uB=
�/=�v�<pО;R���������Ǟn��A��������n�)��=C��[W�gd��i��e�Q{X� �D�w+����n�$����o�����杽8R���Գ<#W=��=H�=�Ǭ=�L�=�   �   �=��=s=*=@g�<�l;��b�*�2"���<���D���9�`����(6���Mm�(�!<���<Ԑ
=�|,=0�==,�7=��=�O�<;>�T�a���b�D�:���9�;v
��(�OiI�ٌf�0�}��B���ꈿ����t~��g�XJ�k)�.c��<;hԑ�-j=�#oҽ��� �G<��F=�ו=��=���=<*�=�   �   �e�=�,�=L�=w�=��d=|5*=�3�<�X�<@6�; �p: ���_� ^�9 ��;Г?<��<���<dy=>*=��;=��==�8*=E�<Pv�;�g׼hW��[��	�j�/Ŭ����;�@�AAe��ق�C����뗿�Ӛ�������՚e���@����5�뾂��vN_�� �RwX� EF;�5=!~�=�R�=j��=&_�=�   �   >g�=�S�=���=�Ʒ=-_�=�@�=h=�"@=J�=x�=|l�<`��<��<m�<���<6�=Z�=� 0=f�==@KC=6�:=��=���<�W�C����	(����D�����E�*��S��!{�����✿�¥��ڨ�zإ�����Y!����z�� S�^�)�����z��=z�����P������F�%=�*�=i��=�S�=���=�   �   (��=�G�=�t�=�]�=5¼=")�=��=�1�=��i=�P=>�==z 1=R'*=�d(=z+=h.1=��9=�BB=�H=H�F=8=2�=P��<�1»��9�0�ϽT6��%��+b;���E5���_�Z����▿T��阮��α�F����S��ɖ�+L����^���3���	�DPǾUɅ�:�������|�,0=���=���=���=|y�=�   �   Da�=�?�=���=9:�=�H�=E=f^�=�c=��H=y6=�?-=B�,=��3=�VA="QS=j�g=bR{=Z��=��=K;�=��l=�/=,��<xl��������!��܇���ξj��B5E��N|�i���z���eͿD�i�ם�h��0�x'Ϳ���K���vz�[�B�����Ǿ�f�����9`�@�;dfN=�u�=���=�	�=�   �   dv�=8��=���=]}�=X�=%܈=DGh=��D=d�(=zp=�=��=ޑ=V()=@�>=�lV=��m=��=|��=FP�=��k=��1=�0�<�)��7p��Bt�����?Tʾ���.�A���w�궗�Ja����ɿO�ܿz�W�쿦��ׁܿ��ɿ�������v�Eh?��L�7�þ0�y��
�NiV�( <jP=�=���=���=�   �   X��=r"�=���=:ږ=�|x=6�B=-=�'�<\�<�P<(�6<�6O<L�<l��<X�<� "=�iD=�#b=�%v=��z=�$h=�X6=��<�a�`���d���#w������G�6��j�P���G^��]⿿��ѿ�ݿ��0ݿ��ѿz���$@������fi��)5��`��8���i�������9�XD<��U=��=���=��=�   �   ��=͒�=��=TH=`=��j<@h��@�l���ü���T�ռH<���.�`�;�ҍ<T��<�',=��P=*td=0`=P�;=�i�<0/��8$Z�w�����Z��&������t&�Z�U�����A��o(�������?˿ Ͽg|˿F��f����y��`���ZuU��%����M륾�3O���ڽ��,J�<B�\=��=d��=��=�   �   �=��_=R�= �N<�87�L����d�n���ޮ����dι��̫�a���d�a�,4�p���l�;x�<�z=�A=(.Q=`�?=�=�D�;$��{�Ž,�6��\����Ӿt��*�;�7�g�?���������Y�������ᴿA���Ǹ���̉�A�h���;�>���Ҿv���Lz.�=Ԯ�0�$��<��b=�1�=|�=K��=�   �   �o:=���<������e���1�Ͻ�����z.�-�5�i3�S�'�R7��$��5W���wy�h3�\����<�4=�8=r>=��=\،<�f��R�������j�eǮ�v��S��AdD���i�@���G����������^���������9k�L�E���U+��%��Lti���	�B�{��߻�~=�e=�7�=~�=��{=�   �   �ao<���.uf�Yr˽��&HA��)j��������@��:ʒ�.�j�v���Q��2'��;�������0%��\���ؓ<D="V4=T?,=���<���:� #��Ƚ*E1�<Q��3��l#��bT���>��Z�}�p���N*��\���Er���\���@�"t!�d� ��Rþ����N�3�
bȽ4����;��=��`=�gv=lv_=�=�   �    4��b��]��z6��Tt�>����3���Hʾ��ؾ&�޾
�ھ�>ξ�⹾�ʟ��P����G����w��n�$������<\�=8C6=F$=P��<�7C��l�BX��E�m��,¾)f������+�.�=�ލI��M��uJ��e?���-��T����}Ǿm��R�N��R �AY����h�E�<�[-=�-T= �J=>Q=��<<�   �   z���D_���G������� ܾ
 �|����X�����N����0E�-Һ����V�U�Ҹ����X��� ��;���<�6=��==��=0�_<ଫ��؊�XZ�w�G����i��	ܾ> �y����K�����gK�8��A⾾κ����-�U�ȵ����Ի��@��;���<~�6=��==��=X�_< ī��   �   �`�BF����t¾1k��´���+��=�E�I�n�M�$yJ��h?�3�-�!W�����"�Ǿ�����N��T �1\���i�C�<�\-=�0T=��J=xX=8 =<��������"�5�\Mt�����4/���Cʾ��ؾ��޾�ھ[:ξ�޹�*ǟ��M���G�����r��P�$�����"�<*�=A6=�=���<�]C���l��   �   �I1�ET���6��(��W���>�g�Z��p�R�,������Hr�v�\�O�@�v!��� �Uþn�����3�eȽf7����;�=��`=lv=�|_=F�=Ќo<X{��df�
h˽��=AA�)"j�k���������1ƒ�p퉾��v�ϔQ��-'�<4��ܮ��b(%��/���ߓ<p=VU4=�<,=���<@��:2+#��Ƚ�   �   �k��ʮ�e����gD���i�+B���I��^���\Ý�������P��*<k�.�E�y��-�'���vi�R�	�n�{�p߻<=�e=�9�=��=h�{=nx:=���<�9��`���v�Ͻ������At.���5��b3���'�2�����O��ly�V*��'�� �<(7=8=>=��=�͌<v���������   �   _����Ӿ_��t�;���g��@��/��N�����������O㴿���������͉��h��;�3��M�Ҿ\���l{.�sծ�����<��b=�2�=x�=�=s�=J�_=��=�O<��6�&��.�d����ծ���� Ź�ī������a�)����0��;���<�}=4�A=�-Q=��?=��=`�;�����Ž̟6��   �   �(��T���/&�h�U�E���C���)������@˿sϿ�}˿\��U���]z������JvU�D%�����륾�4O��ڽ���K�<��\=��=���=��=,�=���=o��=<
H=�'=�k<�ش�x�l��üD��D��t�ռ�&���	��%�;�ލ<t��<
+,=��P=�td=f/`=J�;=c�<�W��^+Z�i���ܬZ��   �   ��������6���j�?᏿H_��j㿿��ѿ�ݿu´1ݿ��ѿ����@��m���gi�*5��`�9���i�`�����9�pD<f�U=��=��=,�=&��=�$�=z��=3ݖ=N�x=��B=*5=�8�<���<�P<�7<�TO<���<� �<�#�<2"=�lD=z%b=V&v=ԅz=�#h=�V6=���<� a���������&w��   �   �Uʾ���:�A�%�w������a��{�ɿ�ܿ�z�١���%�ܿ��ɿ�������v�'h?��L���þ��y�W
�gV��'<�kP=��=���=���=�w�=|��=��=�~�=�=ވ=fKh=ГD=��(=�t=��=��=Ɣ=�*)=(�>=�mV=��m==��=i��=�O�=��k=ܣ1=T+�<01���r���u�ݶ���   �   �ξ����5E�]O|�]i��H{��fͿ@D�i�ٝ�h쿷0�='Ϳy������luz���B����Ǿde����(6`���;ZhN=�v�=,��=X
�=�a�=f@�=��=�:�=�H�=�=�^�=Hc=��H=y6=�?-=�,=R�3= VA=xPS=��g=�Q{=㊅=V�=�:�=��l=n�/=䣐<�q��a����!�n݇��   �   �Tʾ���K�A��w�߶��-a����ɿ�ܿ�y�٠���6�ܿ�ɿ
������v�Ag?��K���þ��y�D
�dV�0<DmP=i�=���=���=�w�=���=��=�=)�=ވ=jKh=ܓD=��(=�t=�=4�=,�=B+)=��>=�nV=l�m=���=ף�=tP�=��k=N�1=/�<<,��q���t�����   �   ߾�������6�b�j��ߏ��]���῿�ѿݿ���/ݿ��ѿr�'?��*����di�Y(5�b_�7���i�@���@�9�8)D<�U=��=���=��=a��=�$�=���=Bݖ=`�x=��B=65=9�<���< �P<�7<�VO<���<T�<�%�<T"=�mD=�&b=�'v=Ƈz=$&h=jY6=��<�a�J���M��t#w��   �   
&�������&�b�U�y����@��~'������_>˿��ο
{˿�������Ux��;���XsU��%����饾|0O�X�ڽ���V�<��\=3�=̜�=�=��=2��=���=p
H=�'=k<�մ���l���ü���L��(�ռ%��`��0�;��<��<-,=��P=Xwd=�2`=:�;=m�<0#��`"Z�?�����Z��   �   �[���Ӿt��٧;���g�>��m��T�܊������3ി����9���Bˉ���h���;�[���Ҿ����v.��ή��஼\��<�b=�4�=v�=���=��=��_=�=PO<8�6���&�d������Ԯ������Ĺ��ë�,���εa�z'� �� ��;T��<��=f�A=�1Q=X�?=��=�Y�;��j�Ž��6��   �   *�j��Ů������WbD�C�i�)?��^F������违����V���R���6k���E���h'�"��Zoi��	�v�{��޻��=�e=@;�=�=д{=Vy:=��<�6��.��ݱ��o�Ͻ������8t.���5��b3�X�'��1����N��jy�(�0��8�<�:=<8=H>=H�=lߌ<�^������+��   �   hB1�[O���0��8 ��eR�J�>�P�Z�h�p�f��(�����GBr�b�\���@�lq!�� ��Nþ����w�3��ZȽ4(��+�;��=�`=�ov=�~_=�  =`�o<Tz���cf��g˽	��?AA�0"j�l���������$ƒ�Z퉾x�v�{�Q�\-'�B3�������%%� ����<�=�Z4=XC,=���<@O�:�#��Ƚ�   �   �R���E����¾Nb������+�5�=���I���M��rJ�yb?�f�-��Q������xǾ�����N�N �R����h��W�<�c-=�5T=P�J=�Z=�%=<X���������5�]Mt�����9/���Cʾ��ؾ��޾�ھJ:ξ�޹�ǟ��M��t�G����rq��l�$�����*�<V�=�G6=�(=`��<�C���l��   �   �ӊ��V���G���� ���ܾ� �cv����F}����nH�j���;�<ʺ� ����U�������X���p,�;���<��6="�==��=��_<�����؊�>Z�j�G����k��ܾA �y����N�����bK�/���@⾖κ������U�:������������;��<��6=�==~�=p�_<,����   �   D��������1�5�NGt�]���+���>ʾ��ؾ̌޾��ھJ5ξ�ٹ����I��X�G�
���i���~$��;�`6�<� =I6=F(=���<(1C��l��W��E�f��,¾+f������+�1�=��I��M��uJ��e?���-��T������|Ǿ<����N�R ��W��x�h�\M�<a-=5T=��J=^=�<=<�   �   جo<�f���Vf��_˽��V;A�bj�����|����������Q鉾��v���Q�~''�i)������,%�@���@��<N=V]4=PD,=l��<���:�#��ȽE1�2Q��	3��n#��cT���>��Z���p���P*��b���Er���\���@�t!�T� ��Rþ������3��`Ƚ>1� ��;�=��`=4pv=p�_=x =�   �   �~:=���<�䠻Pu����"�Ͻ�������m.��5�;\3��'�,�����E���Zy����ę� )�<@=�8=B!>=��=�݌<Lc��Ϧ������j�_Ǯ�s��U��BdD���i��@���G����������a���������9k�E�E���7+��%���si�z�	��{���޻��=�e=L;�=��=��{=�   �   ��=�`=��=�.O<��6�&��F�d�@����ˮ�>�G���l�������0�a���(��P��;0��<4�=��A=v4Q=ک?=0�=@U�;����Ž�6��\����Ӿt��+�;�9�g�?���������[�������ᴿC���Ǹ���̉�<�h���;�5��ֈҾS����y.�dӮ�����<��b=B4�= �=虡=�   �   ���=8��=O��=TH="0=8<k< q���l�h�ü���dr��ռ���8���}�;D�<���<v2,=�P=fzd=�4`=��;=Hn�<`#��L#Z�/���p�Z��&�����s&�Z�U�����A��q(�������?˿  Ͽh|˿G��h����y��`���VuU��%����4륾�3O���ڽ��pN�<(�\=��=���=��=�   �   %��=�%�=@�=gߖ=��x=��B=4<=\H�<\
�<�P<(<7<�wO<x�<��<82�<�
"=prD=�*b=�*v=�z=�'h=�Z6=��<�
a����N���#w������F�6��j�O���G^��^⿿��ѿ�ݿ���0ݿ��ѿ{���$@������fi��)5��`��8���i�8�����9��D<��U=��=g��=��=�   �   �w�=���=���=��=D�=t߈=�Nh=z�D=��(=�x=:�=j�=4�= /)=�>=�qV=�m=���=ʤ�=HQ�=L�k=��1=2�<�(��p��6t�����<Tʾ���.�A���w�鶗�Ka����ɿP�ܿz�W�쿧��ׁܿ��ɿ�������v�Bh?��L�/�þ�y��
��hV��"<
kP=��=z��=���=�   �   ��=>x�=鋶=��=F�=g=H�;= =l�<�B�<���<���<��
=��&=�G=�j=��=�/�=9T�=�Đ=��w=��$=���;d�9��]��~"f��̺��a��HC�����R�� �ǿ�X�ȴ�����4I�����������ƿ���5T��7c@�oV��E��
�W��սh)���<���=f�=T*�=�   �   ��=꨽=ܶ�=)�=.�y=� G=j�=��<�u�< ��<���< X�<���<�w=��,=�S=��w=�1�=R�=���=�=u=�%={�;��0���
�`�:϶����Ş?�<�~�z��y5Ŀ�t����O����P����L��b���Wÿ�_��S9|��<�j��:���d�R�nrϽ�AѼ��<G�=ʟ�=��=�   �   �ǳ=��=�=Ηc=DR$=���<�/< "G��s�p�R�*P��@��E��<Xϳ< [=,8@=��i=��=�݃=�gl=rz'=h0<�4�D�ٽ��P�c>��x� �B�4��4q�4���j���+ڿ�T���]�
���9�r���{�Xl��Z�ٿ�빿�q���Lo��2��Q������ D�𪼽læ�T��<J�|=���=���=�   �   ��=Fz=@�6=�w�<`g�;�Ԉ�d��ZO��z�Z܆����ʥm���=�@M��P1W� ��; ��<�r=�gN=bAe=��[=�E(=X_|<Rܼ������7��>���E�&d$��\��?��'��v�ȿ��<���P�����~�����/��ȿr���󋿘�Z�"�"����,ᔾ -�>���(RM�
G=�?u=*	�=�U�=�   �   |�P=<�=p� <����+J����Tս& �М�����C�a����l������(���:�8<H<$�<�1=P�@=l�$=䷨<�u�yC����j����ȾKZ��&A��sw�Q�������ɿ<ܿ��k��迁�ܿ.qʿ�ײ����&�w���@�����ƾ��nA���v� K�$=25g=�=V�=�   �   ���<��Jr+�<��������&��L�F$j�`~�H��׀�%q��CV��3�$]��<ǽ�q�`�Ƽ���;t��<$�=�= C�<`	�&-C�!��dR��C���Q�n�"���Q��=�����&���U����ǿ'�˿�iȿTM��f=��h������GS��]#�\�����u�N�I�߽&8'��!�;4&=n�O=��T=�X*=�   �   �M��bQj�>Qٽ(�$� L_�4d���G������Ⱦ�ξ��ʾq���`:���|���m��X3������������!�:(�<lz=���<�$<Dtͼ����Cm�&����?��n�Ļ*��S��E{��(�����}���J���������7k����}��V�ޙ,��x���B���Pv�����H宼py�<�=��,=�X=�Qo<�   �   �?�����
�>�uQ���(��L"ԾH*��:�	�����H����<c�m��ھǋ��4؋��aK�m����H0��`�;Ph�<,��<���<��|��X8�5ս�o:�͵����Ⱦ^z���%�yLF�f)c�sz�
z��<��G��|��e��I���(����w�̾�����P?���۽�>�@�^���<�=h��<�L<�<���   �   a��*[F��f��D�¾1%��e*��,��T>��AJ�H�N�tDK��8@���.��	�����UȾ�8�O��z�y��P󚼈�B<���<��<�r<pWh�� p�����TF��b��u�¾���)'�.,�Q>��=J�l�N��@K��5@���.����
���QȾ-���+�O��w����D뚼h�B<���<��<��r<(�h��.p��   �   0u:�X����Ⱦ}��%�PF�]-c��z�-|��,>��P���|�J�e��I���(����z�̾���
T?���۽ >���^����<"=���<x�L<�$���7��s���l�>�lM���#���Ծ;$�� �	����IE�ŷ�C`���h ھ쇳� Ջ�]K��i�J����#�0z�;4i�<���<��<@H}�d8�(=ս�   �   ����C������*�w�S��I{��*���������TL��ڒ������l����}�V�ߛ,�z�F��֎��^x�����h鮼z�<�=X�,=�_=�yo<@3��<@j��Fٽ��$�LD_��_���B�����K�Ⱦ�ξ{�ʾ����6���x��m��S3��w��� ��D������:��<"z=T��<��#<��ͼ����q��   �   �F���U��"���Q�`?�����<��(X��!�ǿQ�˿�kȿ7O��?��֝�����*!S��^#�{�ﾁ���\�N�| �:'��"�;(=:�O=Z�T=�`*=�į< ��da+��1�������&�L�-j��~���Ӏ��q�"=V��3�<X��4ǽ�q���Ƽ@А;��<b�=�=p<�<�h�\6C�����R��   �   )�ȾA\��(A��vw���������ɿFܿ��m����1�ܿ�rʿ�ز�# ����w�'�@�c��P�ƾ�IB���v� K��=N8g=b�=��=P=��=�� <<����J�����Hս  ��������=��[����vc��u���h��h�9��VH<�,�<!1=��@=��$=���<x-u�H��;������   �   zH��e$�\�A������ȿ����=���Q�X��N�V���Y��ȿ5��|�u�Z���"�M�依ᔾr -�o���pOM��H=8Bu=�
�=8X�=��=�Mz=��6=���<`͂;䷈���0JO���y��ӆ�Ǚ��n�m��=�85���W� ۳;���<Bw=rjN=�Be=<�[=D(=8P|< ^ܼ���7��@���   �   �� ���4��6q�%5���k��-ڿV��@^����$:� ��`|�m����ٿ<칿�q��Mo���2�6R�����t D�r���������<��|=���=���=�ɳ=��=�Ŏ=�c=�Z$=��<��/<�zD�0H���R�� P�����B���<�۳<`=�;@=�i=l�=�݃=gl=\x'=�/<:��ٽ@�P�6@���   �   ����?���~��z��G6Ŀ�u忈���O�X ����@�4L��b�A��Wÿ�_��,9|���<�3��ό����R�qϽD=ѼP��<V�=ߠ�=��=`��=p��=���=�*�=��y=j%G=~�=���<$��<p��<`��<�`�<|��<�z=<�,=�S=�w=.2�=R�=~��=v<u=�%=�a�;:�0���(�`��ж��   �   �b�-IC�z���S��`�ǿ#Y�����&��4I����ܦ�����迚�ƿP���S���b@��U��D����W���ս�"���<���=,�=�*�={��=�x�=^��=F�=��=�g=��;=V=��<�B�<���<���<�
=�&=@�G=j=-�=/�=�S�=�Ð=X�w=��$=���;��9��_���#f�pͺ��   �   -����?�`�~�$z��n5Ŀ�t����dO����������K�0b�O��JVÿ_��8|��<����֋��G�R�>oϽ88Ѽ���<��=:��=��=���=���=���=�*�=��y=t%G=t�=���<8��<���<���<0a�<���<({=��,=x�S=��w=s2�=sR�=�=�=u=j�%=r�;b�0���`��϶��   �   V� ��4�\4q��3��Nj��A+ڿT��]�����8�̾�@{�k���ٿ�깿�p���Jo��2��O��=�����C�ۦ��춦�l��<��|=���=(��=Fʳ=��=�Ŏ=&�c=�Z$=���<��/< |D�(H�8�R�P P�����B�h�<�ܳ<�`=�<@=.�i=��=�ރ=:il={'=x0<�4�?�ٽ~�P�F>���   �   �D辄c$��\�?��]��{�ȿޗ⿩:��P�����}�>����㿅�ȿ����t�Z�`�"�¡�ߔ��-�t���H4M�.M=BEu=��=�X�=!�=Nz=��6=̍�<�͂;������6JO���y��ӆ������m���=��3���W� �;࠿<�x=6lN=�De=*�[=�G(=�e|<�Nܼ�����7�#>���   �   ̴Ⱦ]Y�B%A�Grw�F��������ɿ�ܿ	�i����ܿCoʿ�ղ�}���O�w���@�����ƾ��~��=���v���J�B=�;g=��=�=��P=$�=�� <����J�����Hս  ��������=�o[�e��c������D����9��]H< 1�<�#1=*�@=��$=d��<h	u��A���������   �   B���O��"��Q�r<������{��T����ǿ�˿�gȿ.K��V;�������LS�
[#�^������N��߽�,'��i�;(.=>�O=�T=tb*=�Ư<Ѓ�,a+��1�������&�L�;j�	~���Ӏ��q�=V��3��W�4ǽ@q�ԳƼ��;t�<:�=�=�J�< ��j(C����&R��   �   j����=������*���S��B{��&������j����G���������$i����}�	V��,�$v�	��;����q�z��ή�T��< %=n�,=�b=�o<X1���?j�gFٽ��$�OD_��_���B�����R�Ⱦ�ξ{�ʾ�����5���x��Bm��S3�w���������� �:h�<j=���< $<diͼ$����j��   �   Pl:�w�����Ⱦdx�g�%��IF�&c��
z�x���9��&���	|��e��I�T�(�;����̾3�PK?�Ș۽�>���]�8��<(=���<h�L<�!��j7��9���b�>�mM���#���ԾE$���	����KE�Ʒ�@`�	��U ھ҇���ԋ��\K�!i�.��@��;\s�<��<���<�m|�(Q8�0ս�   �   d��PF��_��՚¾��~$�,��M>�7:J���N��<K��1@���.������ MȾ-�����O��r�����њ���B< �<�*�<��r<�Nh�:p�{���TF��b��x�¾���.'�5,�Q>��=J�q�N��@K��5@���.���o
���QȾ���ʧO�kw����p䚼��B<� �<�)�<�r<�:h�p��   �   2��ߋ��{�>�HJ�����;Ծ����	����A�s��]������پ���ы�4VK�d�~w�����Վ;}�<x��<D��<`�|��V8��4ս�o:�ĵ����Ⱦ`z���%�~LF�n)c�zz�z��<��I��|��e��I���(����Y�̾�����P?�i�۽�>��D^�l��<�&=���<мL<����   �   ����3j�N>ٽt�$��=_�\��X>�����"�Ⱦ(ξ�ʾW���1��et���	m�0M3��l������t����@�:�#�<<�= ��<�$<,oͼ�m�����?��m�Ż*��S��E{��(���������$J�������8k����}�~V�֙,��x��������u�]���lޮ���<D#=�,=�e=@�o<�   �   �ԯ<`6�dT+��)��������&�QL��j��~�����΀�pq�z5V��3�R�*ǽ �p���Ƽ�1�;��<,�=�=�L�<`��+C����;R��C���Q�n�"���Q��=��!���)���U����ǿ+�˿�iȿWM��h=��h������@S�|]#�E��磤��N�N�߽b5'� A�;�+=4�O=�T=�f*=�   �   ��P=t�=x<�k���
J�����>ս� �������r7�zU�Ey�Y��*���B��p�9���H<<@�<X)1=�@=��$=l��<u��B����\����ȾKZ��&A��sw�Q�������ɿ?ܿ��k� �迃�ܿ0qʿ�ײ����#�w���@�y���ƾV�A�j�v���J�t=6;g=*�=:�=�   �   ��=&Sz=��6= ��<`!�;\�������:O� �y�4ˆ� ���|�m��=������V��8�;���<�=�qN=Ie=2�[=�I(=j|<�Nܼ"�����7��>���E�&d$��\��?��(��v�ȿ��<���P�����~�����1��ȿp���󋿔�Z��"�v��ᔾ�-�{���PIM�J=
Du='�=�Y�=�   �   6˳=<�=Ȏ=l�c=a$=\��<�0<�B���8oR��O���
��Y@���<�<�g=�B@=
�i=��=��=�kl=�|'=H	0<�3��ٽx�P�^>��v� �B�4��4q�4���j���+ڿ�T���]����9�t���{�Yl��Z�ٿ�빿�q���Lo�{�2��Q������d D�s�������L��<�|=���=���=�   �   ���=��=l��=,�=`�y=�(G=��=���<��<�<,��<�k�<���<�=ޝ,=F�S=��w=�3�=�S�=���=�?u=N�%=���;6�0���� �`�8϶����ƞ?�:�~�z��z5Ŀ�t����O����P����L��b���Wÿ�_��Q9|��<�g��4���N�R�0rϽ�@Ѽ$��<��=���=��=�   �   ���=Ƈ�=��=�T�=�/S=�=4��<�<�&<0 �;0Z�;HGA<욜<P%�<`�#=��R=:;}=��=��=5��=�Lg=ܫ�< w:�&����-��ᙾ���2�c�w������̿����,��X�#��3��f=�0A�Nc=���2�:9#���?���=˿6?�� ut���/� ����"�����w�:.O7=���=��=�   �   �í=�L�=�p�=�0l=N�1=�7�<� �<��;��ֺ`���Q����:��<D��<�r=�6=��f=���=B��==$+c=��<�&��H��VW)��{����1�/�8Ss��$��Ksɿ���f.�x� �f�/�� :� �=��:��/�x� ����`S�
�ǿN���^4p�l�,�9��?琾���P�|���;�p6=��=#h�=�   �   E��=�%�=4Y=8=p9�< �t9l3����������+��4&�v��<c���� G�;и�<�� =�VU=�u=��y=
V=���< �ܻ���|�ʤ��,hྔ�%�pNf��ꗿ�i����翺/�����&��S0���3�x0��'�t����n��7g������C�c��5#�dz۾�����"�֭a� F�;�33=���=���=�   �   h�h=�V/=���< ~�$�м�/M�8���܃����н|۽�6ֽ��½����Des�f��P��f"<���<`Z1=�L=t?>=H��< .𺰫_����@�z�5ʾR�@�Q���������Կ���Y�T7���!�f�$�2�!�j��n���#����Կ�R���c���VP����bƾ��r�����V�8���<�+=Hq=���=�   �   ��<�5<謭���`�.4���G �vf ��/:��IK��R��N�L�?�)(���	�';Ͻ2l��n/	��������<R=��=�7�<��f;�U'�v�߽�YT�m.������8�&Eu�Ѯ��AL���hݿ����N�����x�`����F%��Tm޿�뽿替B
u��h7�.��̢���bN�j(ҽN���K<��=��E=L#8=�   �   ��n���5���u8�
)k�6g��.����Ū�q��&D��g���Mn����t��gC�QA�I\��BxM�@�v�8�'<ܥ�<|�<`r<�%׼���b�)��̎�w�پ+���
P��ℿkY���|���V׿������/�������E\�E�ؿ�迿�q������Z�P��`QپI�����%�����`���/x<Dd=�s=e�<�   �   ��K�J�̽��#���h�����s����۾.~�����L����޷���e�%K���7���t���.�����~q�8��i�;HL�<x�2<�*K��{e�)����	]�ˮ��4I���-)���Y�1��������)����ÿ��οe�ҿ+�Ͽ?ſ�ʴ�Ǖ��]��z \��*�����hl��r]�����J![� ����<��<��P<��@��   �   ]�ٽj%4��W��(t����侔q
� �a21��p<�o�@��p=�N3��|"��?��~��츾�U����<�.�Kn�s��0x�;0?3< �������ӧ�������*����H���*��T�'�{��\��=��JC��{�������"|��m됿��~� W�^q-��1��U��|ꂾ 0!�¸�� G��@��:`ra<�W<��Y��BT��   �   �P2�
ӈ�����TA��� ���?���[���q�81��2悿+ɀ��t��g^���B�t#�/F�
xžx��`%8��{ս�E��_4�K�;P�<���S8���̽�J2�6ψ�����d;�� ���?�=�[��q��.���タ�ƀ�Gt��c^�^�B�� #��C��tž�|���!8��vս�E�PX4��@�;��<���B_8�V�̽�   �   $������lK�K�*��T���{�	_���?���E�����V���m~��}퐿��~�!W��s-�p3��X��p삾�2!�Ļ��L��@��:H�a<�r<�XY�4T���ٽ 4��S��,o����3n
�T��h.1��l<�Y�@�m=��3�Vy"��<�+z��踾�R����<��'�Cn��j�� ��;�63< ����ڧ�����   �   r����M���0)�@�Y�F ������,����ÿD�ο�ҿ��Ͽ^Aſ�̴������^���\��*�����dn��]�����$[������<護<ȬP<�@���K��̽�#�z�h��������}�۾�w��r�HI�b��ӱ��6`�pF���3��mt�ȸ.�C���tq�x�� ��;XL�<��2<�CK�H�e�Ι��@]��   �   F�پ����P�z䄿�[���~��Y׿T�y���Ք��2����^�J�ؿ�꿿s��Ǘ��#�P�p�7Sپ}���d�%�d���<a��8x<�h=�z=�w�<P����]�h榽���Ln8�� k��b��)��������k�� ?������j��_�t�qaC�\<��T���lM���v��'<���<��<�c<�3׼����j�)�pώ��   �   ���b8�Hu�����@N��!kݿ����P����z������'���n޿�콿盿�u��i7����ã���cN�e)ҽH���K<.�=��E=�*8=��<�g<�����`�=)���A ��_ ��(:�RBK�<R�.N�f�?��(�I�	�2Ͻ�d���#	��@��h��<�=p�=�4�<��f;$]'���߽�]T�;1���   �   �S�s�Q�\��/����Կܼ�� Z�r8���!�z�$�.�!�F��&���$����Կ�S��\d��NWP�`��Tcƾ9�r�������8���< �+=LLq=���=��h= `/=İ�< �޹P�м4M������y���н�۽�,ֽ�½R���JVs�dY��O�p�"<H��<(^1=�L=r?>=<��<��𺰲_�6���z��7ʾ�   �   �%�HPf��뗿)k����翂0�����&��T0���3��x0�x'�������濑g��ﻖ���c�6#�yz۾x����"�H�a�V�;b63=+��=���=ɳ�=)�=��Y=�=dM�< �9������^�+�(&����N���� ��;8��<T!=ZU=�u=P�y=PV=D��<�ݻ+��`~�q���mj��   �   O�/��Ts�_%��0tɿ����.�� ���/�:���=�	:�D�/��� ����lS��ǿ7��� 4p�)�,�����搾�����|���;�r6=��=~i�=�ŭ=�N�=�r�=p5l=��1=hC�<��<��;��պ}��0!�� :8�<h��<Jv=��6=T�f=���=o��=���=�)c=0�<h�&��K��:Y)�9}��>���   �   Q�2�3�w�����r�̿���d����#��3��f=�2A�<c=���2�
9#����>��k=˿�>��4tt��/�������"�������:pQ7=���=t�=X��=T��=G �=$U�=`0S=֗=`��<��<�&<  �;`X�;�EA<���<�#�<t�#=��R=*:}=j��=��=r��=�Jg= ��<(�:�*���t�-��♾7���   �   t�/�uSs��$��Rsɿ���P.�N� �&�/�< :���=�H:���/��� ���mR�-�ǿ����3p�U�,�����吾�����|�`;@t6=>�=�i�=�ŭ=�N�=�r�=z5l=��1=PC�<��<�; �պ0}��!�� :��<���<xv=��6=��f=���=���=)=�*c=X�<h�&��I��X)�X|������   �   i�%�"Nf��ꗿ�i�����\/����6�&�S0��3�:w0�'�����
����e������z�c��4#�.x۾ު��_ �h�a� u�;�83=���=��=��=?)�=��Y=�=HM�< �9P������n�+�(&�����M�� �����;8��<�!=�ZU=�u=Όy=nV=��<��ܻ��|�Ĥ��h��   �   �Q�x�Q�y
��ⵯ���Կ����XX�x6���!�V�$��!�T��f���!��D�ԿqQ���b��lTP�/��&`ƾȚr������8�`�<��+=�Nq=O��=r�h=v`/=$��< �޹T�мRM������y���н�۽�,ֽ�½7����Us��X���O�؉"<���<�_1=�L=^B>=|��< ����_���h�z�b4ʾ�   �   ���8��Cu�ϭ���J��cgݿP����M�`���w� �^���"��(k޿�齿Z䛿Zu��f7�S�������^N� "ҽ~z��7K<r�=��E=h,8=��<�i<�����`�H)���A ��_ ��(:�fBK�HR�6N�f�?��(�2�	��1Ͻvd���"	�p6�����<=�=�>�< �f;�R'�f�߽hXT�V-���   �   ��پ����P�yᄿ�W���z���T׿k�N�����������Y���ؿ�濿�o��є��R�P����Mپe�����%�z퟽�K���Tx<Fm=�}=�{�<���$]�K榽���Sn8�� k��b��3��������k��%?������j��H�t�LaC�*<�T��tkM��v���'<L��<��<��<�׼_���|�)�?ˎ��   �   ����FF���+)�)�Y���������|'����ÿ�ο��ҿ�Ͽa<ſUȴ�t���[����[�!�*�����h����\�����[�X��d.�<p��<��P<ȍ@���K��̽�#�|�h� �������۾�w��y�MI�f��ֱ��3`�dF���3��>t���.�����rq�����;hW�<8�2<�K��ue�����]��   �   ���I����F���*��T���{��Z���:���@��򚩿L򦿚y��鐿��~�/�V�n-��.�]Q��炾�*!�����D-��@�:p�a<��<8MY�P2T��ٽ�4��S��0o����9n
�[��p.1��l<�`�@�m=��3�Vy"��<�z��踾�R��/�<��&齊@n�4c�����;pU3< <� ����ϧ�����   �   �F2��̈�_����6��U	 �L�?�~�[���q��,���Ⴟ�Ā��t�p_^�a�B�'�"��@��ož�x���8�rmս��D�P'4����;8<8���P8��̽�J2�,ψ�����i;�� ���?�G�[�!�q��.���タ�ƀ�Lt��c^�\�B�� #��C�{tž�|��d!8��uս,E��D4�@y�;P�< ���J8��̽�   �   ��ٽ]4��P��Lk��?��_k
����*1��h<�L�@��h=��3��u"�~9�2t��㸾�N����<�`齈2n��O��@ۚ;0a3< =�h����ҧ�S�����$����H���*��T�.�{��\�� =��PC����������$|��n됿��~� W�Wq-��1��U��Pꂾ�/!�R����>�� k�:`�a<@�<�9Y��)T��   �   6�K�-x̽�#��h����T��"�۾�q��@��E���X��� Z��@��/��5t��.�P��Bcq�4� �;Ha�<3<�K��xe�I����	]�����/I���-)���Y�3��������)����ÿ��οk�ҿ/�Ͽ?ſ�ʴ�ƕ��]��s \��*�����El��]�M����[�8���)�<Ը�<��P<�q@��   �   �D��dQ�wަ����0h8�Yk�_^�����������f���9������^e����t��YC��5��I��^[M���v�H�'<ؽ�<l�<x�<$׼�����)��̎�o�پ+���
P��ℿoY���|���V׿������4�������H\�G�ؿ�迿�q������T�P��FQپ �����%��򟽐X��pHx<m=:�=��<�   �   ��<،<v��2�`�, ��E< �nY ��!:�;K��R���M�y?���'���	��&Ͻ-[���	��Ԍ��Ø<#=ҵ=�D�< g;S'���߽�YT�`.������8�'Eu�Ӯ��CL���hݿ$����N�����x�b����G%��Um޿�뽿替>
u��h7�%������pbN�Z'ҽ���)K<x�=�E=08=�   �   ��h=�f/=���< �ٹ �мLM�쓽7p����нv۽1"ֽ��½��~Ds��I���O���"<h��<�f1=L=0F>=���<��ﺦ�_�H���z�5ʾR�@�Q���������Կ���Y�T7���!�h�$�2�!�j��n���#����Կ�R���c���VP�݅��bƾf�r�����8�p�<��+=�Nq=q��=�   �   5��=+�=��Y=T =�\�< ��9���l�����N�+��&����h5��X�����;X��<B
!=�`U=��u=��y=v V=� �<�ܻS���{�����(hྒྷ�%�qNf��ꗿ�i����翼/�����&��S0���3�x0��'�t����p��5g������A�c��5#�Wz۾r����"�`�a�pW�;73=���=���=�   �   �ŭ=bO�=�s�=*8l=�1=�K�<��< @�;�պ�J���툻��:�<4��<�{=~�6=��f=y��=5��=yÉ=<-c=��<�{&��H��CW)��{��|��1�/�:Ss��$��Ksɿ���f.�x� �f�/�� :�"�=��:��/�x� ����`S�
�ǿN���^4p�j�,�3��5琾�����|�`�;r6=��=�i�=�   �   ��=h�=a�=X�M=��=���<P#�; �x��5���g���Q�@��@L;�sj<��<*�,=��`=���=
t�=%݂=��F=x��<���ϱ�B�c��¾�+��p[��x���mĿ�����y��.�^F��Z��xh�Drm�sh�aZ�,�E�nD-���J��R¿����-X�#@�fh���nZ�BϽܶü�J�<k=�`�=�   �   (�=A�=��h=zo,=���<��<0O��ߋ�ģ̼��ۼ�̧��L&���U;�e�<8|=��E=��q=���=\p{=��A=�E�<|N���ڽl^��v��4<��gW�ԓ�b��'����~�*��xB��VV�j�c�@�h���c�HJV��.B�2a*��%�C�￑-��K
��:T�)u�Î���vU�0eɽT;����<�Le=� �=�   �   ��{=�LU=��=�M�<��v�P�ȼ$�0���m��Y��l���g���q|��NE��+��85�`�<��<H�1=��W=��[=�1=,ȑ<<a߼�ȽP8O�����4���K��%���l�������
��F"��$8�wJ���V�Tf[�dW���J�X88��"��M
�������}���xI��V	��d��`G�	������H{�<�+S==�   �   ��'=T9�< ��:��Լ:b���f��ě�4��"���
�	���Ap���r��hi��4㻈�<�=�$=:*=�@�<��7���L�7��������d9��!��I��Wӿ�J���	���(��8�дC�ڳG�JD��\9��)��M�dC����ҿ����q~�x�7��J�����1��8��pSt���<ȸ2=~�E=�   �   �q1<4���.�N������_���1��oW�\�u��ㄾ����^���1z�΅]�j�8��s�B�ɽF�p�(-ż��F;0~�<�N�<�a`<,@���e���������po۾�/"�7�a� ����ͻ�4E� ��b��p�#���,�nJ0��X-�0d$����@G���q��8ה���`��#!��پ�"��nm�j,����%��|�<�� =��<�   �   ����O푽�m��D7�v�t�禘��γ�o�ɾm�׾-ݾ+پ"̾�V��Ɯ���}��@��3�}ڡ��M�����<X�<6��U��l��(k`��`�P?��~�[	����ÿn�俢� ����z��]� �������k�7�Ŀ�ۡ�i�~�&?�t��Tϴ��e]��,��+E� �һ@X<�#g<�V���   �   �[�����8a\��w����¾�"�_�	�Q����"�IY&��~#��R�İ���񾹲Ǿs'��T�d��_�����L�4��>h���� �	�����-���y,�Df��bھ����	P��ᄿGW���w��SO׿��꿱���S���J���д�9Uٿ�h��^�����Q�G����ھ�a���d+��P���%
�p]�� j;P(����   �   �*��jo�6b���⾬��Ɨ+�L3E�*�Y�&�f���k�s�g�6�[�P�G�kn.�Q��3��୮�K�v�����Z����0����(3�����F�r�������T�᥾L����"�D@R��m��Ǽ��T������Y/ȿK"̿�ɿc���,��T������y�T�[�$��^�Ǌ��g�V��Z��ҫq�x���pj绨UY���!�� ���   �   �l�7�����򾅲��RE��j��ޅ�1������X����0��9��[r����m��hH��S!�������/gq�E��K�����@�[�p�T��
�����(�l�����������NE�f�j�܅�y���/}������#.���6��p����m�}eH�?Q!����칲��bq�i��
����@�[���T�0�
�������   �   z奾����"�>DR�Hp��^����V������e2ȿP%̿xɿ��/��q���b��_�T���$�b�'�����V�|^���q�����K��6Y���!�%����$��bo�X]����&����+��.E�r�Y�J�f���k���g�Պ[�[�G��j.�m�����C����v� ���U��,�0���0<�̻��r����~�T��   �   �ھ���bP��ㄿ�Y���z��JR׿�����}���O�����쿴Wٿk��+�a��a�Q�����ھ$c��nf+��R��(&
�0F�� �;h�<��vR�����fY\��r���¾���	�q����"�HU&�{#��N����&����Ǿ�#��f�d�.[�Н��|�4��.h� ��
�����3��n~,�yi���   �   ��@?�i~���+�ÿ/��  �����|�D_���x�� ���m���Ŀ�ܡ���~��'?�����д��g]�u.�:,E� �һ�SX<�Bg<@��������㑽na���<7���t�ڡ��	ɳ�j�ɾ2�׾�&ݾ�$پp̾�Q������=�}��@�U/��ӡ�PD� ���0<�}<X!6��U�;s���o`����   �   02"��a�����л��G�r��Ը���#��,��K0�rZ-�ze$����(H�:俘��ؔ���`��$!��پa#��n�,��8�%����<�� = ��<h�1<��� �N�����&Y�21��gW���u�X߄�
�������)z�R~]���8�-n�_�ɽp�p��ż@RG;<��<\Q�<�[`<hI���i��ٹ�����r۾�   �   �f9��"���J���Xӿ�L���
�0�(�z�8�D�C�B�G��D��]9�l )��N�{D����ҿ�����r~��7�QK��X��^1�C8��Lt�4"�<��2=��E=2�'=lN�<@=�:d�Լ�'b��髽�཮��������X|	����Hg��Ok��(]�p��x�<��=t�$=n*=t<�<���F���f�7�S���7����   �   ��K�'���m��6����
��G"�&8�(xJ���V�jg[�XW�f�J��88� "�>N
���L��������I��V	��d��G�C��`������<2/S=�=|�{=TU=z�=�a�<��u�zȼ̝0���m��Q����������c|�&BE�����5�H<��<T�1=B�W=��[=�1=0Ñ<�j߼��Ƚ;O���������   �   �hW��ԓ�S��8����$�*��yB�xWV��c�ظh�t�c��JV� /B�La*��%�5��w-��'
���9T��t�=����uU��cɽ�5��x��<�Oe=0�=�)�=C�=T�h=�t,=���<h�<���Ћ���̼(���ۼ�����5&���U;�m�<T=$�E=�q=Ӳ�=�o{=�A=H@�<�V��#�ڽLn^�x��>=��   �   tq[�y��fnĿF���z��.��F��Z��xh�Drm��rh��`Z��E�(D-�ԁ����<R¿0���^X�{?�^g��BmZ��Ͻ �ü�O�<k=Ya�=��=�=��=Z�M=��=8��<�(�;��x��5�x�g���Q� ��`A;@pj<��<�,=j�`=��=Os�=M܂=��F=��<��-��شc��¾b,��   �   �gW�Aԓ�}��1��x��b�*��xB�jVV���c���h�R�c��IV�>.B��`*�%�;�￪,���	���8T�%t�;���<tU��aɽ 1�����<�Pe=w�=�)�=0C�=r�h=�t,=���<H�<���<Ћ���̼@���ۼ�����5&�`�U;�m�<|=p�E=x�q=��=�p{=:�A=�C�<�Q��:�ڽ�l^�w��<��   �   ��K��%��<l��A�忢�
�HF"�V$8�<vJ���V�Be[�DW���J�R78��"�M
�������n����I��U	��b���G����@�����<1S=�=&�{=vTU=��=b�<��u�Lzȼ��0���m�	R����������c|�&BE����5��<x�<�1=@�W=J�[=1=�ɑ<�`߼,�Ƚ[8O�����!���   �   +d9�&!��_H��<Vӿ�I������(���8���C�x�G��D� [9�>)��L�[A����ҿ����^o~�t�7��G�������0�x3���2t�l*�<�2=l�E=�'=hO�<�B�:h�Լ�'b��髽'�ཿ����������_|	����4g��'k���\�`��T�<��=��$=r-=lE�<l��C�����7�����M����   �    /"�ާa�7����̻��C�6��J��(�#��,��H0�lW-��b$����E�y	�o���Ք���`��!!�9پ8 ���i��&���%�\��<�� =���<��1<���ֲN�����3Y�H1��gW���u�e߄��������)z�S~]���8�n�#�ɽ��p��ż�kG;,��<�X�< q`<T9���c��e��֥��'n۾�   �   4��?��	~�����ÿe��p� �����y�\�������p��
i���Ŀ}١���~�*#?�0���˴��`]�#%E�@tһ�hX< Pg<��������f㑽Wa���<7���t�硘�ɳ�|�ɾA�׾�&ݾ%پw̾�Q������(�}��@�#/�ӡ��B� ���,<�<x�5� �U��i���h`���   �   �ھ8���P�3���{U���u���L׿3�꿸���2���������CRٿ3f����	����Q�o��5�ھ;^���_+�WI��t
� ���#;���6���Q�����`Y\��r���¾$�ʌ	�{�� �"�OU&�	{#��N����"���Ǿ�#��4�d��Z�񜸽Ҙ4� h�@#亘�	����K*��hw,�|d���   �   �ޥ�ܻﾊ�"�`=R�5l�������Q������,ȿQ̿�ɿl���)������G��}�T��$�rY򾶆��7�V�eQ����q�0���`
�"Y���!�2���|$��bo�X]����+��Ɠ+��.E�}�Y�V�f���k���g�܊[�^�G��j.�j��z��-�����v����|T��f�0�����������r������T��   �   ��l�|�����R��zKE���j��م�����z��ԧ��^+���3���m����m�PaH��M!����D����[q����m����X�[��T�<�
��𜽒����l������� ���NE�o�j�܅����6}������&.���6��p����m�{eH�9Q!����й��vbq����P����� �[�p�T�Z�
�휽����   �   � �r]o��Y��s��M��`�+� +E�(�Y���f��k���g� �[���G��f.�ݨ�}��P���	~v����L��ܨ0� ���������8�r�����Z�T�l᥾F����"�H@R��m��˼��T������a/ȿP"̿�ɿg���,��S������t�T�R�$��^򾡊���V�VY��J�q�Ԟ�� 绨Y��!�(��   �   �K��.��pS\�o��c�¾���	���(�"�RQ&�	w#�K�ߩ����2�Ǿ���b�d��T�����(�4�h�g� h���	�J��G,��my,�%f��Uھ����	P��ᄿJW��x��XO׿��꿷���Y���O���Դ�<Uٿ�h��^�����Q�>��|�ھ[a���c+�O��B 
���� 0;������   �   (���uܑ�X���67�`�t�����ĳ��{ɾA�׾� ݾ�پo̾4L������S�}�H@�)�jɡ��3��E���I<��<x�5���U�}k���j`�j�]�Q?��~�]	����ÿq�俣� ���{��]�$�������k�6�Ŀ�ۡ�g�~�&?�i��/ϴ�be]�L+�@'E�P�һ�gX<�[g<���   �   h�1<Ln����N�ݥ���S��x1�``W�f�u��ڄ�����d��� z�v]�d�8��g��ɽ��p���ļ@H;؛�<Xd�<�`<�5���c��������fo۾�/"�:�a�#����ͻ�6E� ��d��r�#���,�pJ0�Y-�2d$����@G���q��6ה���`��#!�xپ�"���l��*����%���<v� =d�<�   �   ��'=�]�<�v�:�kԼ�b��૽�������~����Dv	�V���\��	b��M��{�T�<(�=ȗ$=
2=�K�<�
�������7���������d9��!��I��Wӿ�J���	���(��8�дC�ܳG�LD��\9��)��M�eC����ҿ����q~�r�7��J������ 1�S7���Dt��&�<��2=�E=�   �   ��{=�XU=z�= q�< Pu�LdȼV�0���m��J��ᓓ���~T|��3E�8���@�4�C<��<�1=��W=��[=�1=8ϑ<�\߼[�Ƚ8O�����2���K��%���l�������
��F"��$8�wJ���V�Tf[�dW���J�Z88��"��M
�������{���tI��V	��d��$G�V������\��<�0S=�	=�   �   E*�=�C�=��h=x,=���<�<`諻DË���̼\����ڼ�����&��EV;�y�<�=$�E=��q=մ�=�s{=��A=I�<,L����ڽ�k^��v��3<��gW�ԓ�c��)����~�*��xB��VV�j�c�@�h���c�HJV��.B�2a*��%�C�￑-��K
��:T�'u�����bvU��dɽ�8�����<LOe=S�=�   �   �M�=�$�=�S=@�=�ߤ<@rh; s:���Н��������HBҼ�p��{�8n}<2=��==j=�;|=~�h=r� =@��;��[��S��������M33��݀��p��1���j�Ш,�  L�ܩj�����ˋ�����Ƌ�����.j��K� |+��*��῍_���G~�fc0�6�B,����x�C��!#<�7=��~=�   �   �_�=�5h=��4=�<��<����1м����,A��&O�@]F�H�'����p�W��Ò;A�<�=��Q=�tj=��\=�a=��; �U����0�������/��}��m�����|�)��3H�|�e������%��#Ɉ� ��|�e�*wG�ƥ(���
���ݿ%���5�y��&-��ྰD���[�R>�@Q <Ɯ0=��r=�   �    J=V�=؂�< �,� �Ǽ$�C�#錽�I����Ž�νm�Ƚ�����]����U���@z»��<�9=\4=�58=�=�y;�D�4���5���]׾�&�~�o�Ȭ���տ�$�Z!��o=�p�X��Ip��=��w0��^����p�4�X�H/=��{ �Vf�	pӿC*���m���#���Ӿm�y�����6e.�X1<@�=��M=�   �   t��<PF�;�ҙ� �L�����j����--��<���B��>�&0�$:�R��������c�$�Ǽ`k;�J�<�
�<�k�<@];��+����e��W¾ܹ�L�Z������ÿ���
��P-��EE�"�Y�&�g���l��h�jLZ�t�E�j�-�����f��N�¿!���X�c�>E���_�g�������;���<�g=�   �   �P��<��~W���0��`��	���q��;آ�9 ��;٣��Q��n����lf�\[6����n$����4�`EW��"�;��8<@ꪺ�R���Ž.D���0g��@�7}��Yŭ�aڿ��� ��F.��?��J���N��#K��@�z/�\�����Oڿ���a���?�bM��¥���?�tk��.{ ��B;�C�<��5<�   �   �`��н��#���g�w`���>���پ��<r��|�T������ܾ�Խ���ɛn��r*�hKܽ�t���Ҽ������0��� ���H�����N~۾4�!��Ka�ݾ���������jm��}�<[#���,��0��@-�vi$�֩��t�o�#l��I'���na���!�[wھ�K��vm�,v��طۼp�����s�D����   �   �<�5=��1�����&뾹�k�#��Q5�9�@�(�D�ۄA�u�6�O�%��D�u�ﾀ������v,C��.���Ҋ� }	�$���$n߼ܞs����hGY��������7���t�Zv������ݿ������.��t]��#��	�V���?߿ƾ�����Prv���8����﮾yaX�{���k��*̼hp��0`��ꌂ��   �   RZE����f�ξ:�.*�*/K�j�h�S���u��0C�������+k�~�M�5�,�so
���Ҿ�����I����#e�������ī5�9���:Y ��2��y;ɾCk�s3A�@�w��������l�ɿ�ܿs%�N����i�ݿ��˿���7F���0z�=C����˷ʾ:���t� �`K���^2��ۼ������]���   �   �C��ȞԾWT�0X<��h�G���G�������`1���ʸ���|٬��C���n��I�k���>��L�3~׾�F���=��0޽2 o��	��U��;k���ڽE�:��?����Ծ�P�T<�U�h�����Y����~��3.���Ǹ���֬�(A���l��y�k���>�aJ��z׾)D����=�"-޽:o�`�	��[�ZFk�ҹڽ�:��   �   @ɾEn�<7A�͉w�+��������ɿ�ܿ�(�ū�E�}�ݿq�˿K��@H���3z��C������ʾ����� �JM��`^2���ۼ.�����{�SE�f����ξ��**��*K�V�h���� s��k@��9��y쀿P'k���M���,��l
���Ҿ�����I�d���b����d缸�5�W����] �6���   �   ����7���t��x��|
��ݿ(���V���L_��%��	�1����A߿Ⱦ������tv���8�`�f񮾶cX�� ��k��$̼�b��0J�����2��-=�E-��|���A ���?�#�mM5���@���D�e�A�H�6���%�=A��������X'C��'��Ί�Px	����8u߼��s�����LY������   �   ��!��Na�����������o�r� ]#���,��0��B-�k$�<���u�q俰m���(���pa�
�!�yھ�L��wn�~v����ۼ Е� #s�\歼`�ޕн��#�,g�a[���8��p�پ��n�0y���,����ܾ�Ͻ��
��Ӕn��m*�kCܽ��t�ԠҼ�������<��������K�F���0�۾�   �   =@��~��Tǭ��	ڿ�����!.��?��J���N�Z%K�b@�� /�j��V�>Qڿ��� ���?�N��å�G�?��k��(y � HB;TQ�<H�5<P���������J��*0�V`���dl���Ң����ԣ�M�����Eef�U6����p����4��$W��H�; �8<���X���Ž�D�[�i��   �   ��Z�e�����ÿ'���D���Q-�.GE��Y��g�X�l�Hh��MZ���E�D�-�V���g���¿�����X����E��g�_�#���
����;��<�n=D��<��;촙�@�L����������(
-���<�<�B��x>��0�14�����F�����c��Ǽ �;�U�<x�<Xl�<�8;�+�a�꽓�e�@Z¾����   �   ~�o����	տ�%�^!��p=���X�Kp��>��.1���^����p���X��/=�P| ��f�[pӿt*���m���#�ՃӾ"�y�����b.�><N�=�M=lJ=P�=��< *�X�Ǽ�C�����A����Ž	�ν��Ƚ�����V���U��s�@5»8-�<R>=N	4=�68== �x;0�D�N��*7�� `׾f&��   �   :}��n��"�r�2�)�R4H�b�e����0È����rɈ�n����e�JwG�Υ(���
���ݿ������y�1&-�}��,D���Z�:>� ] <�0="�r=�a�=*:h=(�4=8'�<p�< ��$!м���#A�PO�UF�Н'������W���;dH�<t=��Q=Buj=N�\=B`=���;��U����v������'�/��   �   ހ�hq�����4k�&�,�V L�.�j�����ˋ�����Ƌ�r����j�LK��{+�x*�n��_���F~��b0��^+��ͯ���C�@-#<F7=��~=�N�=S%�=*�S=f�=��<��h;p:� ��<���������LCҼ��p�����i}<�=F�==�j=,:|=��h=$� =���;��[��T�������43��   �   }�n��.���p�)�^3H�6�e�Z��n�����Ȉ�����e�bvG��(��
���ݿB�����y�]%-�Q��dC���Y��>�d <�0=��r=b�=Z:h=0�4=H'�<8�<P��l!м:���#A�pO�(UF���'���뼰�W�0�;�H�<�=��Q=�uj=�\=va=��;ܿU�����������K�/��   �   E�o�����4տ~$��
!� o=���X��Hp�.=���/��Q]��0�p���X� .=��z ��e��nӿ)���m��#���Ӿ!�y�����].�@K<f�=J�M=&J=��=`��<�*���ǼF�C�ጽ.A����Ž%�νֱȽ�����V���U�ts�3»�-�<�>=<
4=n88=j=�'y;̅D�@���5���]׾�&��   �   ��Z�f���V�ÿ���^��6O-�lDE���Y���g���l�� h��JZ���E��-�����d����¿� ����X�� ��B��>�_������@��;���<�p=0��< ��;����F�L����������=
-���<�Q�B��x>��0�:4�����3���2�c��Ǽ��;xX�<��<�r�<��;��+����I~e�W¾g���   �   �@�s|��Oĭ�ڿ�������.�^?�B�J���N��!K��@��/�Ԇ�,��Mڿ(������?�tK�����U�?�e���p ���B;4X�<@�5<���������J��80�r`�#��vl�� Ӣ����"ԣ�M�����Gef��T6�t��)����4��W�p\�;0�8<@b��:O��Ž�D��茶rf��   �   ��!��Ia�����������>l�J|��Y#��,��0��>-��g$����r�Il俸i��A%��~ka�$�!�jsھ�H��i�]o��x�ۼ0�����r��᭼�`���н��#�2g�l[���8����پ3��n�9y���8���#�ܾ�Ͻ��
����n�cm*��Bܽ,�t���Ҽpo������{��0���6F�@���n|۾�   �   �����7�:�t��t������ݿ�~����r���[�"�(	������;߿Bþ�����Env�T�8�p��뮾�[X���񽪳k��̼�V���B��탂�z1��-=�C-������L ���H�#�xM5���@���D�m�A�O�6���%�<A��������'C��&���̊�t	�|���a߼6�s������DY����   �   �8ɾGi��0A��w����������ɿ�ܿ0"���~��ݿt�˿����C��,z�sC�����ʾ����� �C���P2�`�ۼd��L ���z�bSE�Z����ξ��**��*K�a�h����&s��p@��>��~쀿U'k���M���,��l
���Ҿ���"�I����`������缔�5�௰�MV ��0���   �   �<��ڕԾ�N�Q<���h�c���Փ���{��4+���ĸ��뵿�Ӭ�:>���i����k�{�>�G�:u׾@��;�=�i#޽�o�v�	��M��6k�+�ڽ��:��?��y�ԾQ�%T<�^�h�����_����~��9.���Ǹ���֬�+A���l��y�k���>�YJ�z׾�C����=�W+޽�o�Ǝ	��N�`3k�'�ڽl�:��   �   �NE�:
����ξ��&*��&K��h���}p���=��w���逿8"k���M���,�Bi
�
�ҾT
��|�I�|���aY�������漐�5������X ��2��f;ɾ?k�u3A�G�w��������s�ɿ�ܿz%�V����n�ݿ��˿���5F���0z�9C������ʾ������ ��H��:W2���ۼL�������t��   �   ?*�(=��)������뾺 ���#�VI5�9�@���D��{A���6�Y�%�m=�F��h��x����C�,���Ċ�Ti	��n���[߼ܘs�-����FY��������7���t�\v������ݿŁ����2��v]��#��	�X���?߿ƾ�����Lrv���8���Z﮾�`X�t��t�k�,̼�T���8��H���   �   �`���нF�#�Nxg�)W���3����پ���2k��u�B�>�����ܾ�ɽ�����n�`f*��7ܽX�t���ҼP+����Lw������JG�V���7~۾2�!��Ka�ྔ��������lm��}�>[#�Ğ,��0��@-�xi$�֩��t�o�!l��I'���na���!�8wھ�K���l��s��ܨۼТ��`�r��ӭ��   �   ���(�������@���0��w`�� ���g���͢�����Σ��G��T����\f�nM6������R�4�8�V�Ш�;�8<@۩�DM�#�Ž�D�w�*g��@�:}��Zŭ�cڿ��� ��H.��?��J���N��#K��@�z/�Z�����Oڿ���_���?�VM��¥���?��i��^u � �B;�[�<8�5<�   �   $��<���;����"�L�����^�����-���<��B��q>��0��-���������N�c�d�Ǽ��;k�<�"�<}�<��;��+�}�꽤~e��W¾ڹ�M�Z������ÿ�����P-��EE�$�Y�(�g���l��h�lLZ�r�E�j�-�����f��N�¿ �� �X�]�#E����_�����`��;���<�s=�   �   6 J=x�=���<��'�\�Ǽ��C��ٌ�'9���Ž)�νШȽ����\N����U��X�0���dA�<�F=�4=�=8=t=�Zy;f�D�̸�x5���]׾�&��o�Ǭ���տ�$�Z!��o=�n�X��Ip��=��w0��^����p�4�X�H/=��{ �Vf�	pӿB*���m��#�΃Ӿ/�y�"����b.�0A<Ҋ=��M=�   �   fb�=�;h=��4=�.�<�<��4м̵��A��O�zLF�6�'����W�� �;�T�<�$=nR=�yj=��\=�d=�$�;��U����$�������/��}��m�����~�)��3H�|�e������$��#Ɉ���~�e�*wG�ƥ(���
���ݿ%���4�y��&-��ྡD��j[�>��X <��0=v�r=�   �   T+o=H[=�D*=$4�<P-�;��4�D�߼f�$��eG�P�T�*�J��e+�H��xa�@�;�-�<��=ڬM=Ʋa=��K= ��<�������
50�Lᢾy���}K�0Z����Ŀ�����d�B���h��*��t���������y�������ۆ�؏g�"�A�`f�����$�¿ď�� I�����ԟ��C+��S���Q��Lh
=ІY=�   �   ��[=�@=rl=��w<P���܊̼��/�L�i�z	���>���߉���p�b9�c� ��P�B<X��<�3=jN="�>="�<����S���N,�&���;���G��̎�E����������K?�:�c�fE���>��{1��>��b8��4��P���&c�@?>�������������O��v`E�a�n�����'��"�������o=�\L=�   �   @�=(�<�"<�����#-�O��U���FN�E���o�� ��Y8�����񣑽��:�Pu�����;D(�<j�=�x=L2�<x���އ�F!�5���X��f�<��a���淿s��%�~85�j�V��Ex�����X���|S��Ք�4Պ��]x�b�V�l�4��d���x��P)���:����������4������t*�< �#=�   �   HK]<@�껆�����E�ܽ�����4�c�O���`��ag�8b��Q�7)8��O�D��\��t�#�P0���%<�ܟ<xQe<�-��t��$�����w�߾N�+�ߋw�,Ǩ�mvۿ:&	�:&���C��t`��Ry�]A���l�������z��a��D�^&���3�ڿ৿�u��U*��Sݾ'���ZZ�"�f����`�<�@�<�   �   �Ƽ hn�PGѽ:����S�:ۄ�C��Ox��V�������뽾����'��N-��]~X��>!���ٽD~�@b� �ʻ 2��p���W�(���,h� m¾�P���Y�+y��\(ÿ	?��d��8�,�4�D���X���f�Dl�X|g��Y�^�E��-����5����ÿ����Y�4]�����_�d����K���A�@�;��F��   �   ���:���:F��鈾����T�׾K����>��L�b��}��1F�oZ����ھV��������(K�R��֢���*�|���L.����?��˽aB?�����SR����8��V����pҿ>��$l���'��7�H�B���F���C�D9��)��t������Nӿ駿b)��I8�/s������Q=�[ǽ�:6��]��ܦ��@h��   �   �Z�"Vb��ᠾu־.H��"���:�\DN���Z��e_���[�f�O�s�<�φ$��(	�1�پ쵣���f��
�wo��"BO�q�83�!���X��<��ڔʾ���Q�Jt��q��o)Կ ���0��j���!�P9$�X�!�D�����y���M�տ�-��9*��l�Q�5�K�ʾN���9��O��\�,�
��n�E�,����   �   )k�7������B���f�פ���~���ј��ޛ��Y���s��m؄�Bi��^D�u���c��J�n�}�5D����[��8��
��v��\A��Ϛ�6辞$���[��x���5ȿ�͑��\���{��w��8��m��ʿY���.���@]�w%��x�r��pA����`���;4��V�Rj������   �   �ª�&��T=&��:V�cʃ��o��jK��}����e˿�RϿ�̿^¿Lݱ����(5����X���'�s���g��jKa���	������rQ���P� ����D�('_�\���7 ���9&�6V��ǃ��l��,H�����b˿GOϿX̿8¿sڱ�D��3��l�X�I�'�h���*d���Ga�h�	�����*tQ���P�����ZI��-_��   �   4;��$��[�����a���yȿ�	⿔���L ��}��y�9<�� 俷ʿY[���0���C]��%��{�t��|rA�3��*��74�~�U��b��K���!k�H��� �fB�ٷf�����{���Θ��ۛ��V���p���Մ��=i�([D�n ����`��_�n��y��@����[�>"8�z��8�ཌA��Ӛ��   �   ����Q��v�����,Կ������x��!�p;$�^�!������5�����տa/���+����Q���e�ʾ����:��O����,��}�R�E�x����T�4Nb��ܠ��n־~D�ߐ"�
�:�d?N���Z�~`_���[���O�?�<�#�$��%	�3�پ�����f���Oj���<O�fp��;3��%���\��?����ʾ�   �   y�8��������sҿ(A���m���'�@8���B�B�F���C�.9��)��u����<Pӿk꧿i+�LK8�u������x=��[ǽD86�R��̓���Z�������#3F��䈾M���Ȳ׾����:��H�Y������B��S����ھ��������~"K�����Ϣ���*�����X/����?��˽uF?������V���   �   ��Y��z���*ÿ�A�����,�F�D�2�X�6�f��
l��~g��Y��E�(�-���������ÿ����Y��]�����>�d���h�K�ЩA�@T;��E�P�ż�Un��;ѽ,��4�S�lք�����r��f������.潾,����"��)��@wX�&9!���ٽ~�P�Uʻ��1��p��W�C-���0h�0p¾S��   �   {�w��Ȩ�gxۿh'	��&���C��v`� Uy��B���m������\z�La��D�&������ڿ�৿��u�V*�vTݾV���9Z���f� o�`l�<@P�<pt]< z�6u������ܽ���x�4���O���`��Yg�00b���Q��"8��I����v����#���/��&<4�<hSe<(�-�̰t��'�����[�߾N�+��   �   c��跿��&��95���V��Gx�����F���^T���Ք��Պ��^x��V�ڣ4�@e�4��x��m)��.�:����������D3��s��L3�<��#=P�=��<�M<@��� -��F��0����D�.���j�Q���N/���ۜ����:�(b��н�;�2�<��=Fz=�0�< ��ᇽ�!!������Z���<��   �   �͎�H���O�������L?�4�c��E��?��2������8��S4��y���&c�J?>����w��������O��`E��`�܍����'�� ���r��<s=b`L=8�[=ت@=2r=�x<�b��z̼v�/���i����:��Sۉ�R�p��9�xV� ��X�B< ��<�3=.N=��>=��<��xV���P,������<��G��   �   �Z����Ŀ�������B�
�h�0+������������c��g���Sۆ�n�g���A�f������¿�Ï� I�����ӟ�|B+��Q��p8���j
=ֈY=-o=�[=F*=�6�<�6�;��4���߼��$�leG�N�T�l�J�4f+����pa�pل;(+�<��=V�M=�a=��K=��<��ж���60�O⢾&���~K��   �   ͎�s���>�������K?��c�:E��<>��1������7��~3������%c�r>>����s���û��O��(_E�`������'�m��pc��dt=,aL=��[=�@=Hr=�x<@c��<z̼��/���i����:��dۉ�f�p�9��V�0����B<���<�3=�N=��>=X!�<@���T��oO,�����;��G��   �   �a���淿���$�85���V� Ex���������R��%Ԕ�PԊ�$\x��V�F�4�d�B�iw��<(��k�:������f��l0��pV���7�<�#=�=��<N<P���<-��F��M����D�X���{�r���h/���䜑���:��a�� ��;4�<��=�{=�5�<����އ�T!�;����W��M�<��   �   �w��ƨ��uۿ�%	�v&��C�~s`�Qy�Y@���k������xz�a��D��&����F�ڿ~ާ�w�u��S*�Qݾ���,W��f��F�r�<�S�<�x]<�u�u������ܽ����4���O���`��Yg�H0b���Q��"8��I����\�����#��/�P&<��<�`e<�-���t�l$�R�����߾��+��   �   ��Y�Qx��6'ÿ�=��l����,���D���X���f��l��yg���Y�R�E�(�-�R�������ÿ����	Y�[�o�����d�����K���A���; �E���żUn��;ѽ2��G�S�yք� ���r��z������>潾:����"��)��>wX�9!���ٽ~��L⼰@ʻ��0�xp�h�W��%��+h�l¾P��   �   �8������Aoҿ�;���j�N�'�"�7�$�B���F�h�C�9��)��r������Kӿ�槿�%��F8��n��G����=��Sǽ.6��D������*X������3F��䈾X���ز׾���	;��H�d������B��S����ھ��������Z"K����Ϣ�D�*��}���!��{?��˽c@?����?P���   �   a���Q��r�����,'Կk����������
!�87$�<�!�8�������:�տ�*���'����Q�c�	�ʾ����4�H���{,��v�F�E�G���T�Nb��ܠ��n־�D��"��:�p?N���Z��`_���[�ʦO�E�<�&�$��%	�-�پ������f�R��h��l8O�zi�R13�i���V�;����ʾ�   �   �2�g$�Ɖ[�:�=����ȿ��o�������y��u�5�������ɿ*V��O,���<]�%��s�n��jA�Ә����:-4�0�U��`�����Z!k�:���" �mB��f�����{���Θ��ۛ��V���p���Մ��=i�)[D�j �����_����n�2y��>���[� 8��������@��͚��   �   ^���"���6&��2V��Ń�2j��cE�������^˿�KϿ�̿����6ױ�J��e0���}X���'�l����_���@a��	�6� eQ���P�-���D��&_�A���. ���9&�6V��ǃ��l��3H�����b˿POϿ_̿?¿xڱ�G��3��k�X�B�'�Q����c��Ga�v�	����jQ���P�O����A��"_��   �   fk��ꬾ��!����A���f�����y���˘�z؛��S���m��ӄ�s8i��VD����{��[����n��s�47����[��8�����ཤA��Ϛ��5辛$���[��}���<ȿ�ԑ��`���{��w��8��q��ʿY���.���@]�n%��x��q��<oA�j��X���/4���U�O]������   �   �P�VHb��ؠ��i־uA�F�"���:��:N���Z�n[_�y�[�̡O���<��~$�"	���پ鬣���f�R �?`���,O�*b�.3�����W�j<����ʾ����Q�Lt��u��s)Կ%���4��n���!�T9$�^�!�F�����|���M�տ�-��8*��f�Q�)��ʾ���n8�aL��2,��u�МE�z���   �   ق��z��-F�ሾ����&�׾����i7�E�[������>��L��f�ھǱ��̧���K�m���Ţ���*��j��(���x?�{�˽�A?�P���=R����8��W����pҿ
>��&l���'��7�L�B���F���C�D9��)��t������Nӿ駿_)��I8�s��H����=�wXǽ�26��E��d���ZP��   �   ��ż�Gn��2ѽ~��>�S�G҄�-��Om���������Oཾz������C$���nX��1!���ٽ��}��0⼀�ɻ��.���o�Z�W�&���+h��l¾�P���Y�-y��^(ÿ?��f��8�,�6�D���X���f�Fl�\|g��Y�^�E��-����5����ÿ����Y�*]�r�����d���V�K���A� �;�|E��   �   �]<p-��h������ܽN����4�S�O���`��Qg�&(b���Q�D8�=C�Ω�o�<�#��/�h:&<,��<�we<И-���t�P$�����_�߾J�+���w�.Ǩ�pvۿ<&	�<&���C��t`��Ry�]A���l�������z��a��D�^&���5�ڿ৿�u��U*��Sݾ򎄾�Y���f�0Y��s�<�Z�<�   �   r�=*�<�k<$̓�z	-��?��=����;ྲྀ���z�c����%佲俽x�����:�hH��@�;�E�<��=p�=�>�<@��{݇��!�����W��f�<��a���淿v��%�|85�j�V��Ex�����Z���|S��Ք�4Պ��]x�d�V�l�4��d���x��P)���:����������-3��Pl���6�<��#=�   �   t�[=ެ@=>u=�%x< :���m̼<�/���i�- ��[5���։���p��9��E������B<��<�3=�N=^�>= (�<��4S��xN,����;���G��̎�G����������K?�:�c�gE���>��}1��>��b8��4��P���&c�B?>�������������O��t`E�a�_���v�'��!���{���r=�`L=�   �   <T=�>=��
=���<��A������!� �Y��~�����)���]��Q'�Tü�ƚ���o<�=H-7=��L=�P5=�v�<8���BO����F�gJ��%��
�]�n���7տ��	��"-� �T��!��������;ص�wL���ӵ����֕�j�|�S��,�����{ӿ����[��`��*��L�C��
��+���r�<��<=�   �   ?=�Y"=���<�ն;�����a��bf��$���6�������c��tT��BOl��W����� �q;�&�<��=^�7=>H'=xǱ<�ر��B�B����N��M�Y����_wѿ���"$*�^�P� �z������8������������\/������xCz�8�O��9)�Z���п�噿X��������n�?�f��� i�����<��.=�   �   ���<��<`��1�Bge�-����ݽT������ʶ��C�46Ὃ-��b�m�x`���}��4��<x�<�/�<d��<$������[�6� &����� N�g��'&ǿl ���!��`E���k�OV��]8��{������~ߥ�+\���`����k���D�T� ��b ��
ƿ?-����L����0S��j�3��ɟ�[���7�<�=�   �    �v;���̔K�&�����)�~�M��'j���|�������}���k���O��3,��M������U�������:B<��;�������n�$�}���1g����;�߮��"���hv�Rx��h4�8�U��w�A������b����+���O��(�w�:V�Zd4��>�S��|L��<
��V�:������{��l"�ב�t>�����;��`<�   �   P�+ ���C��v�3�PAo�xʔ�c��� �þuKѾ�*־��Ѿ��ľ�c���e���r���6�����@	��س�ڀ��G!���˼j����g��ၾ
�־��$� �m��Z���iӿ0�����<��-W� qn�2y~�/3����<Oo�"X���<��H ��L�ONӿ���}�l��	$��`վÀ�
l�>���ļ�����Hc��   �   ���J����`��I���hľ0��
�W��"��E&��2#����R�Ӯ�Ǆƾ�6���d���������\�~V���{s��F�W�zL����
�N�I��׊��Ե����|�	�X!��6�X�H�JU���Y���U�ؤI�l�7��!�:F
�����!��f势:�I��g
�Ɠ��8V�;d�>�m���� c���AU��   �   >�)����9��:B����s2�N�L�Zla�p�n�Z�s��eo�Lzb�NN���3�\Y���ﾠ6�������+���ս�7����?�
�f���½٢+��A����߾#]$��Od�ү��I�����忮4�����%���.��X2��a/�$`&��q�p�<C�'᾿�;���d���$���߾���\�*����trb�b;�Lt~�o$ҽ�   �   �.��A3�����c+�2kT���{�Jq��2����@���w���흿�[��,�}�j+V��,����\����m��f�,�E�Խg%���Zl�*+�����FZ�,5��� �Z�3���o��_���p����ؿM������X��Te��"�l/��t��{~ڿ@����P���q���4�J~ �ҩ��\_Z����qn��$�i��b���wҽ��*��   �   )����!��]6�S(j���������e��i�пd\ܿ�y࿡�ܿ}�ѿ�����A�����M�k�ۤ7����վ�R�|���9���G���Ճ����E���{�T������Y6�t#j�㠏�s��'b����п�Xܿ$v��ܿ�ѿy���D?��������k��7����Ҿ�:�|����Q�������؃�$������{��   �   �
 ���3�E�o�Kb�� t��ٿ'�����v��ng��$�H1��w��[�ڿ�����R���q��4�� ����	bZ����fn��B�i��]���oҽ��*��*���-��P���^+�OfT�f�{�Cn���.������<���t���ꝿ�X��p�}�h'V���,�:�������j���,�f�Խ<$��4]l�5/��F���Z�69���   �   )`$��Sd�;���'�����忐6�Ԇ�L�%�6�.�<[2��c/�,b&�xs����E�%㾿B=��y�d���$��߾^����*�p����nb�l ;�lg~�ҽȁ)�b�G4��~;���Vo2�H�L��fa���n�Ԛs�R`o�Mub��N���3�V����n2�����N�+�P�ս�4���?��f�w�½�+�E��e�߾�   �   p�I��ي��ֵ����0�	�R!�P�6�ھH��	U�J�Y��U��I�@�7���!�hG
����J#��~抿ΘI��h
����c9V��d뽖�m�f���N��B3U�{�����=�`��D���bľ��!
�"���"�6A&��.#���������ƾ�2��)d�|�Ӫ����\��R����B�s�6L��W��O���
��   �   0�m��\��1lӿx1�<���<�V0W��sn�|~��4��`�tQo��X���<��I ��M��Oӿe����l��
$��aվ�À�0l�$Ȳ��`��H�b�
�N��q7��ֳ3�F8o�DŔ����þEѾ\$־��Ѿ��ľ�^��]a��X{r���6������� ��X΀��?!��˼c���hj�0䁾W�־Խ$��   �   F��������x�y�bj4�$�U��w�������������-���P����w�>;V�.e4�J?�.��M���
����:������{��L"��Ց�@6�� ��;0�`< �w;p�8�K��ⱽ���ϳ)���M�0j���|�M���	�}���k�ĽO��-,�@H�ﶽ�U�$���@��:HB< �;̽�����)�$�����Mj����;��   �   ����'ǿN���!��aE�*�k�FW��j9���������`���\��a��X�k�.�D��� ��b ��
ƿ_-����L����S����3�ȟ��S��4A�<�=���<�"�<�0���lWe�$��̹ݽ��* ��������>�i-��%����m��K�� >����<8�<�2�<��<L��������6�(��e���"N��   �   ���sxѿN���$*�N�P�$�z�H�+9��������j����/��,����Cz�D�O��9)�H��^п�噿�X�=��홮�h�?�����<b�����<��.=�?=$_"=��< �;\}���X�>Yf�r��N1�������^���O��>Gl��P�X�����q;0-�<��=L�7=�G'=ı<��������\�B�����_����Y��   �   �����տ,�	�\#-���T��!�������Tص�wL���ӵ������Օ��i��S�\,�L��+{ӿ�����[��_��)����C�I��d$��x�< �<=T=��>=��
=P��<@�A�d����!�^�Y��~�����5)����]�zR'�<VüpК�0�o<j=�+7=�L=�N5=Xq�< ���Q��4�F�~K�������]��   �   ����wѿ���&$*�L�P���z�q���18������ ��_����.��[���\Bz�L�O��8)����п�䙿�X��������&�?� ���@^��@��<��.=?=d_"=4��< �;�}���X�bYf����f1�������^��P��TGl��P�t���@�q;�-�<�=̘7=�H'=�Ʊ<��򲮽�B����������Y��   �   E���%ǿ7 �J�!�"`E���k��U���7���������qޥ�"[���_����k�f�D�H� ��a �E	ƿ,����L�G��4Q����3�mş�L��F�<~�=���<x#�<�.��异We�)$����ݽ#��? ��������>��-��%����m�tK���;����<(��<�5�<$��<@������l�6�)&����� N��   �   s��������u�w��g4��U� w�A���x������*���N���w�28V��b4�r=�B���J�����4�:�Ԏ��Iy��"��ё�l+��P�;X�`<��w;8��K��ⱽ����)���M�Lj�ҧ|�]���$�}���k�ٽO��-,�DH�ﶽ4U�����@�: #B<@/�;����Q��΁$�����f���;��   �   ҭm��Y���hӿ@/�~��"<�,,W��nn��v~��1����Lo��X���<��F �dK�Lӿ���u�l�x$�}]վ����Dh�ꂽ����8����b������Z7��޳3�Y8o�SŔ����þEѾr$־��Ѿ��ľ�^��fa��\{r���6��������x��$ɀ��.!�؝˼A���kf�&ၾؤ־��$��   �   ��I��֊�ӵ����P�	��� �@�6�0�H��U�
�Y���U�Z�I�.�7��!��D
�Φ�l��k㊿�I�ae
�F����2V�=\뽢�m�h��(F���0U��
�����4�`��D���bľ*��+
�-���"�BA&��.#���������ƾ�2��d��{�������\�N�j��us��C�W��J��z�
��   �   c[$�iMd�A���N���)��63� ���%���.��V2�^_/��]&��o����?�K޾�K9��4�d��$�4�߾���A�*������cb�^�:�c~��ҽt�)�=�D4���;���`o2�R�L�ga���n��s�_`o�Xub��N���3�V����b2�������+���սq2����?�ܔf�қ½h�+�A@��y�߾�   �   8 ���3���o��]��zn����ؿ�����\��>c�� �`-��p���zڿ!���N��Hq��4�x{ ������XZ����@f����i�TZ���mҽ&�*��*���-��P���^+�XfT�r�{�In���.������<���t���ꝿ�X��u�}�j'V���,�4��x����j��D�,�E�Խ� ���Rl��&�����Z��2���   �   �����W6��j��������(_��j�пUܿlr�C�ܿt�ѿ���<��沐���k��7�n���;��z|����*�������Ѓ�����^��^{�6������Y6�z#j�砏�z��/b����п�Xܿ,v�
�ܿ#�ѿ���J?��������k��7����Ҿ���|����6�����_у��������:{��   �   �'��*������[+�[bT���{��k���+������9���q��睿�U����}��"V���,��������f��v�,�R�Խ����Ml��&��^���Z��4��� �Y�3���o��_���p����ؿU�����\��Xe��"�p/��t��}~ڿC����P���q���4�:~ ������^Z�U��<j��.�i�Y���iҽ��*��   �   })� �0��'6�V��rk2�եL�ba���n�b�s��Zo��ob���M�H�3�R�ϝ��,��J��n�+���ս,����?�^�f�<�½̡+��A����߾]$��Od�ԯ��M�����忰4����
�%���.��X2��a/�(`&��q�r�=C�'᾿�;���d���$���߾���D�*������gb�L�:�*]~�.ҽ�   �   �������`��@���]ľ }
�B���"��<&�w*#�m�������_yƾ\-���d�:u�����$�\� D�D���rs�*D��W�BL����
�L�I��׊��Ե����~�	�\!��6�\�H�NU���Y���U�ڤI�p�7��!�<F
�����!��e势5�I��g
�����D7V�~a뽤�m����`>��F(U��   �   �������-����3��0o�����v鮾�þ�>Ѿ־Y�Ѿ��ľ�X��-\��Brr���6�0�������B�������!���˼%����f��ၾ�־|�$�"�m��Z���iӿ0�����<��-W�qn�4y~�13����<Oo�$X���<��H ��L�PNӿ���z�l��	$��`վ��k��삽$������X�b��   �   `)x;�ޖ��uK�ڱ�p����)���M�bj�V�|�����U�}�B�k��O��&,��A�V䶽��T�Th���r�:�DB<�_�;����3����$�H���g����;�ஆ�#���kv�Tx��h4�8�U��w�B������d����+���O��*�w�:V�Zd4��>�U��}L��<
��Q�:����`{���"��ԑ�X0����;��`<�   �   ��<�.�< ��@��Je����=�ݽJ����R��4��|9��#������m�(0�������<D��<�A�<�ǃ<���"�����6�&����� N�g��)&ǿm ���!��`E���k�PV��]8��|������}ߥ�-\���`����k���D�T� ��b ��
ƿ@-����L����S����3�gȟ��Q���D�<�=�   �   �?=\a"=���<�1�;�r��R�pQf����,�������Y���J���=l��G����@Tr;�9�<.�=N�7=�L'=�ͱ<�쒼���
�B�����L��M�Y����_wѿ��� $*�^�P��z������8������������\/������xCz�8�O��9)�Z���п�噿X����z���6�?������d�����<Z�.=�   �   �B=��,=���<�24<8��S@��z�R����,�������{��B�P��(�!���(<@��<�*=VB@=�&(=X��<@ڿ���ý�@T�xy��W���h������k޿D�� B5�^�_� ������������p��c���n�����Mf���c��bT_��4����{�ݿQa����g���1����R��Q��Tȸ��ȥ<z�*=�   �   �B-=�d=��< ܸ�4׹� D7�5����}��
��� ��jߤ�IB���&:��� ^���$�<h�=�}*=�=hy�<����(ʿ���O����!k�xbd��(��V�ڿz��
2�ڍ[�麄���Xܯ����{���H���ׯ�%؛�Ď���[���1�l2�&ڿ���F�c���������N�q�����|�<b=�   �   @A�< [T<H��j������Ͼ��T�Dx����Ν �1��	����Ԉ���ⅽ4E�h��G<pc�<$}�<,A<0XƼ%Q���jC��į�M��ICX� ����п��|)�eO��Dy���}��-w��մ������*���ȑ��'y��&O�T�(�rp���Ͽ4���5�W��i��﮾>%B��Q������xM<$4�<�   �   @e�(iм6�m��Iƽv��ha7�S�\��az���t"��I����"{�n�]�@~8����xȽ<�q�\�׼��H���;�%�:p�ּmU��s0��򞾀��FRE�����_��\(���O��L=�~�a�΂�_����T��64���r����������a��K=��3�c������Aˌ��D�h�bE���_/����8�м���:��<�   �   ��5��E���d�kB�[#�����s幾ŏϾ��ݾ9w��ݾоd����[���〾BqC�����`��rA9�~��(�x�́��m>��oz����B�⾕G-�(^y����ݿ�F
���'�̸E�^�b��C|� ц����������|��tc��F���'��V
��ݿߩ��	y��,��
�߇�������������m�XS���   �   ��ѽ��%��&q��h���о���������!� �+��/�6�+�>�!��m�����a�ѾTP��n�r��&��ӽrEz�|%�|�!�����N��-f�н�6��T�-����l��M��,�B�(��?��aS�J�`�XZe� �`���S�x@�RI)��y����ɕ��ާ����S���W}����e�|� ��և�z�Ho�w��   �   �-7��a��f����P���h�[1<���W��m�L�z����,{��m��0X�*�<����y���{������G8��	��ܑ��~\�J{���Mս�T8��A��ˇ��$-���o�6���ǿ������z��Э-���7��;� �7�,.�ZN����~��ǿ�\���;p��B-�	��)���8���Խ����xZ�d����b��   �   �"���̾�c��4�Ŵ_�qv��9���礿i	��?��>��7E�������`�K�5�p��\�̾����9�LN轠Y�����G���*��<+i������C�{=�|��񟿁o¿H\�|@ �����U�������'�� �m�_ÿ�k��V�|�8�=������Ui�H���>���.�������5�>O8��   �   \4ɾ����;@��Zv��䖿�Z��m�ȿ�ڿ��{��l��udۿ�<ɿn���o��7w�a�@��=���ɾ\����)��jӽ�����_����ҽ�s)�����O/ɾ����7@��Uv��ᖿUW��Λȿ-�ڿ�濏�꿧���`ۿ�9ɿ�����l��>3w�T�@��;�]�ɾ�Y���)��hӽE����b��>ӽ�x)�p���   �   �F��~=��|������r¿�_㿀B ����X�������)��� �i"��ÿ�m����|���=�ހ������Wi�����>��E,�������-�,I8�^��h ̾`���4���_��s������㤿����;���:��B�����i턿��`��5����b�̾ش���9�8J�_X��x���q������1i������   �   (-���o�����ǿI�𿸗����<�-�(�7�:;���7�P.�6P�X�?���ǿ`^��>p�RD-�p�쾑*��b8���ԽJ����pZ������X��&7�]�������I���d��,<�_�W�4
m���z�*��'{���m�,X�
�<�W�,t���w�����QC8���ّ��}\�^}���Rս�X8�E��q���   �   T�A����o��S���-�Z�(�r�?�ZdS�(�`�6]e���`�$�S�z@��J)�{����N��������S����~���e�ò ��Շ��s��d���v�i�ѽ��%��q�0c����оO������S�!���+��/�ѻ+� �!��i�~����Ѿ�K����r��&��ӽ�<z�x!���!����^Q�]2f��ӽ��8��   �   Xay���"ݿHH
���'���E��c��F|��҆�-���������|��vc�:F���'�nW
�>ݿ�ߩ�Ky���,���c���&��򿔽����H�m��;���5��;��N^�sB��������g߹�H�Ͼ�ݾ~p⾍�ݾiо捺��V���߀��jC����2Y��&79��q��h�x�P���xA��R}�
������I-��   �   o��[a���*��8Q�hN=���a�Vς�Ì��@V���5���s��(������Ԩa��L=�j4�L���j	���ˌ���D�Mh��E���_/�ݏ����м���:H�< ���Kм�m��>ƽ���Y7��\�Yz����������F{��]��w8�:��3oȽ`�q� {׼ #H� ��; ;�:��ּ�X��Vv0������TE��   �   Y���:п����)�vfO�vFy��Ñ����Px��ִ������+��]ɑ��(y�d'O���(��p��ϿW���M�W��i�u﮾�$B�iP��,����M<�@�<�P�<؁T<��6�����Tƾ�VJ��r����$� ��+�������݀��>܅�`:�(���G<�j�<X��<�)A<�^ƼJT��mC��Ư����1EX��   �   l)��u�ڿ&���2�܎[�����1��ݯ����������Rد�Z؛�ݎ���[��1�Z2��ڿߙ��܈c�������x~N������繼<��<f=PG-=^j=�(�< "��Hƹ��:7����^ꣽ`x�����������ڤ�>���:��濼@ʏ�l+�<��=z~*=��=v�<�����̿��O�����>l��cd��   �   ���hl޿���nB5���_�C���牟�����q��c���n��Y��f���c���S_���4����Чݿ�`���g�F��~��-�R�lO��\���(Υ<��*=��B=R�,=��< 84<� �܁R@�z�)����,������{���B�x����!�h�(<T��<L
*=�@@=�$(=��<4ῼ�ý8BT��z���W���h��   �   �(����ڿ���2�ʍ[�κ��J��ܯ�}��������Jׯ�vכ�(����[�*�1��1�ڿ-���Їc�������&}N�鞽�T㹼䆖<�f=�G-=�j=�(�< ��`ƹ��:7�(���wꣽux��Ż������ڤ�#>���:�翼 ɏ��+�<=�~*=��=�x�<X���F˿���O�����~k��bd��   �   ����wпؾ�$)�~dO��Cy�:����<v�� Դ������)���Ǒ�&y�r%O�6�(��o�5�Ͽ����M�W�lh���2"B�7M�����!M<tC�<�R�<؃T< ��<�����uƾ��J��r���:� ��+���������I܅�J:����G<�l�<���<�3A<\VƼQ���jC��į�I��-CX��   �   ����^��s'��<O��K=�6�a�<͂�G����S���2��q������j����a�J=�t2�7�������Ɍ���D�Zf��B��9\/�m���t�м@��:��<����Jм��m��>ƽ���Y7�"�\�%Yz���������`{� �]��w8�C��&oȽ�q��y׼�H����;���:H�ּ/T���r0�n�&���QE��   �   �\y� ��Kݿ�E
���'�P�E�n�b�PA|��φ�&��������|�drc��F���'�"U
��ݿݩ��y���,���@���������L���xqm�7��x�5�F;��<^�wB��������y߹�[�Ͼ
�ݾ�p⾢�ݾ}о�����V���߀��jC�|���X���59��l��`�x��w��'<��.y�����⾦F-��   �   0T����wk��Z���*���(��?�R_S���`��We�&�`��S��u@�<G)�x����E���ϥ����S���y��F�e�U� ��χ�Nl�<`��v���ѽ��%��q�1c����о^������_�!���+�/�ܻ+�*�!��i������Ѿ�K����r���&�:�ӽ�9z�����!�����L��+f�{ν�S5��   �   #-�h�o�����ǿH��4�������-�B�7�0;���7��.�$L���={��ǿ?Z��x7p�[?-�<�쾎%����7��Խ����<iZ�i����W罊&7�	]�������I���d��,<�j�W�A
m���z�8��'{���m�
,X��<�Z�-t���w��~���B8��齡ב�zv\��w���Iս�Q8��?��8���   �   �A��x=��|��m¿RY��> �����S�� �j���%�� ���ÿ�h����|�o�=�)|�!�qNi�4��/6���&��3���m+罎H8�6��X ̾`���4���_��s������㤿���;���:��%B�����m턿Ď`��5����L�̾����69�H��T�����������'i���   �   �+ɾ2���4@��Qv�;ߖ��T����ȿ��ڿ8�濯�����!]ۿ6ɿW��i��*.w�!�@�E8�,�ɾ�U���)�<_ӽ�x���Z����ҽ�r)�����//ɾ|���7@��Uv��ᖿZW��՛ȿ5�ڿ��濗�꿭���`ۿ�9ɿ�����l��A3w�S�@��;�8�ɾ�Y���)��eӽB|��'[����ҽ0p)�^����   �   h��`�˾k]�R�4���_�q��M����ि���L8��d7���>������ꄿ��`���5�5����̾w���%9��?轩O��w���򅯽���p*i�P����C�{=�|��񟿄o¿M\㿀@ �����U�������'��� �p�bÿ�k��V�|�3�=�	�U���>Ti����[:��(��菘�N'��D8��   �   �!7��Y��I���D��#a��(<��|W�m��z�|��_!{�&�m��&X�I�<�,� m���q����*<8�����Б�Nn\��u��iJսnS8�sA������$-���o�8���ǿ����~��ԭ-���7��;�"�7�..�\N����~��ǿ�\���;p�B-�݌��(���8��Խ����:hZ�]����Q��   �   ��ѽs�%��q��^��-}о���)��F}!�=�+��	/�Q�+���!��e����{~Ѿ|F����r���&�įӽ�*z�^�:�!�t��0M��,f��Ͻ�r6��T�.����l��O��,�D�(��?��aS�L�`�\Ze��`���S� x@�TI)��y����˕��ߧ����S���}��̈e�� �|҇��l�"\�J�v��   �   4�5��3��8Y� �A����ݐ��ڹ�L�Ͼ�}ݾ�i���ݾ 	о釺�VQ���ڀ��bC����N���%9�XU���x��m��	;��^y�|���⾍G-�*^y����ݿ�F
���'�θE�`�b��C|�"ц����������|��tc��F���'��V
��ݿߩ��	y��,�h
⾐��������������hm��*���   �   �-�d6м�m��5ƽ����S7���\��Pz�����P��J|{���]�Gp8����dȽƜq�X\׼�WG��5�;�u�:��ּS���r0���t��ARE�����_��](���O��L=�~�a�΂�`����T��74���r����������a��K=��3�f������Aˌ��D��g�-E��
_/�������м �:��<�   �   4Z�<��T<�_�v��������bA��m������ �&�l�������w��ԅ�(,����H<x|�<؏�<XGA<�NƼ�O��jC��į�F��HCX� ����п��|)�
eO��Dy���~��.w��մ������*���ȑ��'y��&O�T�(�tp���Ͽ5���3�W��i��﮾�$B�MP��@���pM<�F�<�   �   �H-=�l=D/�< ٲ�캹��37� ����壽fs��p�������wդ�9��N:�(ֿ� ܎��8�<D�=��*=��= ��< ���bɿ���O����k�ybd��(��W�ڿz��2�ڍ[�麄���Wܯ����{���G���ׯ�&؛�Ŏ���[���1�l2�'ڿ���G�c��������NN�����깼l��<�f=�   �   >3==�&=,��<��<P5��0���I��n���擽�4������� ���+H����>0��<�u�<~T(=�>=<�&=�4�<��Ƽ�tƽ��V��c����D�j��`��SA�>5���6�~Fb��P��]�������/��P���l0��Ǔ��?ˡ�a��dlb��7��U��u࿣���R�j�������n)W��\ǽ Xʼ���<X�$=�   �   �F'=�	=<W�<�	�<�ʼ�O@�����n���,5���2Ľ�
�� p��|P���;?��$ȼ����l8�<N�
=J�(=
�=�ǋ<�ȼ(�½dIR�M���o���sf����?�ܿb��2�3�:�]�mh��R���h��kͿ��k��RͿ�>k��%���u���^�<�3�����ܿ������f�a��Ἶ��R��ýxf˼��<J?=�   �   � �<�~7<3,�����>���tĽ�R��:������}#�A���^�������ýؚ������n&�hi=<� �<D0�<��6<��ͼT<����E����0_��KZ��Y����ѿ���j�*�R�Q�8r|�3ғ��������u��w��3���zғ�h}|���Q�(�*��	��ҿ�y��|Z�ӈ�|㱾b7F������мh�0<p*�<�   �   ƈ��$⼼x�T̽Z!�*:;�\�`�K�~��㈾+��,ֈ�`w~�d�`��:����'�˽�v��:߼@}z��$�; \�9$�޼�@���2������/�:IG�~v��x-��������bo?�(bd���������⪟��������׬������:\d�>s?���������G������tqG��Q��󠾔3������� t9p��;�   �   �0?����z�
��.F������T���ڼ���Ҿ\��4j�;�ྰ�Ҿj���z$��[��7�E�8x
��?����=�t;��x���V��./��(��ǳ��')�"/���{�<���Bd߿p���)��7H��f�`�����i܋�R���&��X�e�%H��x)�ȿ��l߿hʫ��|��=/�|[�uዾ���љ����䀆��۸��   �   '�׽~)���u��F��L�Ӿ97 �^�v�#�6�-�,1���-�X�#����  �ɰӾ����nu�D!)�e׽ޥ�8�#���&�|��0f�AGi�L"�����+uV�y<��J����K�����*�jvB��3V���c��6h�:sc�~V��XB�2�*�<��<񿿃�� ?����V�����B��Çi��������'��%��j���   �   ��:��ڊ�׳��<�������>��nZ��p��}�UO����}���o��IZ�#�>�ޘ���� {��ī��v�:���콵����Cb����mXٽ�,;��U��5��;F/�d�r�����Wpɿ0��$R��� �2�/�0�9�0=�p�9���/�� ��9���SYɿH럿��r�F/�_�ﾽe���R;���ٽ��@c��h��8M��   �   �����=Ͼ�x�pn7�I�b��<������&ꦿ���@%������tզ�9z���"����b��F7��Y�@Ͼ�i����;��a�q֜�����������T�l�SV���	���?�S�_���h�Ŀ�2�^���|�"�������Hi�ʽ���Q�Ŀࡿ�3��?�/	�oP���l��������S������.�;��   �   |8̾����B�x�y�ᘿ顳�˿�|ݿ�2�"3��!��_ݿ8�ʿ����Ø�Q}y���B����i̾���&�,�s�׽�[���a��E�׽��,�h/��`3̾B����B�U�y�ޘ�����f˿	yݿ�.�-/��T\ݿ�ʿ�|�����hyy���B�o��̾�����,�^�׽"\��e����׽��,�3���   �   �	���?��W�7�����Ŀ�6�h���~�d�������@k��������Ŀ+⡿87���?��	��R����l�n�����|Q���������;�{���'8ϾZu�j7�!�b�:�������榿���!��r���UҦ�gw��6 ��S�b�5C7�W�=
Ͼg���;��]�$՜�� ��͇��p��2�l��Z���   �   gI/�~�r����Wsɿ���$T��� ���/�Ŀ9��2=�ܰ9���/�� �T;����k[ɿ�쟿j�r��G/�љ�<g��T;��ٽ@����c��a��`C���:�L֊�����4��m����>�ziZ�,p�K�}�pL��,�}�M�o��DZ���>�\��`����v��y���ީ:���콛򔽪Bb� ���^]ٽ1;�8Y�����   �   rxV��>��׊��O������*��xB��6V���c��9h��uc��V��ZB���*�~��>�G���*@��7�V����	D��*�i�^��Ǉ��Z�'�D�$�4c����׽ w)���u�A����Ӿx3 �7
��#���-��'1�<�-�2�#�/��� �I�Ӿ	���gu�()�D׽��"�#�V�&�'���h��Ki��%������   �   &�{�?����f߿����)��9H�zf�T�������݋��������Vf��&H��y)����n߿\˫��|�}>/��\��ዾ����ϙ�����p��ĸ�� ?����
��&F�����O���Լ���Ҿ���fc徦�ྈ~Ҿߪ�����W����E� s
�[8��r�=�/������@2��������,徉$/��   �   �w��K/��S������q?�Ddd�Ԧ�����Z�������N������������]d�*t?�������0H��i���rG��Q���y3�������� �9��;�i���2x��H̽���2;���`�M�~�߈�a&���ш��n~�ϑ`�v�:�.��,�˽�v�D&߼�z��B�; ��9P�޼�C����2�Ż��)1�wKG��   �   [���ѿr����*�ıQ�t|�Cӓ�ᅦ���$v��m�� ���ӓ�D~|�<�Q���*��	��ҿz���Z�Έ�S㱾�6F�A����м�0<�6�<��<H�7<�,�P���6��
kĽH��������0x#����]Y�������ý������M&�X�=<d�<�3�<h�6<P�ͼ{?����E�����`��MZ��   �   ���^�ܿ���3�@�]�i����mi��ο�4l���Ϳ��k��U%���u���^�6�3������ܿz���A�f��Ἶ��R�5�ýd_˼t��<bC=�K'=  	=Pd�<����ʼ�E@�}��������/��X-Ľm��bk��AL��R4?��ȼ C��?�<j�
=B�(=��=lċ<�ȼ��½�KR�痼����uf��   �   Ca���A࿠5���6��Fb� Q������쎶�6/��P���R0�������ʡ��`���kb�&7�4U�-u����Z�j�$��\����'W�;Zǽ Qʼ,��<��$=5==��&=0��<��<5�\.���I�hn���擽�4��ͽ��� ��L,H�,���C0��<�r�<�R(=F�>=~&=�/�<� Ǽ	wƽ0�V��d�����;�j��   �   U���q�ܿt��:�3�*�]�Sh����ah���̿�k���̿��j��k$��u���^�j�3�@����ܿô��1�f�?
�
༾G�R���ý[˼<��<2D=L'=r 	=�d�<����ʼF@���������/��n-Ľ���rk��KL��h4?��ȼ B��|?�<��
=��(=��=ǋ<LȼO�½>JR�㖼����	tf��   �   �Y��Z�ѿP���*�ƯQ�`q|��ѓ���������s��S�����jѓ��{|�<�Q��*���ҿ�x���}Z�_��b᱾N4F������мH�0< :�<`�<P�7<0,�B���6��$kĽ2H��������Ex#����pY�������ý������ L&���=<(
�<�6�<��6<�ͼF<���E�&���,_��KZ��   �   v���,��3������xn?��`d���������������������m���t��� Zd��q?�~�������E������3oG��O�6��3�,����� ^9 �;`_�����x��H̽���2;��`�f�~�,߈�r&���ш�o~��`���:�:��'�˽Εv��$߼`�y�0T�; x�9�޼�?��@�2����-/��HG��   �   ��{�J����b߿����)�6H��f���������ڋ�Ĳ��4����e��"H��v)�N��Sj߿gȫ�m|� ;/��W��ދ�����ʙ���h�����R?�=��
��&F�����O���Լ��Ҿ���{c徻�ྞ~Ҿ𪼾���W����E�s
��7����=�*��|郼D���,����񲋾�'�.!/��   �   zsV�P;��Æ��J������*�rtB�b1V��c��3h�Rpc��V�VB��*�n���8�4����<��>~V�\���>��R�i���������'���$��a��Ʊ׽�v)���u�A����Ӿ3 �?
��#���-��'1�G�-�=�#�8��� �R�Ӿ	���gu��)�x׽@����#���&�a��xd�Ei�� ��Y���   �   cD/���r�����?nɿ���P��� ��/�Ⱥ9��-=��9��/�ȳ ��7�v��TVɿ�蟿��r��B/����)b��DM;��ٽf�����b�~_��B��:�5֊�����4��p����>��iZ�7p�W�}�vL��9�}�X�o��DZ��>�`��c����v��d���|�:�D��V�>;b�K���`Tٽ5*;�$T������   �   	�t�?��O�K�����Ŀ�/濤���z���H�����g�Ļ����ĿAݡ�-/�C�?�9	��K��b�l����s����K��U��e��k�;�P���8ϾXu�j7�%�b�:�������榿���!��y���[Ҧ�kw��9 ��Z�b�8C7�W�)
Ͼ�f��`�;�q[콣ќ�T��B�������l��S���   �   �/̾�����B�p�y��ۘ�ś��:˿�uݿ�*�A+�%�|Xݿc�ʿuy��'���Mty�n�B����̾�����,�ҭ׽�S���\���׽��,�#/��>3̾:����B�W�y�ޘ�����l˿yݿ�.�5/��[\ݿ�ʿ�|��"���lyy���B�k���̾~����,�6�׽W��c]���׽ �,��,���   �   {���4Ͼ�r��f7���b��7�������㦿���a������Φ�;t��P��4�b��>7�qS��Ͼ�b��@�;�S�h̜����?��L����l�V���	���?�S�a���i�Ŀ�2�b���|�$�������Li�̽���T�Ŀࡿ�3��?�#	�7P��D�l������DM��	��>�콻�;��   �   ��:��Ҋ�����=/������>��dZ��p���}��I��k�}���o��?Z�2�>�*��F����p��ޣ����:�h�콙锽�2b�u����Tٽ�+;��U����2F/�b�r�����Xpɿ3��&R��� �4�/�4�9�0=�r�9���/�� ��9����UYɿJ럿��r�F/�7��ne���Q;��ٽ~�����b�i\��<��   �   ��׽�q)���u��<��N�Ӿ:0 ����#�9�-�]#1���-�͙#��� �ͤӾ���	_u��)��׽܊���#�p�&����d�eFi�"��y��&uV�y<��K���L�����*�lvB��3V���c��6h�<sc��V��XB�4�*�>��
<���?����V����lB���i��������d�'���$�h]���   �   �?��殽��
�* F�����@J��ϼ��Ҿ�ྴ\���xҾפ��3��RR����E�}l
��-���=����ك�*���+����w����(�"/���{�=���Dd߿p���)��7H��f�b�����j܋�S���(��Z�e�%H��x)�ȿ��l߿jʫ��|��=/�U[�'ዾ����͙�����c�������   �   �(��8�� �w��?̽<�,;���`��~��ڈ��!��͈�f~���`���:������˽l�v�t߼�Ay�0��; ��9��޼V>��$�2�V���|/�6IG�~v��z-��������bo?�*bd���������䪟���� ���׬������:\d�>s?���������G������qqG�}Q�q��3�q���D�� 96�;�   �   ��<8�7<��+�j���/��$cĽ�>����\���r#����S�Q���2�ý΋��rv�P&���=<��<C�<�6<��ͼ�:����E�����)_��KZ��Y����ѿ���j�*�R�Q�8r|�4ғ��������u��w��2���yғ�h}|���Q�*�*��	��ҿ�y��|Z�ˈ�^㱾�6F�#���м��0<H=�<�   �    M'=�"	=,k�<�G�x~ʼ�>@�`���a����*��(Ľ	 ��f��5G���*?��ȼ�S��HL�<4�
=p�(=��=x΋<�ȼd�½-IR�@���m���sf����@�ܿb��2�3�:�]�mh��S���h��kͿ��k��SͿ�?k��!%���u���^�>�3�����ܿ������f�_��Ἶv�R�V�ý�a˼���<�C=�   �   ��B=��,=��<��9<�D�X��7;�vws�荋�
i��A���xp�� 7�tWݼ0R��xP<�N�<t�2=�H=$	1=�=�<�ߥ�ר���M��ڹ�h���c�7㡿�kڿ~p���1�:�[�)��P\���z��2ν�Xi���ҽ�ʑ��0����B��dd\��2����ۿfĢ�3Ie�F
�Ki���XP�P���ٳ�Tu�<��*=�   �   r?-=Π=Σ< ��8�@�2�?��g3����r�����|���h�}���-�dŨ��"�:h¯<p�=�<3=��"=��<���y���I��*��"-���_��&��^�ֿ�&���.�z�W��/������{�����������������s��]r��T-X���/����x�׿6���1(a��&�����L�U����Ҵ��j�<$�=�   �   4��<��X<�� ���Ё������<�v����&�~U���F��'ϸ��r}��O���ջPrq<���<��<��j<���l�h�=�T�������T�s.��Ն̿��G&�F�K�D�t�.��P��.���d��������R���u�CL�f�&�R���WͿ!ܗ��)U�`���߬�M�?�떰����qR<���<�   �   ���<:˼��i�O�ýN����4���Y�_�v�����ʗ���5���pu��X�?03�*�	�6���b���� ���X�"<�3|;D!��w���+�"��FE���A�秊�;F��@[��f�V{:�n
^����#������+���\���ԏ�%�����]��:��/�P����˼�"��<mB�;����?���,�)���!ʼ`;�8<�   �   V�1�nʦ�Ѳ���?�cD}�����^���в̾�4ھ�޾��پ��˾4���ʓ��]{��=�����<��Z�+�,���ؚK��W�������3���t޾G!*��<u��j���ڿ�q��k%�%C��_�V�x�����ł���i��v�w��?_�<�B��-%��a�jڿ蠟�f�u��*���޾Ւ��a5�9���(＠Ua��9���   �   D�ν�#��Yn�����8ξe���c3�Dp��")�b_,���(�������9���̾�C��d
l���!��?˽8Sl��������d���\���`�e��7����P�������w������&���=�x�P��P]���a�h�\��P��=�ta&�&$�FL뿢»�u���[�P�\��q�����a���������������q��   �   ��4�����_�������Q&:��U��.j�Ύw�|�(w�tui��)T��*9�������F������ �2�B�ཤ���P���x��Oνj�3�]H����|�*�ԯl��$����Ŀ�T��,��.���+��)5�X8�~�4�+�(�� �
�k�2;Ŀ9ɛ�\Vl��m*�_�����{4�ɸϽ�|��+T�OK��Wg��   �   �1��Ђɾ��	�H�2�c]�G�����T���٫�Ǯ�鐫�����	g���p���0\���1�%	�WȾ?X���4�Ի��8��h��]���5v
�g�d�L����P�V;�, y��9���}��	)�����*P
�|������G�X�	�����O�ڠ��6����Dx�o~:���?{��Ԇd���
��J���	��Z����}⽪T5��   �   ueƾu��>�~�s�_��������ƿрؿ��㿑���m���׿��ſ����Q���z�r��(=�2k�Нž�`��T�%��
ͽM��	{����ͽ�&&�\ڃ�}`ƾ, ��>�y�s�\��_�����ƿ}ؿ��㿶��9j�i�׿f�ſ2���������r��%=��h���ž�^��Ք%��ͽ�M��K~��9�ͽ�+&��݃��   �   vS�	;��$y�R<��Հ���,῿���JR
��������I�B�	�	���@!�X���@����Gx��:����}����d�F�
��J��H��D{��Yu⽬N5�r-��L}ɾ_�	���2��]]�i�������B֫��î�����u��Ed���n���,\�q�1��	�SȾxU��
4�ŷས7�����q����y
� �d�qĳ��   �   ��*�ӳl�l'����ĿX��.�(1��+�,5��Z8���4�*!+������
��m�>=Ŀ�ʛ��Xl��o*�Ĝ辉����|4�:�Ͻ.|��#T��D���]��4�����LZ��������!:�QU�_)j��w�`�{��"w�Spi�	%T��&9�@����������������2�w�ཚ��ЃP���x��Tν��3��K������   �   ֻP�����G���q��ƍ���&�R�=��P�xS]�N�a��\�>P��=� c&�`%�6N�#Ļ�������P�y��̚���a�����̗�����$����q��ν>�#�@Qn�D����1ξ���P/��k�+)��Z,���(����F���3����̾,?���l���!� 9˽�Jl����:��Dg��b��d�`��������   �   �?u��l���ڿbs��m%�4'C���_�&�x�5���?����j����w��A_���B��.%��b��ڿᥧ���u�Ө*���޾[����5����0�5a��"����1�;���\��ƹ?�;}�5���b~��f�̾.ھG�޾7�پ��˾́�����t�z���=����*5��.�+�����K�H[�������x����޾�#*��   �   R���H��g]�����|:�p^�:���|�����s,��$^���Տ�������]�҄:��0�9���>̼��"���mB�Ӡ���?����,�����ʼ`t; [< �$˼��i�L�ý���b�4���Y���v����=���\1��khu�}X��)3���	�o꿽>�b���� 3�� �"<�?|;L&��(z��H+�:$��oH���A��   �   �/��M�̿����H&���K���t�0��j��+/���e����z�������u��CL���&����$XͿDܗ��)U�_��{߬�İ?����\��0�R<ԩ�<̟�<��X<x������ȁ�Y���N2� ��g����P���
�6��JǸ�fe}�$E� Wջ��q<$��<��<��j<���|��=�>���^���T��   �   �'��u�ֿ4'���.�v�W�b0��N��j|������F�����	������xr��d-X���/����G�׿ ����'a�h&�T����	L�x����˴��q�<0�=D-=B�=�ڣ< ��84߳���2�,��.���볽�l��w��֛��&�}���-�Ĺ�����:�ȯ<��=�=3=D�"=p�<`��3��<�I�',��8.�	�_��   �   �㡿=lڿ�p� �1���[�j���\�� {��Kν�Xi���ҽ�������{B���c\���2�z�^�ۿ�â�@He��	�-h��WP�����ҳ��z�<��*=��B=��,=��<H�9<h?���6;��vs�����i��c����xp��!7��Yݼ [�sP<0L�<ز2=2�H= 1=D8�<�楼)�����M��۹�%���c��   �   '����ֿ�&���.�n�W��/��p��i{��o���*����������
���q��V,X��/�R��]�׿K����&a��%�U����L������Ǵ��t�<�=�D-=��=ۣ< ��8@߳���2�;��%.���볽�l�����盞�H�}���-�๨�@��:8ɯ<Π=f>3=�"=�<4������I�++��}-� �_��   �   Q.����̿���RG&���K�v�t�������$-���c���������M��.u��AL�L�&�j��cVͿ�ڗ��'U�����ݬ�H�?�J���L����R<��<���<��X<p��֛��ȁ�j���l2���|����1P���
�X��fǸ�xe}�E��Uջ��q<ж�< ��<��j<���]�z�=�\�������T��   �   y����E��^Z��� �vz:�4	^�1�����p����)��z[��bӏ������]�J�:��.�%����ɼ�� ��kB����==����,�����`ʼ��;�c<���˼H�i�@�ý���n�4���Y���v����L���j1���hu��X��)3���	�o꿽
�b�|�� �����"<`v|;T���u���+��!���D��b�A��   �   2;u��i��Rڿq��j%��#C�4�_��}x�[���L���h����w�=_�"�B��+%��`�ڿ����D�u���*��޾>���z1�غ�����x$a�d��,�1�Կ��F��¹?�;}�<���o~��v�̾$.ھY�޾K�پ�˾݁��%�����z���=�����4��̔+�(�����K�N优���޲�b���<޾_ *��   �   ��P�a���J𻿎��Ί� �&��=�0�P�N]���a���\�R�O�X =�h_&�f"�MI�"���k���!�P����ӕ��n�a��������n~������q��ν�#�)Qn�B����1ξ���Y/��k�4)��Z,���(����N���3����̾0?���l���!�B8˽�Gl�,�����a��SY����`�������   �   ��*�^�l�W#����Ŀ"R�j+�*-�t�+�:'5��U8��4��+����0�
��g�C8Ŀ�ƛ�ZRl��j*���输|���u4�`�Ͻ��{�T�eB��R\㽂�4�����AZ���������!:�ZU�f)j�&�w�l�{��"w�_pi�%T��&9�E����������t���B�2�(��b���|P�|�x��Kν��3��F��|���   �   �N��;��y��7�� {��&�]���BN
�h�����tE�>�	������࿧���r����?x��z:���v��J�d��
�B������w��.s�	N5�G-��5}ɾ[�	���2�^]�l�������H֫��î�����z��Jd���n���,\�t�1��	�	SȾPU��p4����>4��N������s
�ͦd������   �   "]ƾ�����=���s��Y������אƿ�yؿ��ފ�]f㿨�׿ܷſ񻮿�����r��!=��e���ž�Z����%���̽oE��v��Ӝͽ�%&�ڃ�W`ƾ$ ��>�x�s�\��a�����ƿ
}ؿ��㿻��?j�o�׿m�ſ7��� �����r��%=��h�w�ž�^���%��ͽ�H���v��ךͽ%#&��׃��   �   �*��Lyɾ��	���2��Y]�����������ӫ�_���L���.|��-a���k���'\�-�1����MȾ-Q��t4�{�� /���������t
���d�����P�O;�* y��9���}��)�����,P
�~������G�\�	�����T�ޠ��9����Dx�l~:���
{���d���
�FF��(���v��'o�oJ5��   �   �4�W����U����������:��U�F$j���w���{��w��ji��T��!9�*������N���
�����2�������~tP���x�9LνN�3�	H��׊�p�*�ϯl��$����Ŀ�T��,��.���+��)5�X8���4�+�*��"�
�k�5;Ŀ;ɛ�\Vl��m*�8������y4�J�Ͻ��{�(T�h?���V��   �   )zν�#�mJn�팡�J,ξ�����+��g��)�tV,�)�(�n��C��E,��_�̾�9����k�Þ!��-˽�8l�������F`���Y���`�%��(����P�������x������&���=�z�P��P]���a�j�\��P��=�va&�&$�IL뿣»�w���V�P�P��7�����a�2��������~����>�q��   �   �1�}���N��]�?�"3}�����y��y�̾�'ھ��޾��پ��˾�{��ȉ��4�z�Ί=�@���*��<�+�$���paK�D�w�����⹆�I޾>!*��<u��j���ڿ�q��k%�%C��_�X�x�����Ƃ���i��x�w��?_�>�B��-%��a�nڿ񤧿h�u��*�}�޾����V4�ὑ� �a�p���   �   ���˼��i��~ýn���4�>�Y�}�v��{��Ď���,���_u�rX��"3�`�	��߿���b��轼 ����#<��|; ���t���+��!��*E���A�槊�;F��@[��f�V{:�n
^����$������+���\���ԏ�&�����]���:��/�S����˼�"��:mB�$���n?��P�,�ʷ���ʼ �;@r<�   �   ��<�X<���4����������h)�������J�f�
�:��0���JU}�(7���ԻX�q<8��<<��<�k<h����묽��=�3�������T�s.��Ն̿��G&�F�K�D�t�.��P��.���d��������S���u�CL�h�&�T���WͿ"ܗ��)U�Z���߬�ذ?�e����	���R<��<�   �   xE-=��=��< ��8�ӳ���2�!���)���泽�g��7������J�}���-�T������:�կ<(�=�B3=��"= �<,���
���I��*�� -���_��&��^�ֿ�&���.�z�W��/������{��ᆹ������������r��^r��V-X���/����w�׿7���0(a��&�檷��
L�����\δ�$q�<��=�   �   mR=�w==Ԃ
=4Q�< �`2���n�PzM�*�n��Cy�r�k�zH���3�� }�9䝟<~=��H=��]=)G=$,�<�M>�[2��>�:�ȍ��3���+U�
�����Ϳ)��"'��M��v��[������'����R������Ţ�������w��HN�R(��9��OϿx_���\W�g7��/��v?�ZT��x�p�\��<��;=�   �   v�==*�!=���<��;8�q�|��P�[�2+��p���Ur�����V�� �S�>m�WH� �<<-�<��,=�-I=�l9=��<h�@�5ҝ���6�q����	��YQ��a���2ʿ��8`$��qI�d�q�E�����h���9��G���|���z����r�FqJ�4m%������˿Y���jnS��y�٢���;��ʤ���r�XS�<F.=�   �   �Z�<�2�<@�ʺhۼ�`]�%t��p%ֽzY���;
�>��^	��!����ѽH���R��ü@�:$4�<.v
=�+=��<��L��`���+�������>F�lލ�kv�������l���>�|	d��������⮟�냣�,���=���)���Qd���?�x!�������������H�|���f��pG/��䚽Hd|����<=�   �   ���;�׎��E�������
"%���G���b�(-t���y��s���`�GE�4"���������n8�(�m����;���<H�5<��n��憽R7�����I6�m�4����v#��OM濘(��3/���O�oo��x��Ԏ����f��������n��UO��?/��o�H����>ӂ��46�6w�Ӥ���x������8���<�Yi<�   �   �������1�Nw/�Ôi�b%���k���R����ʾϾL@ʾ���򺨾[;����e�J�+����qK��$� K$�Pː�����Rq�
F��:w�x�;�����e�_p���}ͿW� ����K7� kQ�|�g�Ftv��{�X�u��f�:xP��6�nz�� �ӧͿ̝���f���L�Ͼ�z�J����z�����а໐�N��   �   �<�����^|[��ӕ�@�����x����2-��"!�N��z;�֡������������rW��O��K����A�P"ۼ��@�Y��~޽�5M��#�����]hC�M܆�h��|޿����i��i2��C�jO���R��rN�X�B��U1�n�����ݿ�ð��Ն�6�C�ZG�w��V$O�u^�0�a���=�~'L��   �   4�$�*�x����� �)��}~.���G�Q�[�?nh��l�&�g�íZ��oF���,�='��9�\ì���t�C�!�$�Ž�lj�L�(�2SO�(B��++#�����s6ؾ�f��^���G����῔u�W� �!��u*��G-�F�)��� �R�"��M�߿����a[���|]��4��Jؾ'���1$�ķ��*�T�hh/�Jr���ʽ�   �   ����g��L� �l�'���O���v��M�����*١�و���c����6G���tt���M�,�%�Z����f��8~�)#��xƽ.�z�^W�����;���|�Q���������G"/�3
j�[������ĩԿ���d��2Y	�D��v������2�ӿg;��}���ԟh�6@.�^������8@Q����o��4LZ�|c���ɽR>%��   �   ^Q����g2�f
e�����	����i��k[̿-�ֿ�iڿo\ֿ	>˿����9���r���c��0�Z��Z���@7q�)��i��Jjt��u�y{��Ю�|�r��L�����x2��e�Ǥ��瓥�Of���W̿~�ֿAfڿ�Xֿ�:˿	���6���p��c�@�0�6��O���83q�̩� g��`kt�u�`���y��E�r��   �   �����%/��j�������5�Կl��d��@[	�L��j�����6��ӿ�=��m����h��B.���������BQ�����z���GZ��Y�۔ɽ�8%�/}��db���� �Z�'���O���v��J��߅���ա������`��
����D���ot���M��%�f����b�� 	~��#��tƽ��z��W�h��+����Q������   �   �i�N^�������hw�Y�P�!��w*��I-�j�)��� ��S������߿�����\��]�/6� Mؾ����`2$�*�����T��`/��=r���ʽ�$�Үx�p����@��z.���G��[��hh��}l���g��Z�?kF���,�$��4�K�����t��!���Ž*gj�H�(��VO��F��/#������:ؾ�   �   bkC�<ކ�����~޿2���k�l2�D�C��O�l�R�
uN�j�B��W1�ހ�D����ݿUŰ��ֆ�ĬC�fH�����%O��^⽼�a����)�(L��2��&�� t[��Ε�6�����辟��i��(�E!�5���7�c������}��ۆ���kW��J�fE��h�A��ۼ���&�Y��޽�9M��&������   �   ��e�;r�� �Ϳ�� �����M7�^mQ��g��vv���{���u�.�f��yP�F�6�v{�� �
�Ϳ�̝��f����P�Ͼ~z�t����z�민0s�P�N����󬑽���o/��i�J ��If���L����ʾ�Ͼ>:ʾ���ڵ���6��A�e�E�+�;��|D��h��3$� ��������q��H��>w���;���   �   ���!%��UO��)�`5/�P�O�*qo��y��GՎ�2������� ��t�n��VO��@/�Np�'翪����ӂ�56��w�����x�ܷ���0���&<zi<��;L����E�q��ƈ��%�6�G�n�b��$t���y�`s��`�JE�!"��������a8� gm�0�;��<�5<�n��醽�9�����B9�{�4��   �   �ߍ��w�������m��>�d�䎄����䯟���������������Qd�x�?��!�L����������H�x���f���F/�2㚽�U|�茖<�=�i�<�D�<@Aɺ��ڼHQ]�Kk���ֽ"O��86
����Y	�8���ѽ�@��LR���ü��:\?�<�y
=l-=��<�M�dc��G�+�� ��&!��@F��   �   �b���3ʿX��`$��rI�r�q��E��o�����	:���������{���r�VqJ�0m%����s�˿'���nS�4y�B���� ;��Ȥ��r�lZ�<:.=��==L�!=���<P�;wq������[�'&��H���Mm������Q��N�S��f�(AH�@<p3�<��,=t.I=Hl9=���<�@��ԝ���6������	�W[Q��   �   ����8�Ϳr)�H#'�
M�V�v��[��ޤ��?����R������Ţ�y����w�lHN��Q(�p9�`OϿ�^���[W��6��.���?�R��0�p����<"�;=�nR=8y==P�
=�S�<���<0���m��yM���n�vCy���k��H����5�� ��9p��<�|=�H=�]='G=$'�<�Z>��4����:�Ҏ�����,U��   �   &b���2ʿ��@`$��qI�:�q��D��������9���������Ez����r�`pJ�vl%�J����˿{���mS��x�O�����:�gǤ��r�]�<  .=`�==��!=(��< �;�vq����Ƥ[�?&��\���cm������Q��f�S��f�XAH�X<�3�<8�,=�.I=m9=h��<0�@�@ӝ���6�����	�^ZQ��   �   Mލ�3v�������l�^�>��d�z���l����������)���=���?����Od���?�p �-��p������H�$���d���D/�#���PF|����<t=�k�<4F�< 8ɺ`�ڼ>Q]�]k���ֽFO��J6
���Y	�X��"�ѽ�@��jR���ü��:(@�<�z
=�.=T�<��L�q`����+�������>F��   �   ���"��{L�(�3/�h�O��mo��w���Ҏ����!��������n�TO�R>/�vn�:�Y����т�p26�t���fu�����&���4< �i<���;����E�a������%�G�G���b��$t��y�xs�"�`�bE�4"��������a8��dm�@�;��<@	6< �n��冽�6�J����5���4��   �   ��e�o���|Ϳ�� ���XJ7�liQ�f�g��qv�p�{���u���f��uP� �6��x��� ���Ϳ4ʝ�óf�����Ͼ�z������z�(ޯ�PR�МN�~���������o/��i�P ��Tf���L����ʾ�ϾQ:ʾ���굨��6��O�e�L�+�"��.D����*$����8z��q��D�9w�Q�;���   �   �fC�<ۆ����Jz޿j��^h�,h2�ΪC�O�h�R�.pN���B��S1��}�x��&�ݿ�����ӆ�%�C�E���BO��V�лa����!�nL��1�����t[��Ε�5�����辥��p��(�N!�?���7�k�����}��߆���kW��J��D����A�ۼ�r�v�Y��{޽�3M�?"������   �   8e�1^��Y���h�$t�^U�*�!��s*�jE-� �)��� �P�P���߿ݩ��Y���x]��1�dFؾ��,$�������T��Y/�9r�P�ʽ��$���x�a����?��z.���G��[��hh��}l� �g���Z�IkF���,�$��4�G�����t���!�m�Ž�bj�d�(�8LO�b>���(#�뛉�4ؾ�   �   3����/�#j�m��+�����Կq�￘��@W	�:��l�����/�ҿ\8������q�h��<.�������
:Q�����p��=Z�S���ɽ8%� }��Jb���� �W�'���O���v� K��⅙��ա������`������D��pt���M��%�f����b���~�,#��rƽ6�z���V�y���@����Q�>����   �   �I��Ы��2�e�����M���Zc���T̿��ֿ�bڿEUֿ67˿����3���m��Rc�X�0������+q�;��<^���[t�Lu�jx��ޭ���r��L����s2��e�Ǥ��铥�Sf���W̿��ֿFfڿ�Xֿ�:˿���6���p��c�C�0�2��1����2q���5d��
bt��u��v�������r��   �   fz���^��x� �*�'��O��v�^H�������ҡ�u����]����A���jt���M���%������]��� ~��#��jƽv�z���V�g���������Q�k���z���>"/�.
j�[������ĩԿ���f��4Y	�D��x������2�ӿj;�����ןh�6@.�F������{?Q�����i���?Z��P���ɽ�4%��   �   B�$���x�N�������-v.���G�<�[��ch�1xl���g���Z�efF�M�,�) �.�����O�t�d�!�U�ŽpVj���(��HO��>��*#�C���F6ؾ�f�^���F����῔u�W� �!��u*��G-�F�)��� �R�$��R�߿����c[���|]�z4��Jؾ�����/$�l�����T��X/�t3r��ʽ�   �   h+��8���m[��ʕ�$￾���.�����$�!����3����&{� x��Ձ��vcW�QD��:����A�x�ڼ�f���Y�|޽�4M�|#�����UhC�L܆�g��|޿����i��i2��C�nO���R��rN�Z�B��U1�p�����ݿ�ð��Ն�3�C�NG�A���#O��[���a�����XL��   �   �������\��i/�r�i����:a��/G����ʾ� Ͼ4ʾ����P����1����e��+��齔:��b
���#� ^���p���q�E��9w�K�;�����e�^p���}ͿV� ����K7� kQ�~�g�Htv��{�Z�u��f�<xP��6�nz�� �اͿ̝���f�ޢ�'�Ͼ�z�L��\�z��᯼pB່�N��   �   P)�;ȧ��4�D�����~���%�N�G���b�dt���y��s���`��E�C"�����gu���P8�.m��m�;$��<� 6<8�n�}䆽�6�~���-6�g�4����v#��NM濘(��3/���O�oo��x��Ԏ����f��������n��UO��?/��o�L����@ӂ��46� w���x�����(+���6<x�i<�   �   �r�<8Q�<�>Ⱥ<�ڼ�D]��c��Tֽ�E��81
����T	�"����ѽ8��R�T�ü o�:xR�<ԁ
=�4=`(�<��L�_��u�+�������>F�kލ�kv�������l���>�|	d��������⮟�샣�,���?���)���Qd���?�x!�������������H�v���f���F/�㚽8R|����<�	=�   �   �==��!=P��<�.�;�aq����[��!������gh������L����S��]� "H��#<�?�<N�,=83I=�p9=H��<��@�|ѝ���6�c����	��YQ��a���2ʿ��8`$��qI�d�q�E�����h���9��F���}���z����r�HqJ�4m%������˿[���knS��y�̢���;�ʤ��r��Y�<�.=�   �   R�i=�NV=�<'=Г�<H3 <�L�lvȼ����2���;�\].� ~��б�0�����><ly�<��8=gh=��{=xAg=� = �n:X�x��O��ݖ�����?�{}���ɺ��w�����9���\�����[��1��e�������t}��>��Z�]��\:�f&�u����ݼ�00���gB�t����_���9%�����z��O=,�T=�   �   8�V=̰<=�l=��{<��0���z�!�mW�
�x��O���Ht�@O��T��^�� @)7�.�<D=p�N=�i=|�Z=�;= C:քr�ڷ�����*���N7<��!��[�������d���5�FkX���z��H��݄���#������U���{�r<Y��7�؏�z��������C�>���������w!��}�� c����=j;H=�   �   b�=�^�<��< �t�6�#�&������Yӽ(�3�ｱ�潇�ν>����x�^���H-���O<�t =��.=|R3=0�<  �5�a��g�������羧2��A��,Ѯ�4^�<S�h�,�D�L�� l����>����������x��|l��M�Ή-�,�?�OW��ʒ��gL4�zf�:������ެt�`j���Q�<0l!=�   �   8�a<@�л<��o7���Խr}��-�ԷE�0BU��Z�H�S�dC��U)�V'	�Ѡʽ����� �����\��<0��<��< �6HI������y��Ѿ/F"�N�j��Ġ�_�ѿ�R�� �$n;���V�ȿm�
l}��f���|�Fm�<�U�� ;�.�����ҿu�����l���#�1�Ծ��~�KW��tZ��Zǻ���<x+�<�   �   `Ƹ��d�X�ɽ���L�d���▾)� W����p��MD������z�ףF�����A���Q�@]�� �;���;�λ�/��ݽT�V��y��*��;O���������������Y&��=�x�O�ֈ\���`��[�@�N��<�l�%�Ԇ��k꿹)�� ���HP�%>�T�����Z���6@>� �"� yd;@��   �   ?I��f��4?��3������gоeJ�������L��R����i���̾�_�������9��!�	����� \��Bi��5��µ�i�0�ї���_�/�&�s�ޠ���ʿu���j�"��51�;�x3>��[:�� 0�� ��d�� ��}�ɿI�����s��0���e���k3��H��B�&����|����~��   �   X����Y�25���&Ͼ���~ ��F4��vF���Q��U�`Q�f E��c2����� �˾��|�T�̷��枽�V*��4ݼ�[��x����
���p�E+�����`VH�S/��)ᨿ�3Ϳ���RF��Z����w��p�,[�F ����Q�˿�����z��a�G�����C����q�������������	6�?諒�   �   >$a�DX���R�p����;��_�)U~��N���蒿/R���\���R����{��{\�'&9�}�����w���?]�N=
�.�����:�X>�rc�8�ν�D5���_�ݾ�m��rS��)��+8��������ڿ�Q����v\��B���'����ؿs㿿���m酿x�Q�DR���ܾ�a��\�4�~Ͻ�f�h��bA�ϋ���F��   �   Dd��]��4< ���N�c��w������l!��E�ÿ��ƿ�ÿ0Ӹ������Ք�c|�1�L��o�F�N�����Q�P��������5��6�����{��UT��_����뾛8 ���N�F�~��t����������ÿ��ƿ�ÿ/и�
�OӔ�T|���L�(m�^�辇����Q����������5��7���������T��   �   E�ݾ�p��vS�!,���:�� ���<�ڿFU���(`��̒��m����ؿ濿.���6녿G�Q�eT���ܾ�c����4��!Ͻ�f�0��YA������A�a��S���L澹��1�;��_��O~��K���咿;O���Y���O����{��w\��"9���������|]�,:
�����r�:��@�xc���ν�I5�����   �   ����YH�{1���㨿�6Ϳ���*H��\����y��r��\��!�I���˿k����{����G�����E��J�q�������������^�5��楽����Y�O0��� Ͼ-��g��B4�rF���Q���U��Q���D��_2�v��� � �˾R����T����ួ�Q*�3ݼZ_� }��0�
�"�p�./���   �   !�/���s�@࠿6�ʿx��\l�"��71�D;��5>��]:��"0��� ��e����/�ɿ������s��0������l3�#I����&����\x���q�;@������,?�//��-���о]C�;����k��FN����Wc�W�̾9[�������9��������[�(Di�B:��ǵ�:�0��ӗ����   �   �>O�C�������#�꿀��Z[&��=���O��\�4�`� �[��N�`<���%�ć�5m��*��� ���IP��>�@�����Z��@>>�(�"���d; ������2d�)wɽ����L���Zݖ��쨾gQ�����j��'?��a����z��F�(��D9����P��K�� �;`��;0ϻ�/���ݽ6�V�u|��,��   �   ��j�^Ơ�9�ѿ�S� "��o;�Z�V���m�(n}��g�� �|��m���U��!;��.����~�ҿ���v�l��#���Ծ�~�2W��rZ��<ǻ��<�:�<H�a<paлZ���-����ӽw���,�<�E�V:U��Z���S�T�B�0O)��!	���ʽ쌁�����y�8��<ȿ�<\��<�:��MI�A��S�y���ѾH"��   �   �B��tҮ��_�&T�|�,���L�t"l�ٟ����^��m���|y��bl�rM�>�-�v��忋W��ꒁ�|L4�vf������Z�t��O��tZ�<�q!=H�=�o�<0<��t���#�	��ӏ���Oӽm齋��^��۶νG6��:�x�����#-�0P<z =�/=�S3=D�<  ��@�a�j�,���*��C2��   �   R"��N���ɜ�pe�X�5�*lX���z�nI��^���$�����V��" {��<Y��7�ԏ�]���么���>�����9���v!�R|���I����=?H=R�V=��<=rr=��{<��~�������!��cW���x�WK���?t�:	O�|M�XR��  z7�6�<�F=P�N=l	i=N�Z=R:= PB:��r������������8<��   �   �}��Eʺ�Nx�R��69��\�����[��E��f�������O}���=����]� \:�
&�����Sݼ��/���fB�'����^��"8%����� �z�0R=�T=��i=PV=>'=D��<8 <�H��tȼ ����2�t�;��].��~�8ұ�`�����><w�<��8=�eh=�{=�?g=T�=��m:n�x�JQ��ޖ�8�����?��   �   �!������Л��d���5�$kX���z��H������0#����KU���{��;Y��7�.��W�� ���E�����>�����Z���u!��z��P:��2�=�?H=��V=�<=�r=P�{<��~�̧����!��cW���x�eK��
@t�^	O��M��R��  x7�6�<
G=��N=�	i=��Z=n;=��B:r����'��������7<��   �   tA���Ю��]��R� �,���L� l�q����������ھ��x���l�zM���-�>���V�������J4�d�p���ޮ���t��2��D_�<s!=B�=�p�<p<Ȥt���#���ߏ���Oӽ�齧�ｃ����νg6��j�x���p#-��P<�z =�/=0U3=�	�<  6�a��g�������羑2��   �   ��j�JĠ���ѿ4R� �2m;�J�V�2�m�*j}��e����|�<m�f�U�0;��,���̖ҿ佡�-�l���#�V�Ծd�~�1T��jZ��ǻ��<�>�<h�a<�Zл���-����ӽw���,�K�E�k:U�Z���S�l�B�BO)��!	���ʽ򌁽d���h�D��<���<X��<���FI�T��ߊy�}�Ѿ�E"��   �   �:O�����l���F��&���X&�t=���O�Ȇ\�ĺ`���[��N��	<���%�`��Di꿠'��_���EP�<�?����Z����4>���"��)e; ������Hd��vɽ����L���`ݖ��쨾uQ�����j��7?��p���!�z��F�0��39��2�P�0I���;P�;�λ
�/���ݽ��V��x��?)��   �   ��/�0�s��ܠ���ʿs��`i��"��31�;�P1>��Y:��0�0� ��b������ɿ���+�s��0���@	�� g3�\A����&�̗���o��o�f?����p,?�%/��(���оcC�@����r��NN����fc�d�̾@[�������9���X�������[��*i�n0������0��ϗ�����   �   G��=TH��-��aߨ��1Ϳ���D��X����u��n�:Y�r�X��]�˿���lx���G�A���?����q���#������L���5��好+��ƻY�@0��� Ͼ*��g��!B4�
rF���Q� �U��Q���D��_2�|���� ��˾M��ԍT���������M*�X&ݼnU�\u��n�
���p�)���   �   D�ݾdk��oS��'���5��A�����ڿVN�\����X��������쿐�ؿR࿿6���煿p�Q�	O���ܾ0^����4��Ͻ��e�P�xSA�����A��a�hS���L澳��/�;��_��O~��K���咿?O���Y���O����{��w\��"9���������4]��9
�����j�:�7��c���ν�A5�����   �   ]������5 �I�N�3�~�Cr��É������ÿI�ƿ[ÿ�̸��yД�J|���L��i����#���Z�Q���������5��6�����?y���T��_����뾕8 ���N�C�~��t����������ÿ��ƿ�ÿ3и��SӔ�[|��L�)m�V��j�����Q�Y������5�d�6����u��.�S��   �    a�P��(H�̰���;��_��J~��H���ⒿLL���V��M��P�{��r\�D9�����O���]�u4
���Z�:��2��c���ν�C5����>�ݾ|m��rS��)��*8��������ڿ�Q����y\��F���,����ؿw㿿���q酿y�Q�BR���ܾ�a����4�(Ͻf���zQA�K���=��   �   R��H�Y��,���Ͼ6�����>4��mF�)�Q��U��Q�9�D�B[2�r��o� �|˾v��<�T�ݭ�`؞� B*��ݼR��u����
��p�+�����XVH�Q/��(ᨿ�3Ϳ���TF��Z����w��p�.[�H ����T�˿�����z��`�G����C��<�q���{���h�� ���5��ॽ�   �   r9��|����&?�j+��������Ͼ=����V�����qJ���r\��̾�U��h��A�9��j|�������[�`i��-�d�����0��З���V�/�"�s�ޠ���ʿu���j�"��51�;�x3>��[:�� 0�� ��d�� ���ɿK�����s��0���0���j3�.F��x�&�Ԙ��,i���g��   �   ����� d�Qnɽ���L�����ؖ��稾�K��(跾�d���9��V�����z��F�n�� .����P�.��`�;`J�; �λ�/��ݽ��V�hy���)��;O��������������Y&��=�x�O�؈\���`��[�B�N��<�n�%�ֆ��k꿽)�� ���HP� >�1����Z���J:>�`�"��Ee; ���   �   ��a<�л��&&��>�ӽ~q���,�>�E��2U�8Z��S���B�BH)��	�z�ʽ�������@�����<d��<d��< ���CI�6��8�y���Ѿ)F"�L�j��Ġ�^�ѿ�R�� �"n;���V�ȿm�l}��f���|�Fm�>�U�� ;�.�����ҿx�����l���#��Ծ0�~��V�fpZ�0'ǻx�<E�<�   �   p�=4{�< /<�t�`�#�G�����GӽF����潦�ν�-��v�x������,��>P<� =x	/=�Z3=�<  �68}a�~g�f�����羥2��A��+Ѯ�4^�>S�h�,�D�L�� l����>����������x��|l��M�Ή-�,�A�QW��˒��eL4�of���� ��&�t�0I���]�<nt!=�   �   ��V=��<=lu=��{<�J~�������!��[W��x��F���6t�@ O��D�pB��  �7�C�<�L=<�N=�i=��Z=�>=��C:��r��������$���L7<��!��[�������d���5�HkX���z��H��݄���#������U���{�t<Y��7�؏�{��������D�>���������w!�H}���R����=x?H=�   �   �P�=D?s=�;I=DP=t/�<��;pb�Dq���/м��ݼ�=ļ l�� ���`�<`��<�~*=e=*	�=��=G��=2�J=Le�<���>���J{���վ�g%�Feo�7����bտ���j"�8*?�l[���s�]<���5���A��� t���[�@�b&#����׿�˥��r��Y(��ھx����c��I;��<N�-=r=�   �   ��s=�[\=��+=���<3<��񻀏��̞	��S&��$.�R> �����0R������x<�=��G=�y=_�=hف=��D=��<��;�����u�=NѾ�W"��5k�������ѿ�}�N`���;�XW���n����f�� ��o��W�6�<�Z ����ԿV�X�n��$%�1־�~��	��b5��<��'=6�f=�   �   @=�H=�"�<����̺�6��D��.���؋��A�SP������s�Φ ��։�`��;ܿ�<�2=�p\=�A`=�21= r}<��	�_��`f�ž_o�o_������ǿ��������j2���K��Oa���o�� u�ܯo�Na��K��2�"S�e%��ٖɿ����P�a�#���4ɾ��m����<�$��<@�=�JD=�   �   h�<p��;d���mC�������3��!�,3/�&:3�e-�9G��N�I+ս5:���(�p}8���b<��=0u"=&u=��]<����ǽy�M�B籾����K�Ȋ��E���Y翎���$�dp:��M�̐Y���]��%Y�b{L�J�9��#�Z���翮'����t�M�nV��G����S�s�ӽr ��@�; ��<6�=�   �   P��v���똽���.�'��7U���}��������������x������/ x�;�N��� �9{�ȹ���v�� <l��C�<��<�<����y��O/��љ�͠�kb3��x�A��H�ο����6��o%�R5��G?�|�B��>�.4�ą$�R���R���Zο�3����y�ۀ4����:A��P04�df���+缰��;�̓< j8<�   �   ��R�Vƽ�]���\��O���5��-oξ�U�8��B8���g�����"˾%l���Y���)U��
��ݸ��4:��5_���F;@�;4���H������2�}���˾Ә�<T����j"��:ؿ�������z�V�#��]&��"#������N�����ֿ�O��o]��]T�����̾�k��~J�p��w���I����8����   �   �߽3�3������r��uC�oQ�l����+�#�5�(9�$5��X*������۾A)���}�h-�%$Խ��]�p���������HFF�$ٽ=�F�Ĭ���O���r-�Q$h���f��7Rӿ�t�����y�*�
����� �YI�Fѿ�����m�f�ͮ,�:����Ǣ�:H�<�ܽ��O�������R���׼�,q��   �   R�9��b����ľ����^"���A���]��"s��P���n��F���q���Z��
?��������k���#.��N�4�}׽p-a�Ԭּ\D���b��������v�)��ٍ�oe7�~�k�=���8D��=�����ѿm�ܿS���ۿSп-����W�����%)i���5�%U�����M�t�	�����s��������m���߽�   �   ɢ��&Iɾ�
��z3��,^�򋃿_z��=_��g	������YP��<��ܓ��ށ�i[�|�0����Sƾd���x+��ýҐF���Ѽ�zԼ��J���ƽ.����)Dɾ�
�w3�T(^�^����w��E\��_������uM������ٓ��܁��[���0���}Pƾ����8+��ý��F�H�Ѽ��Լ8�J�i�ƽ�	.��   �   z�����i7���k�µ��G��Q����ѿ��ܿ����ۿ�Uп˯���Y��~
��R,i��5�W�K����t�.	�#����s����(�鼎�m��y߽�9�m^��n�ľ����Z"�`�A���]��s�*N��Pl��4��q���Z��?�Ԯ�����n���*+���4��w׽('a���ּ0H���h�(	��؏��v��   �   LT���u-�&(h���Ui��0Uӿ)x���{��
�d���� �	L�\Hѿ���9Ē���f���,������ɢ�sH�l�ܽ:�O�$���زR�(�׼�q��u߽x�3�E���;m��&=��M�n��Z�+���5��#9��5��T*�j�����۾%��^�}���,�BԽ��]��y��X������MF�jٽ�F�6����   �   D��` T������$���<ؿ���`���|�(�#��_&�X$#���J��������ֿQ���^��&T�Q��w�̾�l���K�����r��@�� ������R��Kƽ�V���\�K��d0���hξ�N�]��i1���`����@˾Qg���U���"U���;ָ��):��_��1G;��;���Y���H��F�}�y�˾�   �   �d3�!�x���y�οG ��:8�Rq%�5��I?�D�B���>��/4��$�V��UT��I\ο�4���y��4��	��	B��14��f��p(�`��;`ڃ<h�8<�4����ᘽo���'��/U���}��������������s����� x��N��� ��q�.���4`���Cj�M�<��<��<��/~��xR/��ԙ�^���   �   ��K�'����F���[翰���	$��q:��M�z�Y�R�]�
'Y��|L�V�9���#������e(��D���$�M��V�H���S�C�ӽ���[�; ��<
 =P/�<`L�;����\C����!����]�!�>,/�?33�X^-��@��H�!ս�1���(�PS8��c<��=*x"=�u=8�]<x��E�ǽ��M��鱾����   �   I_����1 ȿL�������k2���K��Pa�F�o��u���o�<a���K���2��S��%��.�ɿǖ����a�8���4ɾ��m�����$� �<"�=pOD=: @=�P=L5�<���h����6��<��ȯ��5����丽H��\��
s��� ������;���<r�2=�s\=C`=�21=�h}<��	�3��Ff�"ž�p��   �   <7k�Z ����ѿ~��`�r�;��XW���n����f����	o�T�W�X�<�Z ����Կ0��n�x$%��־�~����_5��'<��'=��f=��s=.`\=��+=���<�M<�������	�zK&��.�~6 �����dE������x<��=r�G=ty=f_�=Lف=t�D=L�<^��y���4�u��OѾ�X"��   �   (fo�����cտ���"��*?�Nl[���s�m<���5���A��b t�~�[��@�&#����N�׿5˥�3�r�<Y(��~ھ�Gb��E;�H"<��-=�r=TQ�=�@s=�<I=`Q=�1�<p�;H_�p��/м��ݼP>ļ�l��� �<t��<�}*=�e=��=��=o��= �J=�_�<b���@���L{���վ|h%��   �   ,6k�������ѿ�}�F`���;��WW�`�n�,�+f��R��o�F�W�z�<�ZY �b���Կx좿�n��#%�|־~���4]5�8/<��'=B�f=,�s=�`\=4�+=Ԝ�< N<�������	��K&��.��6 ������E�� ����x<��=|�G=�y=�_�=�ف=~�D=��<Ж�������u��NѾ�W"��   �   @_�i����ǿ@���x��nj2��K��Na���o�D�t���o��a���K��2�2R��#��s�ɿf���l�a�����2ɾ��m�����$���<N�=�PD=*!@=0Q=6�< ������6��<��֯��I����丽-H��x��2
s�� ������;���<ԥ2=�t\=DD`=t41=0u}<��	�s��pf�žKo��   �   ��K�M���qD���X�����$�`o:��M�P�Y�
�]��#Y��yL���9���#�4�����%��[���7�M��T�
E����S�ݵӽv�`��;4��<
=�1�<�S�;����&\C��������d�!�N,/�N33�j^-�A��H��!ս2���(��R8��c<��=�y"=~x=x�]< ���ǽ̧M��汾����   �   da3���x�K��	�ο)���5�~n%��5�F?���B��>�Z,4�&�$����#P���Xο2����y�j~4����~>��J,4�9`��T�0��;��<��8<p(����ᘽ<����'��/U���}�明����������s�����x�1�N�ʯ ��q����,_�� �i��P�<�<��<�����w���M/�љ�i���   �   ���|T�෌�� ��88ؿ˸��h��Fy���#�0\&�� #��~�R��S���E�ֿ;M��z[��.
T�����̾i��VF����P`�� ���$�ۛ�N�R�Kƽ�V���\�K��a0���hξ�N�e��t1��a����L˾Zg���U���"U����ո��(:�H_��jG;��;t�������8����}��˾�   �   �L���p-��!h��쓿�d���Oӿ9r�V��Rx�p�
����N� �!F�Cѿ{���S�����f���,�l���Ģ��
H���ܽ$�O�\w���R� �׼Fq��t߽3�3�0���-m��=��M�n��^�+���5��#9��5��T*�q�����۾%��V�}�h�,��Խֵ]��r��P������?F�6ٽ��F�ת���   �   j������b7�R�k�K����A��������ѿG�ܿ�}�ۿ�Oп"����T�����$i��5�HR�2����t���1���df����H�鼪�m��x߽��9�M^��Z�ľ����Z"�^�A���]��s�-N��Tl��:�q���Z��?�ٮ�����m���+����4��v׽�#a���ּ$7���[�i�������v��   �   t����@ɾ;
�t3��$^�:���u���Y��{������tJ������֓�Dځ�P[���0�m�vKƾ}��I+��ý�~F�ЌѼjԼ:�J�"�ƽ�.�ڞ��Dɾ�
��v3�P(^�^����w��G\��a������xM������ٓ��܁��[���0���tPƾր���+�Dý��F���Ѽ�lԼv�J���ƽn .��   �   ~�9�\[��a�ľ���W"���A�u�]��s��K���i���y��q���Z�v?����������&����4�\m׽�a���ּ�.���[�5���Cv���͍�he7�y�k�:���8D��=�����ѿn�ܿU���ۿSп0����W�����*)i���5�"U�������t�d�����m�Ĩ���~�m�6s߽�   �   n߽`�3����h���7ྶJ����j�+���5�S9�p5��P*�}��^���۾���Ϫ}���,�xԽ�]� ^��(k����D@F�.ٽ��F�����|O���r-�J$h���f��6Rӿ�t�����y�,�
����� �[I�Fѿ"�����n�f�̮,�.����Ǣ��H�x�ܽ��O�,~���R�8׼�q��   �   җR�tCƽ�Q��\��F���+��lcξ�H�̬�*��6Z�I��,˾�a��$Q���U�,���˸��:�(�^���G;�K;Ģ��⩃�(����}���˾ɘ�6T����i"��:ؿ�������z�V�#��]&��"#�������R�����ֿ�O��q]��^T�
����̾�k���I�5���h�����@��Λ��   �   ���j|�ژ������'��(U�d�}�Z�����������n��?���x��N��� ��e�@����?����f�8c�<��<�<����x��|N/��љ����cb3��x�@��H�ο����6��o%�R5��G?�~�B��>�.4�ƅ$�T���R���Zο�3����y�ۀ4�v��A���/4��d��0!��Ӊ;��<�8<�   �    <�<���;(铼�NC��	��O��R�.�!��%/�p,3��W-�m:��B�`ս'(����'��8�H5c<��=��"=~}=�]< ��ϔǽ�M�%籾����K�Ɗ��E���Y翐���$�dp:��M�ΐY���]��%Y�d{L�J�9��#�\���翱'��Ĉ��v�M�lV�~G��Y�S�F�ӽ�� o�;���<�=�   �   �#@=�U=�B�< ��螺��6��5��5���{��Iܸ��?��6w����r��� �|���@"�;D��<h�2=�z\=(I`=X81=`�}<b�	����$f��ž[o�n_������ǿ��������j2���K��Oa���o�� u�ޯo�Na��K��2�"S�g%��ږɿ����P�a�"���4ɾ��m�"����$��<��=�QD=�   �   ��s=�a\=��+=���<0_< ��$s����	��C&��.�p. �����06�� 4���x<V�=��G=�y=ia�=8ہ=R�D=H�<ܓ�������u�5NѾ�W"��5k������ѿ�}�N`���;� XW���n����f����o��W�6�<�Z ����ԿV�Y�n��$%�-־�~�x	��a5��#<l�'=��f=�   �   /}�=��=�j=�9=�0=�˟<@�< u�������_ѻ`\V�`�w;x^h<(��<��(=�&c=*��=ȑ�=�s�=N�=M�=�V
=8�c�!尽��C��㬾}��H�m���/�����J�	��t!���7��J���V�~[��V�8JJ�4 8�%"���
���4�����efK�	���f���jN��Ž@Ǽ�<cR=A��=�   �   �A�=�Qz=^�P=L�=X��<��<��U�(�P��햼0:��0���ؖ��a,;l��<~�=Z�C=Pl}=�x�=��=�0�=|
{=*�	=@8R�t���OT?��N��8���kD������9��1�߿<�����q4��zF�8�R�L�V��R���F��4��^��S���Ῐ��9z����G�������twI��Ͽ��h����<*�M=Ł=�   �   �@b=�>=�n=`m<�
�����TS��9R��q���x�lrh��_A�j����y��;4��<��.=$Ck=z�=��=�i=�P=�o!��g��� 2��잾>����9��ۀ�t����fտ�.�V2��m+��<�v5G�pK�G��;�,d+�&h������ֿV���vB����<�3� �8��� 5;����䦞��e�<�w>=4/f=�   �   \�=���< <.��ռ�,X��,��  н�T��
Z�fo�{��뽦~ý"�����3� u��HV<�� =�a@=P�\=�J=�T�< ^��/c��r��Ď�����)�rl�󛿇�Ŀ"o�0g�����x,��*6��p9�*�5�L ,�@��1�ą�jCſ����?�m�~+�4�������@%�=�����g� ��<*#=��2=�   �   ��<�����4I�I���� �d�&���H�=hc���s��x���q�B�^� B��~�q��윽�� �� ݻ`k�<
�=*F=�s�< ֪��S�1��|�t���ƾ��ubP�_d��JO��c�Կ����b���U�t�!�b@$��!!���V��M����CԿg ��?���8Q������ɾ�jz�M�	�p�m��x���<�1�<���<�   �   �\켖��O��io-���f�X������t��M�Ǿ�B˾\)ƾ�Ƹ�Xh������}\]���#�vٽ�p�㥼 
�;�x�< �<�;r���2Ͻ�SG��)��U�����0�N�l�����Q����(׿���RI�h'��Z�F�
�ȁ�*���տ\}��C��k���0�\����s��w�J�,�׽*�,��es�(se<�g<��\��   �   �ɟ���	��O������\����޾q� ����%���-?�x��ex����پ�C��B����LF��n��c��8g漀 S�H�%<@�I;4�üƙ������O����Ⱦ����B�\y�s����n����ʿ#ݿ��S�T�翵�ۿ�ɿ8���m+��}�v���@�m��^Ⱦ�j���:����ݼ�J�� �;`ٻ����   �   ,����_�"퟾�Nվ/r�!T!� 9�y�K�40W���Z�F%V���I�*�6�o��L��R2оm���'X�au��%��LT�����@g�:��S�0D��ؽ�uA�J ����޾0P��=E��}s��ݏ��;���<��(���뇾�"Ӻ��۰�����B#���hp�9�B��u��NܾpT����?�\Y׽��E���i�@ũ� ��	��ߞ��   �   ��Z�Җ���l���t�9���\��{�g剿�e��C���?���G����x�Y�Y���6�q��2߾5E����U��� ������ƼP���0����Ӽ؈��U�+�Z�����Cg㾠���9��\�>�{��≿!c����������򷈿��x���Y���6��n��.߾EB��t�U�ę �ʬ��X�Ƽ ���`ૻ Ӽqވ�QZ��   �   �����޾BS�zAE�߁s��ߏ�m>���?����������պ�dް�����?%��lp���B��w��Qܾ�V��̒?�]׽*�E���i��]����
v	��מ������_��蟾Iվ�n�WP!��9��K��+W�H�Z�� V�w�I�|�6�<������-о�i���"X��q�� ��\I�@ꚻ@3�:��S��9D�|�ؽ�zA��   �   ��Ⱦ���DB�Uy�����Xq��x�ʿݿ���F�%��N�ۿAɿ=���#-��H�v��@����ȾCl��� ��;��̾ݼ ��J�;�ػ�|������	�áO����.W����޾� ���c�R���;���Wr��a�پ#?�������FF�Zj��]���W� R�X�%< �I;��ü(������R���   �   �����0���l���������O+׿���J��(�@\���
���m��տ�~�����k�(�0�����u��<�J���׽��,� Is�8�e< �g<�(Z�PA켡������th-�N�f�FS��{��/o��v�Ǿ=˾�#ƾ^����c���򊾒U]���#�]mٽ��p�xХ� 9�;0~�<��<��;h��;8Ͻ,XG��,���   �   ��eP��e��0Q����Կ3 �����PW��!��A$��"!���^�����@EԿ�!�����J9Q�����ɾ3lz���	���m��r�Р�<�<�<(��<��<`Ň��#I������ �b�&��H��_c��s���x�?|q���^�B��x�/��V䜽^� �0�ܻ y�<0�=�G=xq�<�Q��S�����t���ƾ�   �   �)��l�|���7�Ŀq�Dh�ܫ�(z,��+6�2r9�V�5�N,��@�n2�ن�>DſO���!�m��~+����Z���A%������g�Ե�<r#=��2=�=h��<�-+���Լ�X��"��>�ϽJI��T�i���U���tý�~��J�3��]���z<�� =rf@=�\=��J=`Q�<�~���f���t��Ǝ�����   �   ��9��܀������gտ�/�23��n+��<�x6G�fK��G���;��d+��h������ֿ�����B��ס<�F� �4����4;�;������k�<�z>=|3f=
Fb=\>=�v=`4m<P���(l���E�6+R��	q�
�x�:dh��RA�r��Yy���;x��<h/="Gk=��=���=��i=�N=�!�Fk��l2�\�����   �   ,mD�U����:��*�߿Č�>���q4��{F�КR���V���R��F��4��^��S���῀��z��X�G����z����vI�Xο��c����<ʘM=sƁ=�C�=�Uz=��P=f�=ܙ�<��<�KU�p�P�lߖ� ,���煼 ~� �,;̜�<`�=f�C=�n}=�y�=L�=�0�=X	{=�	=�FR�=���TV?�:P��)���   �   oH����	0��*�㿌�	��t!��7��J�؟V�~[�̧V�JJ���7��$"�V�
���志3�������eK�g���e��$iN��Ž��Ƽ��<eR=��=�}�=C�= j=�9=�1=|͟<�< 3��ྮ��^ѻ _V��w;X\h<Ď�<��(=�%c=���=3��=�r�=LM�=)L�=PT
=��c�A簽��C�w䬾�}��   �   AlD������9��?�߿6������p4��zF�ΙR���V�x�R���F�J�4�(^��R���ῷ��yy��d�G�������JuI��̿�_�����<�M=�Ɓ=�C�=0Vz= �P=��=8��<��< KU���P��ߖ�,���煼p~� �,;���<\�=f�C=�n}=�y�=~�=1�=B
{=F�	= >R�����U?�JO��}���   �   ��9��ۀ�0���"fտv.��1�tm+�<��4G�|K�G��;�6c+�Dg���%�ֿ ���rA���<��� �Y���>2;����ę��Tq�<�|>=�4f=�Fb=>=@w=�5m<𯐻�k���E�B+R��	q�$�x�^dh��RA����xYy��;���<�/=xGk=�=��=B�i=ZQ=�n!�h��� 2��잾����   �   ~�)��l�w���Ŀnf�ީ��w,�`)6��o9���5��+��>��0�уAſ8�����m� |+�F��ʗ���=%�\���0�g�x��<`#=��2=j�=`��< +�t�ԼpX��"��1�ϽII��"T��i���p��uý�~��f�3��]���{<2� =Zg@=V�\=�J=�X�<�O��Fb��rq�!Ď����   �   -��7aP��c��5N���Կ���`���T�"�!��>$� !�����������AԿ{������X5Q�����}ɾfz���	���m�pT�(��<�C�<���<8�<Ç� #I������ �T�&�
�H��_c�(�s���x�O|q���^�,B��x�G��Y䜽@� �`�ܻ{�<��=�J=�z�<�p��Z	S�����t�q�ƾ�   �   -���{�0�M�l�_��������&׿w��H�&�HY�į
�N��a�m�տ{��@앿V�k��0����ep����J��׽��,���r���e<H�g< �Y��=�������Lh-�.�f�?S��w��0o��z�Ǿ=˾�#ƾf����c���򊾞U]���#�Emٽx�p�TΥ�pH�;���<��<��;�~��/Ͻ�QG�b(���   �   G�ȾX���B��y������l��Z�ʿ�ݿ�|�^�W��ɋۿ(ɿ����")����v�h�@����=Ⱦ�g��X��2���ݼ �}��w�;�ػdz�(�����	���O��W����޾� ���d�V���;�!��`r��j�پ(?�������FF�:j�]���S� MQ���%<�%J;��üT������BN���   �   ������޾N�;E�'zs��ۏ�y9��@:��p������Fк�ٰ����� ��jdp���B��r��Iܾ�P����?��P׽ʟE��i� Y�� ��br	��֞�f��t�_�|蟾
Iվ�n�RP!��9��K��+W�L�Z�� V�|�I���6�A������-о�i���"X��q����\C�PÚ��"�:(�S��(D�<�ؽ@rA��   �   ƹZ�����Kc��l�9�f�\� �{�~����`�����$���h���	�x�J�Y���6�7k�X)߾�=��˨U��� �Ȥ��,�Ƽ�4�������ӼUֈ�U�нZ�w���.g㾘���9��\�<�{��≿#c������¾��������x���Y���6��n��.߾<B��A�U�d� �m�����Ƽ@[������(�ҼQӈ�xR��   �   ���~�_�!埾�Dվ$l�M!�@9��K�C'W���Z�^V��I�]�6�~��T��k(о.e���X�l����-� ��� ��:p�S��+D���ؽ&uA�" ����޾'P��=E�}s�ݏ��;���<��)���쇾�#Ӻ��۰�����E#���hp�;�B��u��Nܾ[T��n�?�5X׽ީE�ȸi� ������zm	�'Ҟ��   �   p���w�	��O�^����R��h�޾�� ����������7�����k��P�پ�9��8����?F�vd�>T���9� O���%<�SJ;4�ü󗖽V���O����Ⱦ���B�Xy�r����n����ʿ%ݿ��T�V�翸�ۿ�ɿ:���o+����v���@�n��QȾ�j�����8����ݼ �~��y�;0�ػ$s��   �   �+켜���콼b-�O�f� O������i��܇Ǿ=7˾�ƾͻ��p^���튾qM]��#��aٽl�p�����`��;$��<�$�<�;�1ϽfSG��)��?�����0�H�l�����O����(׿���RI�j'��Z�F�
�ȁ�,��տ^}��E��k���0�W����s�� �J���׽6�,�@s�(�e<��g<�'X��   �   0�<���I�\}��� �D�&��H�=Xc���s��x��sq�_�^��B�r� ��ڜ�>� ��@ܻd��<��=NP=��<�5��v	S����#�t���ƾ��pbP�]d��KO��c�Կ����b���U�t�!�d@$��!!���X��O����CԿi ��A���8Q����րɾ�jz���	�v�m��e�<��<F�<l��<�   �   ��=`��<��(���ԼnX�w����Ͻ�>��zN��c��
�}�|jý*u��d�3��@���<� =o@=^�\=|�J=$_�<@A��b���q�xĎ����	�)�nl�󛿇�Ŀ"o�0g�����x,��*6��p9�.�5�N ,�@��1�ǅ�kCſ����B�m�~+�/��♒�h@%�5���p�g�H��<x#=��2=�   �   TIb=�>=�|=�Qm<`k��XW���9� R���p���x��Uh��DA�4��H(y� >�;t��<�/=&Nk=��=H��=��i=
T=Xf!�Bg��� 2��잾2����9��ۀ�s����fտ�.�T2��m+��<�v5G�rK�G��;�.d+�&h������ֿY���vB����<�2� �,����4;�M�������l�<<|>=�5f=�   �   D�=fWz=.�P=z�=���< �<`�T�h�P�hҖ�8���م��b��#-;0��<��=f�C=�r}=�{�=�=�2�=�{=ڃ	=x3R����4T?��N��5���kD������9��3�߿<�����q4��zF�8�R�L�V��R���F��4��^��S���Ῑ��9z����G���򛮾^wI�tϿ��f����<��M=�Ɓ=�   �   �<�=v$�=*��=��Z=��0=��=�s�<�G�< �q<0�n< E�<���<�,
=X�8=*�k=`I�=�٥=)a�=�9�=�>�=/��=�jT=�"=<j�I�3������~D־���jX_�����=����Z7�J\$�`�-�l�0��-��y$����D�eE�ꑼ������b���"�S�ܾ`$���S�D_������P�=
�m=�ʎ=�   �   m^�=��=�tl=��@=*�=T�<H�t<Pj�;`�y; �b;���;�d<L��<
�=�}L=o��=$�=���=���=�̱=��=̀S=�	K<��@�8���̀���Ѿc���g[��p��4���=P߿���T����!�@�*�t�-�N�*�d�!�H���6v��\��^��r^����ؾ� ��.��z���K�*3=��i=��=�   �    �z=��\=
�,=���<XO< ����p� )Ǽ�����.��8�ۼ�����"���G<��<d�2=2s=�V�=��=�0�=�o�=B-P=Hhq<v](�H��S�p�`�ž�$��O�<)������Կ����|����N'"��%�b"���l���A��Bhտ�
��N���cR����\�ʾN�{�*8	�4�]� �k9��=Б^=֣~=�   �   �X<=�=Pww< ���S༆�E��b��<���R���6��i;������wm�pK�p�g�H�<� =6�K=��=���=�Մ=��H=�F�<^-���ؽ�`V��<��
��p�=�@d}��
���ĿX��h���}����������*��d��M��"Ŀ�s����~���?�|��_����_�`��$2�`��; �=��I=��U=�   �   �1�<��;��ʼjIb�~�����P���B)�	Y6�u�9�O3��J#�J?�_�ڽ�G���)��a"�@��<P:=|�S=�5`=�':=$�<����#���,5�Ȱ��n��(�&��_����������̿�t��X��J�����x��|`���j���˿���6Վ��D`���'�1����<������(�(<�M=n4(="=�   �   �8�Q#�x�������4c-�O�Z�W����+��蚾G���3V����{Lz��P� !�0?�����)ؼP�;�s�<R�%=�y!=�+�<p��4����0|���þ��_Z>�\�t�����Pz����ǿ}�ٿ!/忷�����ؿ;`ƿ_@�����FOs���=�~����ľ���^����ؗ��@�t<@8�<4��<(Ą<�   �   ��B�����@�_Z�P?��#t���˾OV�wL�܇�l���޾}ƾ9��I��F�M�o��������K���_�<XT�<���<��:?&�.Խ�AC�����
�"�7�H�j�w�Am���'���y������¿�f��_K�����K ��.cu���F����Hx��욾oC��{׽��2��e�P��<�R�<� K< �:��   �   �XȽ��&��u�^���NԾ> �����#�^�,��/�ָ+�tM!�c������tξ����]	k�x���������PK��%�<�-�<��<�ۡ������l��Ai����i�����>D�-i��҄�p���T���ћ�Y���kR��Vj��Y8f�.~A��{����1I��9@e�Z�	��������� ��;@ϕ<��I<��z�=��   �   "��R{����.�fD�bj1��%K��2_���k�
�o���j�Y/]�Z�H�&�.��d���Zs��ns�����ઽ�7� ��9��<`�<����������"��K{�P���(�+A��f1��!K��._��k���o�j�j�q+]�׀H��.�b����p��2is�=���۪�2� Ƶ9��<��<����j(�?���   �   �Gi��"��n�����BD�+1i��Ԅ�jr��W��-ԛ������T��@l���;f���A�
~�:���K���Ce���	�ѡ���������;xԕ<��I<�����=�PȽ�&���u�ɱ���HԾ�: �����#���,�<�/�4�+�J!� `�J���Qpξ$��k�D�򒶽h�� K� )�<+�<X�<�롼����%q��   �   ʟ��h��$���H�D�w�ko��1*��|��d��o"¿*i���M������ ��fu���F�����z���qC�׽�2��e���<�[�<p=K<8�:�L�B������:��Z��:��o���ʾPP�DFﾯ��x��8޾xƾ���vE��^�M�����橽��� y��g�<�U�<���<@a�:�G&��4Խ�FC��   �   C�þC��,]>���t����w|��ڵǿ��ٿ�1�'��c��?�ؿbƿB�����yQs�y�=�±�h�ľD�`�����<�����t<$?�<���<�Ԅ<����B#����v���n\-���Z�|��M'��3㚾|����Q������Dz���O�j!��5⽦�ؼ�)�;�}�<%=�y!=&�<����8����5|��   �   ���U�&���_�u���f��� �̿,w�[��r��������ib��zl�d ̿ ��(֎�F`���'������/<�G��������(<�P=�8(=�=0C�<`p;��ʼN8b�e
��5������;)��Q6�f�9�DH3�;D#��9�N�ڽ?�� �(�6"��ʎ<@=�S=\7`=�&:=��<�����'��Y05�G����   �   ���j�=��f}�����Ŀ��\���~��������h+�Je�O��#Ŀ�t����~�]�?��|��`��4�_����#2�p��;L�=t�I=T�U=�^<=�=ȟw<л��$7�`�E��Y�����%I��+-���1������gm�h=��Pg�H�<� =��K=�=դ�=�Մ=��H=@�<P3���ؽ<dV��>���   �   �%���O�:*����W�Կ-���<��ְ�("�z%�"�x��ީ�aB���hտA��VN��dR�ӯ�z�ʾI�{��7	��]� 2m9��=��^=\�~=��z=z�\=Đ,=p�<X<O<`� �8�p��Ǽ8��������ۼ�╼�Ҿ��j<|,�<h�2=�s=@X�=��=01�=�o�=�+P=�Zq<�b(��L��9�p�`�ž�   �   b���h[��q�����Q߿$����� �!���*���-���*���!�n���Gv��\��K񒿑r^�y���ؾ4 ��n-���z�@mK�B5=4�i=�=�_�=�=�xl=��@=�='�<8u<P��;��y; Xc; *�;� d<���<��=4�L=���=�=$��=ɺ�=�̱=p�=�~S=@�J<��@�����΀�Ҿ�   �   ;��'Y_�3�b�����<���7�j\$�t�-�l�0��-��y$�r���C��D�{��������b�W�"�H�ܾ�#��mR�i]�����p�=΅m=�ˎ=}=�=	%�=���=��Z=��0=\�=4u�<�H�<@�q<��n<�D�<<��<z,
=��8=r�k=�H�=~٥=�`�=�8�=N>�=a��=�hT==< �I�i��z����E־�   �   ����g[��p��?���3P߿���0��N�!��*��-�ܭ*��!������Qu�\���𒿄q^����sؾe���N,���z��KK��6=R�i=o�=`�=��=yl=* A=L�=\'�<�u<К�; �y;@Xc; *�;� d<���<��=.�L=���=�=:��=꺶=ͱ=��= �S=�K<��@����΀���Ѿ�   �   n$���O�)�������Կ ���������&"�
%��
"�$�����C@���fտ�	��M��bR�Q��G�ʾ3�{��5	�*�]� Dq9��=��^=ܨ~=��z=T�\=r�,=��<8>O<�� �x�p��Ǽ��������ۼ�╼ Ӿ�hj<t,�<r�2=s=fX�=��=�1�=~p�=�-P= iq<~](��H��F�p�C�ž�   �   �����=�Ec}��	��ĿE�忾��$}���������)��c�0L�?!Ŀ[r��	�~���?�vz�{]���_� ���2� Ҥ;B�=T�I=f�U=t`<=�=��w<@����5���E��Y�����I��+-���1������gm�~=�Qg���<� =R�K=p�=z��=�ք=�H=�I�<�+���ؽ!`V�<���   �   ���!�&���_�����l�����̿Ts��V��:��z��P��/^���h���˿����ӎ��A`�_�'���y���<�6y��x����(<xU=H<(=
=�F�<��;��ʼv7b�

���������;)��Q6�j�9�LH3�GD#��9�_�ڽ?����(�X5"��ˎ<A=��S=�9`=�*:=�$�<�z��#!��v+5�̯���   �   �þȽ��X>�2�t������x����ǿ_�ٿ�,�I�还�俰�ؿ�]ƿ7>������Ks���=�6���ľ���Z�諌�새�`�t<�I�<�< ڄ<���<A#���� ���<\-�a�Z��{��G'��2㚾~����Q������Dz��O�p!��5⽐�ؼ�1�;4��<��%=�}!=(3�<��w1����R.|��   �   ����f�O ���H���w��k���%��mw�����~¿Md���H������#���U_u�G�F����s�z难�iC�t׽��2�@cd�4��<Lf�<�LK<h�:�H�B�ȭ���:��Z��:��o���ʾLP�DFﾲ��|��A޾xƾ���yE��]�M�����橽��� D���l�<�^�<���<���:9&�*Խ8?C��   �   �=i�&���e���<D��)i��Є��m��[R��gϛ�򳘿P��h��F4f��zA��x����%E���9e���	�E����|��H <�<�I<��=�*OȽ��&�a�u������HԾ�: �~���#���,�A�/�6�+�J!�`�Q���Vpξ&򠾹k�,�~���ܬ���J��1�<�7�<0 <ϡ�n����i��   �   ("��F{���u$쾕>��c1�/K��*_��k�Q�o�
�j�0']��|H�p}.��^�v�澢k��bs����`Ӫ�l$� h�9%�<P�<@4����z��n"��K{�2���(�!A��f1��!K��._��k���o�n�j�v+]�܀H��.�b����p�� is���R۪��/� ��9��<@�<� ����2���   �   �IȽ��&���u�!���!DԾ@8 �r��q#��,�{�/�n�+�kF!��\�����jξ��9�j�@�u���l��@CJ�>�<�>�<�	 <�ӡ�)���Ll�.Ai�����h�����>D�-i��҄�p���T���ћ�[���mR��Xj��^8f�2~A��{����*I��@e��	�����$���� <�ޕ<h�I<����w=��   �   �B�&���6���Y�67���j���ʾ�J�Q@ﾇ{�Q��I
޾�rƾ����A����M�����ܩ����⳺4|�<�h�<$��<���:�;&��,Խ�AC�^����	�"�0�H�d�w�@m���'���y������¿�f��bK�����M ��3cu���F����Ex��욾�nC�{׽�2���d����<Hf�<�WK<8�:��   �   ����6#��x�������V-���Z�x���"���ޚ������L��&��$<z�>�O��!�d*�ꆽ��׼���;��<Ƥ%=�!=,7�<@���2����0|���þ���YZ>�W�t�����Oz����ǿ}�ٿ!/忹����"�ؿ=`ƿb@�����HOs���=�}����ľ��D^�����쐈�p�t< H�<|�<��<�   �   LQ�<�;��ʼ�)b������&���5)�.K6�f�9�FA3�|=#�83���ڽ5����(��!���<J=|�S=�>`=.:=,(�<�z���!��x,5�����\��"�&��_����������̿�t��X��J�����z��`���j���˿���7Վ��D`���'�.�����<�Y~��������(<
T==(=�=�   �   �c<=B=��w<Pj����8�E��Q������?��}#��E(��d��
Vm�^-�g���<' =�L=��=��=�؄=��H=HM�< +�7�ؽ�`V��<����j�=�=d}��
���ĿY��h���}����������*��d��M��"Ŀ�s����~���?�|��_��h�_�׉�J"2� ��;^�=2�I=��U=�   �   ��z=Z�\=ȕ,= �<`ZO<�k �xlp��Ƽܑ������T�ۼ˕��y��ȓ<�>�<|�2=� s=G[�=J�=�3�=r�=B0P=�pq<\(�	H��(�p�Q�ž�$��O�;)������Կ����|����N'"��%�d"���l���A��Dhտ�
��N���cR����W�ʾ:�{�8	��]� pm9d�=�^=d�~=�   �   4`�=-�=�zl=�A=D�=�.�<�&u<���;@Tz;`�c;0Y�;�7d<���<:=��L=� �= �=ֺ�=T��=Pα=��=X�S=�K<N�@����̀�~�Ѿ`���g[��p��7���=P߿���T����!�@�*�v�-�P�*�f�!�H���7v��\��^��r^����ؾ� ��.���z� �K��4=
�i=3�=�   �   �V�=�Ȍ=C�=�1i=�/L=z�0=��=�=��=Z�
=�e=xo4=ZW=�\�=-��=��='�=���=j��=���=gl�=�~�=R�=�[��
��/=9�������l,�`Bg�����0���vӿ�8ￆ���	�L6���	�ڳ���ￅ!Կ���ٵ����i��Q/��������@�I�6�ҽ����7<,W*=.it=쉌=�   �   H��=��=^;t=��T=��3=��=���<DV�<�a�<4��<���<Hr=V�6=lRc=���=���= Ķ=���=pP�=�$�=0A�=���=*,=�A��5��/�4��$�����FA)��2c�6��k7��4пPX��~ �z�t�	��w��� ����r�пJ�������e���+�i������D���˽����J<8�+=�Wr=��=�   �   (=0g=�YB=v�=���<P�w<P�; ���\Y� 
:�@��:�b<�<\R	=l�D=R�=��=���=���=|��=�=&3�=0=Pt��V��Vt'�#b��$��	 ��]W��ŉ�����ƿ��u����� �B(��� �^w���Z<ƿG������\>Y��E"�x]徦���B6�{���h�ݼ�<Hr.=�k=���=�   �   <P=(6%=X��<��)<p/ɻxt���R��K9���O���Q�̱=�����������@Uq<><=��V=�ӊ=P��=�~�=��=cb�=`j'= |@���v����j&��a�ʾ'����D���|��皿E��Bcο�Qῴa��m��E�࿴�Ϳ�������AB}�Y�E��#���ξ�����C������ 3�<�1=�\^=0�e=�   �   �
=�6�<����1�$Z�K����ƽ��>i���	������սLխ��.y�)����/�<��'=,�n=� �=#��=ri�=�=0=�'<�~5�ã��]��v��\s���-�Z4_�N^���	������G�ȿ�mӿd�ֿMӿȿ����n������+�^�R-�Z���F屾	�d��'�~�e���ѻ��<$�0=�H=��8=�   �   `(%<�G��h�B����0 �gE�|E;��9S���a�k�e���]�{UK�Ǻ/�|�� ϽKp���J޼ ��;���<��J=��p=�l=�f5=�3�<�6ܼ����Lg2�Hѐ�[�Ծ��+�=�T�j�A܊�oѝ�ܘ���鵿��6q��+ɫ�hۜ��i��<�ݏ�J�Ծo���&6�B�ý:U�pP�;���<�K)=i%=�&�<�   �   ������p�\�ӽ(-��TP��[��z������u���\Ӷ�!ڱ�dD��>E���@u�c�@�Z1��/���B)��������<�'.=2HJ=��3=���<ȫ�0�x����!Tb�/�T,�Ԛ��i@�2�d��q����wΖ�NT���O������V����b��L>�����y�L���t`����<Ѐ��>g���<��=:`=�^�<��
<�   �   (�u����Y�1�˩v��@���¾��������<U���gi���۾�Ỿ<_���0h��"�u|ɽ��@�`Zػ���<�=е(=��<�Q�;<������jF%�\���������D��4�P�N�M8c��p�St��o��ka�ppL��2�Gl�������y���������W�;�$�<=ܿ�<��C<����   �   �Y۽��4�T����𱾜����͉�)�,�y�6���9��5��*���.�G�۾�髾�w|�z>*���Ƚ�1���>�(Ŀ<D�=l�=�b�<(����P�jQ۽h�4�����q챾~���������,��6�J�9���5���*����+�(�۾�櫾�r|��:*��Ƚ\�1���>�lȿ<�=��=8X�<X����P��   �   #K%�?_���õ�t��+�g�4���N�$<c��p�6#t�Co�8oa��sL�^2��n����冱�.�y����,���� �B�;$�<�=H��<��C<��J�u���彀�1���v��<���¾b������	�6R���c��0�۾�ݻ��[��
+h���"��uɽ �@�0%ػ���<��=��(=��<  �;���z����   �   PYb������0�{���l@���d�xs���󎿃Ж�TV���Q�����mX��V�b�SO>�����|�v���w`����Ҁ�8Jg�(�<"�=vc=�i�<h�
<�����p��ӽY'��MP��W�����T�������tζ�fձ��?��EA���9u���@��,�2(��|7)� V�����<�*.=�HJ=�3=���<���ȑx�����   �   �Ӑ���Ծ	 ��=�x�j�ފ�Xӝ�ۚ���뵿��s���ʫ��ܜ� �@i�Ѧ<�>��R�Ծޜ��6���ý�W�J�;���<(N)=Xm%=T3�<�K%<�0����B����u��>?��>;��2S�Q�a��ze�^�]��NK���/��v�Z�ν�h��(3޼`�;���<��J=��p=�l=�d5=�*�<�Eܼ]���Dk2��   �   @y���v��"-��6_��_��x��a���#�ȿjoӿ5�ֿ	ӿ�	ȿ���o��������^�7S-����w汾��d��(���e�Њѻ���<�0=8	H=��8=d
=<H�<H����Z� ����ƽ<���]���������ܯս̭�vy�B�`9��A�<��'=��n=#"�=���=&i�=\;0=X<"�5�^���]��   �   زʾ���}�D��|��蚿�F���dοS�Lc�o������Ϳ�������dC}�/�E�U$�N�ξ���P�3D��̟���4�<R1=|_^=޶e=:P=�<%=d��<P�)<@�Ȼ�Z���D�d<9��O��Q���=�J��n��p^���{q<:D=B�V=)֊=���=��=J��=�a�=�g'= 2E��v�V��A(���   �   4&� �n_W��Ɖ�)����ƿ࿭���.� ��(�^� �9x�����<ƿ���ނ���>Y�F"��]�����E6�<�����ݼ��<�s.=�k=뛁=�=n4g=&_B=،=���<��w<@L�; ��`�X�`k9� �:��<h(�<|Y	=��D=H�=��=���=���=솾=ڊ�=y2�=p=`��%Z���v'��c���   �   8��CB)��3c����%8���пY�: �\z���	�x�)� �2�뿕�пV��}����e���+���.��-�D�|�˽�����J<Ј+=�Yr=��=[��=U��=p>t=*�T=��3=�=D��< `�<�k�<��<(��<�v="�6=�Uc=���=̉�=�Ķ=���=�P�=�$�=�@�=��=�)=�+A��8���4��%���   �   ���&m,�Cg�X���r0��wӿ39￞���	�L6���	����p��3!ԿT������i�!Q/�����H�����I�>�ҽ����7<�X*=�jt=���=CW�=Ɍ=�C�=�2i=�0L=. 1=0�=n�=�=p�
=�e=>o4=�YW=�\�=ᣖ=���=��=X��=���=��=�k�=�}�=�=��[����x>9�⁞��   �    ��tA)��2c�>��d7��пX뿱~ ��y�(�	�rw��� �/�뿯�п������~�e���+����A��۾D���˽0��h�J<:�+=�Zr=-�=���=���=�>t=��T=�3=d�=���<D`�<�k�<��<P��<�v=.�6=�Uc=���=Љ�=�Ķ=��=�P�=�$�=A�=���=+=�"A��6��ʯ4�%���   �   �#ྊ	 �t]W�zŉ�����ƿ;࿢���� ��'�F� �&v���	�3;ƿ5
�������<Y�jD"�N[������6�������ݼx�<�v.=(�k=���==�5g=*`B=��=��<��w<�O�; �� �X��h9���:��<l(�<|Y	=��D=f�=��=��=䜽=N��=v��=p3�=\=t��V��Ft'�b���   �   ��ʾ�����D�~�|��暿1D��3bοFP�N`�wl�����'�Ϳh��|����?}�Y�E�"���ξ����=?�������>�< !1=pb^=8�e= P=(>%=��<�)<��ȻY���C��;9���O���Q���=�L��n��P^�� |q<`D=|�V=\֊=S �=l��=.��=<c�=�k'= ?�؃v����%���   �   hu���q���
-��2_�]]�����?�����ȿ�kӿ��ֿnӿCȿ���
m��@�����^��O-�����~ⱾЦd��$���e��Fѻԝ�<��0=�H=��8=�
=L�< ;�����Z������ƽ���]���������߯ս̭�|y�D��8�0B�<6�'=��n=�"�=Я�=�j�=R@0= 2<H{5���y�]��   �   �ϐ�W�Ծs�k�=�%�j��ڊ��ϝ�#����絿�1o��.ǫ��ٜ��i�L�<������Ծ�����6��{ý�J�@��;8��<8S)=:q%=h9�<�U%<�,����B�N������?�w>;�f2S�=�a��ze�\�]��NK���/��v�V�ν�h���2޼��;D��<.�J=F�p=^l=j5=0;�<$.ܼΐ��=e2��   �   �Pb��p)����?g@�l�d��o������̖�IR���M������T��
�b��I>����6u����Zo`�����ɀ��g�$�<�=�h=�q�<��
<�����p��ӽ�&�LMP�mW������I�������qζ�dձ��?��GA���9u���@��,�(��7)�0O��x��<"-.=�LJ=��3=d��<x��h�x�����   �   7C%��Y��޼�����h�4�4�N��4c��	p�rt��o��ga��lL�`2�`i������q�y���+y��X�Ч�;�6�<�=8��<��C<�야��u�����1�;�v��<���¾P�� ����	�6R���c��2�۾�ݻ��[��+h���"�wuɽP�@�pػ��<�=T�(=$�<�}�;:���ﵽ�   �   WK۽^�4�/���鱾W�ᾃ������,���6�ǿ9���5�n�*����(��۾6⫾ck|��4*�ڛȽ&�1���=��ۿ<��=��=�k�<x��
�P�dP۽��4�����N챾_���������,��6�L�9���5���*����+�.�۾�櫾�r|��:*���Ƚ*�1��n>��ο< �=6�=�m�<x����P��   �   N�u�����1���v�9��{¾z�ྛ�����3O��#^����۾�ػ�[W���#h���"��kɽ�q@���׻³<z�=^�(=�%�<�q�;F��}��E%��[������p��8��4�N�N�L8c��p�Ut��o��ka�spL��2�Jl�������y�����������m�;x-�<�=���<��C<╼�   �   ����ȩp��ӽs"��GP�T���������˶���ɶ�|б�>;���<���1u���@��&�N��b')��큻���<�3.=QJ=�3=��<X����x�j���Sb��8,�ʚ��i@�,�d��q����wΖ�OT���O������V����b�M>�����y�H���t`�����π��5g��
�<Z�=8h=Du�<�<�   �   @k%<����B�8�����9�\8;��+S��a�-se���]�JGK���/�gp�q�νx_���޼�k�;���<��J=��p=�l=�k5=�;�<t1ܼÒ���f2�&ѐ�?�Ծ��$�=�P�j�A܊�pѝ�ݘ���鵿��8q��.ɫ�iۜ��
i�	�<�ޏ�H�Ծe���6���ýlS�pg�;���<4R)=4r%=�?�<�   �   x
=�W�<P�������Z�����}�ƽ���S��d������ �ս�����y��
�@���Y�<��'=d�n=�%�=�=>l�=�A0=H3<l|5� ��Զ]�|v��Is���-�U4_�M^���	������J�ȿ�mӿg�ֿOӿ"ȿ����n������,�^�R-�X���B屾�d��'�$�e��tѻ���<0�0=�H=v�8=�   �   �"P=B%=D��<0�)<�ȻpC��|7�
.9���O�D�Q��=����Q��`�����q<nN=�V=�ي= �=���=ண=rd�=Xm'= X>� �v�l��P&��M�ʾ!����D���|��皿E��Ecο�Qῷa��m��H�࿶�Ϳ�������CB}�Z�E��#���ξ����?C�������7�<H1=b^=6�e=�   �   8=�7g=rcB=�=,��<��w<���; �	�@$X� �8�@ �:(�<�:�<�a	= �D=�=	�=���=ݞ�=䈾=ʌ�=|4�= =�i�fV��&t'�b��$྽	 ��]W��ŉ�����ƿ��y����� �D(��� �`w���[<ƿG������^>Y��E"�x]徢���.6�4�����ݼ8�<�t.=D�k=ל�=�   �   ���=���=@t=V�T=L�3=X�=���<@h�<�t�<T��<���<J{=��6=Zc=���=���=`ƶ=r��= R�=�%�=B�=���=-=A��5���4��$�����DA)��2c�5��m7��4пPX��~ �z�t�	��w��� ���s�пK�������e���+�i������D�o�˽J���J<T�+=�Yr=��=�   �   Hnx=p�r=L�f=�nX=�J=
�?=��8=��7=��==,�J=&_=�z=�+�=b�=
��=���=�=���=���= ��=gJ�='�=��q=D �<�����彰Y�i������,��F^��􈿓���������ȿiԿ�׿�ԿɿU񷿽7������<`�wk.�b4��ᴾ��k�p�
�.S��@�v�(�<��&=6Z=�rr=�   �   6	s=�jj=�5[=�I=ċ8=H*=�� =:Q=�m!=��-=ndB=�_=�<�=�I�=<S�=���=��=���=vB�=���=L^�="y�=j�s=���<n���߽b�S��Щ�4�����(��UZ��������������ſI}п�9Կ{п��ſ
δ��g��1���[��+��7��D����;f����-��kW���<��(=��Y=��o=�   �   b,b=��P=��7="�=�� =8�<t3�<0U�<L�<�0�<���<a
=(_3=v�b=⬊=���=M�=V��=e�=J��=nr�=Eu�=x�w=��<�!�TJ˽*<E��_���v龼����N�5r�W��<���A绿�>ƿW�ɿz(ƿͻ�g����9������P�o!��'�W�����U�l���V�]� ��� �<�8/=�X=vg=�   �   ��C=�8#=h��<��<� �;��0�.�ꄼ����s9��T� b*<|�< �(=HAj=E��=���=���=z�=$�=e�=�|= D�<;��~{��FM.����TWӾ?P�~�<���i�8���j���X����0���e������_���h��;l����i��j=�o^�Я־����?�;�@�н�(*��rX:,[�<��7=�U=�V=�   �   b�=�ѽ<P��;�H&��J��	4���l�#���J�������,��� �a���pD�� 0;�2�<�h7=�R�=�}�=�f�=�R�=^b�=jj�=�t=7�ƅ�^��u��R���	��h�%�CN��u�񵋿4&��E���4��ce��|���S1���0t��M���%�%���O����A{�(�������Ѽ(�8<�X=Z�>=��K=��;=�   �   �s�< @˸�xļTYL��'���XϽ�������V(�����\����ٽB��*�M���� a<@c	=�i]=%�=7��=�s�=n�=�;%=��;x�5�G�oG�1ᗾ��Ծ �}�.�v�P��pn�4䂿 F��ఌ��[K����l�O�Ӕ-�n�
���Ӿ>���a�H��j콮�Y�(�(#�<�Z%=B=��9=�=�   �   ��Ǻ����0���&ѽ���L�4�;�U�o�n��~��Ӏ��y���d���F�H�!���#[���:���d�� �<N9C=$�{==b�z=b9=茏<���C���&��Ao�!H��T⾪J��|*�xC�
W�'ec�&`g���b���U�S�A��f(�~1�,l޾�릾d�i�l��>ǟ��)ټ ;(<�
=j�9=t>=�=,��<�   �   �0�1����e�/ ,��Hb�[E��!]���V��.s��K�¾�@���������Q��h�O����f+ĽD�G� a��<�j4=�<e=J�k=L�F=���<�1^��B�s�Խ��0�G���U��4/ݾ*K��n��5)��$3��D6�hH2���'� /�����j׾�|��6Nw���&���ý�*� �!�`��<��2=�G=�t0=���<��[;�   �   �ׂ�t��8��}�xF���iƾM������[�����\��4��o?�Fֿ��ћ��n���'�XCѽ��K��������<L�/=t�S=�K=��=��b<Tɢ�fт�E��n8���}��B��NeƾS�徦������'����� /��;�zҿ�RΛ��n���'�:=ѽ
{K��������<P 0=��S=n�K=4�=��b<ۢ��   �   ��Խ\�0�
J���Y���3ݾ�M�|q��8)��'3��G6�TK2���'�k1����wn׾����Rw�B�&�q�ý�*��	#�|��<4�2=�G=Zw0=`��<@T\;�j���]��,�\Bb��A���X���R���n����¾q<��m������N���O�J��[$Ľ��G��A��<2n4=$>e=��k= �F=���<`�^�BB��   �   
��go�lK��+X�M�^*�{C�DW�chc�Zcg���b���U�؜A�
i(�K3�o޾��i�����ʟ��2ټ�0(<�
=ܘ9=t>=��=ȕ�<�{ƺy��y)���ѽV��F�4���U�2�n��~�*Ѐ��y�5�d�s�F���!���S�� /� �c�$.�<�=C=��{=^��=x�z=8_9=���<��������   �   �G��㗾 �Ծ7���.�8�P��sn��傿�G��s���:񉿻L���l�!O���-���
��ӾҒ����H�n���Y��"� !�<�Z%=�B=z�9=j =`��< H�� cļ�KL����;OϽ2������"�Ň��V�� �~�ٽ����ȉM�|�����<�j	=�n]=�&�=��=t�=^m�=68%= ��;��5�E��   �   �u�KU�����l�%�jEN�]u�[����'�����������f������j2���2t�o�M��%���������xC{�o�A���|�Ѽ��8<Y=V�>=�K=�;=.�=�޽<���;H &��2���3�<�l��튽����3󔽽y���a�F
��*�� �;�D�<�o7=�U�=��=$h�=}S�=<b�=i�=Fq=pe��ʅ�a��   �   ����YӾ�Q�N�<���i�^�����������52���f������`��hi���l����i��k=�_���־E����;�5�н�)*��YX:�[�<l�7=:U=|�V=6�C=v=#=,��<L#�<�E�;@i���.��҄�8֖� ډ��D9������*<|1�<��(=�Gj=Պ�=���=��=I�=[�=�d�=�|=�<�<4F�����P.��   �   �a���x�����N��s�?��-���4軿�?ƿ6�ɿC)ƿ�ͻ�����k:�����P�mo!�(���֪U�����&�]����,�<�9/=n�X=Jg=�.b=��P=f�7=�=d� =�<�A�<Hd�<��<@@�<��<8h
=�e3=�b=N��=���=��=|��=�e�=���=^r�=�t�=X�w=L��<�+��M˽�>E��   �   �ѩ�������(��VZ�>���[��G����ſ�}п:Կ`{п�ſ<δ��g��1���[�|+�G7�� ���-;f�n��,�@fW���<��(=�Y=�o=�
s=�lj=08[=��I=ގ8=rK*=R� =U=�q!=|�-=hB=R_=>�=K�=TT�=b��=���=<��=�B�=���=�]�=xx�=Z~s=���<����߽J�S��   �   Jj�����,�G^�������,����ȿ}Կ�׿~Կ�ɿ �~7��f����`��j.��3�ᴾ��k�r�
��Q����v��+�<�&=`Z=�sr=,ox=>�r=�f=FoX=��J=��?=�8=&�7=�==J�J=_=�z=�+�=,�=̶�=k��=��=J��=~��=���=�I�=k�=��q=��<�������Y��   �   �Щ�{����(��UZ������������E�ſ�|п9Կ{zп�ſpʹ��f���0���[��+��5�� ����9f�\���(��\W���<"�(=d�Y=&�o=�s=~mj=�8[=Z�I=~�8=�K*=�� =^U=�q!=��-=:hB=j_=>�='K�=ZT�=l��=���=J��=�B�=���=<^�=�x�=�s=d��<����߽��S��   �   �_��nv�s��2�N��q���������滿�=ƿ|�ɿ�'ƿ̻�t���9�����P��m!��%����U�q���$�]�����L	�<�</=��X=Vg=�0b=b�P=��7=<=�� =��< C�<pe�<��<�@�<|��<^h
=�e3=4�b=[��=���=��=���=f�=���=�r�=�u�=��w=\��<t!�2J˽�;E��   �   ��pVӾ�O���<�q�i���������]����/���d��N ��V^��Qg��k����i� i=��\�H�־����3�;���нD!*� �Y:�e�<`�7=�U=h�V=��C=�?#=T��<�&�<�R�;�T�8�.��Є� Ֆ�@ى�XC9����h�*<�1�<Ν(=�Gj=�=���=d��=��=�=�e�=j�|=�F�<�7��az��xL.��   �   �u�UQ�����:�%��AN��u�޴���$��쩡��}���c������/��.t���M���%���������D={���|���x�Ѽ�8<�^=�>=�K=��;=0�=�<���;�&��.�d�3��l�Y튽G����򔽓y���a�&
��*�� �;�D�<
p7=�U�=��=�h�=\T�=�c�=�k�=4w=P �ą��\��   �   �F��ߗ���Ծ�	���.�a�P�Vnn��₿�D��N���!�I����l�<O�X�-�L�
�:Ӿk�����H�d� �Y��� ��1�<Za%=� B=��9=($=��< T���]ļlIL����mNϽ����·�V"�����V�� �j�ٽ������M������<�j	=�o]=}'�=��=�u�=�o�=�>%=��;v�5����   �   ����o��E��5Q��H�yz*��uC�LW�bc��\g�a�b���U�S�A�d(�/�h޾q覾��i��������ټ�](<&'
=��9=�>=B�=d��< ƺs��((���ѽօ���4�2�U���n��~�Ѐ��y�.�d�n�F���!����S���.�@�c��/�<?C=��{=伇=�z=�e9=ܕ�<p��x����   �   ?�Խ8�0��D��"S���+ݾI�@l�3)��!3��A6�WE2���'�/,� ��wf׾�x���Gw�ߝ&���ýP*� e�l��<��2=:G=�|0=���<`�\;�� ����[�7,��Ab�nA���X��gR��vn����¾k<��j������N���O�B��@$Ľ"�G��>�L�<p4=Ae=Z�k=~�F=X��<��]�&B��   �   ]̂����:8�;�}�Y?��waƾ�徾������k������)��6��Ϳ�Xʛ�� n��'�04ѽ�lK��N����<p0=2T=
�K=��=��b<�¢��ς����8�
�}�cB��*eƾ7�徕������$�����#/��;�zҿ�RΛ��n���'�=ѽpzK�0���h �<�0=� T=h�K=��=��b<๢��   �   �	�{{���U�,��<b�G>��&U��KN��j����¾�7����������J��3�O�����Ľ��G�H�t+�<�v4=�Ee=.�k=��F=��<��]�&B�;�Խ"�0��F���U��/ݾK��n��5)��$3��D6�iH2���'�/�����j׾�|��/Nw��&�b�ý*���!���<f�2=G=&|0=��<��\;�   �    wź�d��#��ѽ�����4�@�U�P�n��~�_̀��x���d���F���!���aJ��L� ,c�dC�<�FC=X�{=̾�=P�z=�f9=��<���������o��G���S⾚J��|*�xC�
W�&ec�(`g���b���U�U�A��f(�}1�-l޾�릾W�i�R���Ɵ��'ټ�B(<�"
=М9=�>=��=���<�   �   ��< T��Nļ?L����FϽX��������ف�Q�����ٽ����xM�����<u	=�w]=�*�=k��=w�=�p�=L?%=`��; �5�T�
G�ᗾ��Ծ�s�.�q�P��pn�5䂿"F��Ⰼ��\K����l�O�Ԕ-�n�
���Ӿ:���M�H��j���Y�@��'�<<^%=PB=��9=�%=�   �   ��=��<�%�;��%�t⼢�3�\�l��劽	���aꔽ�p��
va�@�������;L[�<|y7=�Y�=���=(k�=4V�=�d�=Ql�=�w=0%�Ņ��]��u��R��q	��`�%�CN��u�񵋿6&��G���8��ee��~���T1���0t��M���%�&���L����A{��L���|�Ѽ8�8<�[=V�>=��K=b�;=�   �   �C=LB#=��<�1�<���; ��@k.����� ���@����9�@��`�*<�F�<$�(=�Oj=l��=���=���=��=��=�f�=��|=,H�<�7���z��M.����@WӾ7P�x�<���i�8���l���Z����0���e������_���h��=l����i��j=�p^�ϯ־����0�;���н�'*� �X:_�<j�7=�
U=��V=�   �   01b=��P=$�7=\=�� =��<�N�<�r�< �<P�<���<�o
=�l3=��b=f��=j��=B�=���=�g�=X��=t�=tv�=F�w=���<���I˽�;E��_���v龸����N�4r�Y��;���A绿�>ƿZ�ɿ|(ƿͻ�h����9������P�o!��'�U�����U�H�����]�����X�<�:/=��X=g=�   �   �s=�mj=�9[=��I=�8=N*=R� =bX=u!=B�-=�kB=*_=�?�=�L�=�U�=ߺ�=���=p��=�C�=���=_�=�y�=B�s=��<���w߽L�S��Щ�/�����(��UZ��������������ſI}п�9Կ{п��ſδ��g��1���[��+��7��D����;f�ޜ�h-�HjW���<b�(=4�Y=t�o=�   �   v�=�D=��=~=r=H�&=��3=�E=�HZ=8_s=E&�=�g�=Y�=FR�=�Y�=��=��=x�=��=4&�=���=*Q�=x��=�VC=p1�;`[�.����d�]}��a������E�<�k���������t��@`���x������膿��l�!G�� ��(��	մ��ny�q|��˵�pE$�0 ׻� x<�u�<D=\=�   �   bc=�[=�[=��=J�=j%=��"=B�1=~qE=p�]=V�z=Wٍ=��=</�=�5�=���=�&�=X=�=�Z�=�f�=0�=H��=fޡ=�OF=0��;4~Q�9 �(�_�`ꩾ�T�`��e\B��g�`���i����������M����q�� ���P9h�9_C�Ak��&�$밾�xs���3���:��ᙻX��<,��<m=(�=�   �   ��=2�=d�<$X�<�[�<�<���<���<��=�x=@(8=`0[=Q��=�]�=�v�=���=�*�=���=���=��=���=�+�=⌢=ءN=h(#<B�5��o�d�P�U�����߾a8��7�*}[�8{��Y㑿0���6ԑ�Pቿ{��[���8�>i����E����,b���y���L�� a7:Tt�<�/=L�=�J=�   �   �a=���<�ð<0��<�1,<p��;���;@�l; �;"<E�<8�<��=26O=c�=�=@��=��=���=*��=�C�=N��=a�=��Z=l��<��r�ʽVV9�H~����ʾ����'��tH�ԕe���|����A��zn���|��)e��2H�c�'�]���̾ᓾ�/G�<{�&�z�(���h=<�1�<��=��=Z;=�   �   0%�<`_�<�'�;@�Q���^�l��\��('�^I����Zɼ@�`� ��9���<>E=@�R=��=;�=���=���=�)�=@�=M��=P�g=��<X����s������v�Bͯ�Ŀ����?0�K;J��^�ޭk�tp��Bk�n�]��XI�pb/��V��4R��C�z���$�ڿ�$%-��^�����<�1=�?%=ܨ%=^-=�   �   ��<P�;X�G�(p��ނA�~��K����ʯ�K�����������s����AO����p�ϻX�<��=�o=�Y�=X�=ټ�=�=�Ş=��r=T� =@T�v�k��/���I�^���c�þO�������I+���<�xH�0�K��qG���;�9�)�z\�Ur��\������nH�u���Z�����x�.<���<��*=
i6=j�'=��=�   �   `�;0Xn�� �OC��,i��
[�Ǝ�-��x�&�Lz'��Q�������P���Z�m���ܼ��0;Ds�<r�P=�=��=xӢ=�Q�=.�y=	= ��;R��rd�������f��Ɯ�C�Ǿ�T��+�4���"���%�a "�FD��+	����an¾v���$]�����ʫ��Y��M�:��<�.=ZcH=F�B=��!=���<�   �   (��( $�*a����ɩ�օ=���]��nv���������~�B7j��K�RG&�����n���"*��л6�<��<=<�|=�W�=6�=Șy=��4=��<��{�x�n������,���n�����Iͺ�A2ؾC5�X���l� �&����l�4�Ҿ^���瑾L6^�m���8�� 9��:��(��<x�/=ƦY=F�`=ԥG=rx=���<�   �   ���y\��];�Ú+�/`��S��d�������q���߄��1��N"�����(H����J�e�� �����C�(��8�<�3=xQj=N�~=�eq=�-C=�F�<`];h���V���3��+��`��P��¡�����e���Ӏ��8-�����Ό��QE����J��������*�C������<p3=�Sj=.�~=,eq=�+C=(?�<� ;�   �   T�n�W��C�,�>�n�Į���к�c6ؾ�9������ �����q���Ҿ��nꑾ�:^�����=���'9��g��d��<�/=p�Y=,�`=�G=*{=��<8����#�[��&�"��m�=�t�]�hv�V�������~�1j�n�K�rB&�����Fg��*��@л�B�<T ==F�|=�X�=^�=��y=��4=H��<`�{��   �   �i�������f��ɜ�ŴǾ�X�6.������"���%��""�fF��-	�ڈ�q¾Jx��(]����hΫ�X_����:���<.=�bH=��B=��!=l��<�/�; ;n�j� �5=���a��fR��������&��t'�tL�������B�����m�<nܼ�p1;���<��P=���=9��=Ԣ=�Q�=��y=�=0Z�;H���   �   �5����I�����s�þ������,L+�M�<��H���K��sG���;��)�^��t��r��e��ZqH������\��tĪ�P�.<г�<��*=,i6=��'=�=t&�<�;pG�t]��rwA�hw��ë���¯��������������z3O�\��pnϻ��<�=�o=�[�=��=���=��=�Ş=��r=�� =����k��   �   ����v��ϯ���龹��A0�q=J�#�^�"�k��p��Dk�U�]�rZI��c/��W�� 龕S��E�z�B�$�,ܿ�(-��o��Џ�<&1=�?%=��%=�.=�*�<Lg�<PS�; �Q��^���Х����<���@Aɼ0�`� �9,ć<�M=D�R=a��=s�=X��=���=*�=G�=���=�g=��<l����w���   �   Y9�����ʾ+����'��vH���e���|����-��Vo��/|��*e��3H�D�'��]���̾�ᓾ�0G��|���z������9<�0�<��=n�=p<=�c=T��<T˰<���<�I,<���;0��; m;�1�;�7"<�V�<L��<b�="=O=b"�=��=D��=���=���=���=�C�=��=��=�Z=l��<^!���ʽ�   �   ��P�ؑ����߾~9�O�7��~[��{�9�䑿ژ���ԑ��ቿ�{�ĺ[��8��i�;�㾒���-b�,�������� \7:pt�<�/=��=`K=2�=
�=\�<�^�<�c�<@
�<���<ȧ�<��=�~=�-8=�5[=ծ�=�_�=�x�=*��=2,�=x��=���=2�=���=7+�=��=^�N=�#<p�5��s��   �   ��_��멾IV�*��C]B�ͦg��`�� j��-���V��������q��F���z9h�J_C�>k��&��갾�xs�j�����9�pۙ����<<��<�m=�=Ld=�\=]=��=x�=�'=P�"="�1=|tE=b�]="�z=�ڍ=��=70�=d6�=T��=z'�=�=�=�Z�=�f�=�
�=ɔ�=�ݡ=�MF= �;x�Q�v: ��   �   ��d�~��*	�\���E���k�ݺ��<����t��A`��wx��l���膿:�l��G�}� �0(��ZԴ�xmy��{�ʵ�C$���ֻ�x<�w�<<==6�=BE=X�= ==��&=
�3=�E=IZ=b_s=E&�=�g�==�=R�=�Y�=d�=��=,�=:�=�%�=���=�P�=���=�TC=��;t[�(���   �   ��_��ꩾU�h��Y\B���g��_��{i���������澙�q������d8h�Y^C�uj�\%��鰾ws�D�����6��ə����<���<@o=\�=�e=<^=F^=��=h�=�(=��"=��1=�tE=��]=^�z=�ڍ=�=E0�=r6�=d��=�'�=�=�=[�=�f�=*�=��=ޡ=OF=��;�Q�o9 ��   �   �P����G�߾8���7��|[�e{����⑿�����ӑ������{���[�J�8�h�ѝ㾮���<*b���R���<����l8:�{�< 3=·=,N=��=��=��<�b�<�g�<l�<h �<Щ�<h�=B=t.8=*6[=�=�_�=�x�=D��=N,�=���=���=~�=��=�+�=��=(�N=p)#<��5��o��   �   ZU9��}����ʾ)��3�'��sH���e�&�|�=���U���m���|��'e�1H�̷'��[���̾!ߓ��,G��v󽤐z����� R<�:�<(�=��=R@=�g=0��<�Ѱ<���<�S,<���;��;@$m;�:�;(;"<0X�<,��<��=h=O=~"�=��=f��=���= ��=D��=vD�=��=�=�Z=���<���ʽ�   �   0�Вv��˯������g>0��9J��^�ͫk�B�o��@k�.�]��VI�q`/��T��龡O���z�|�$��Կ��-��(��D��<N7=E%=��%=�3=D3�<|o�< q�;�YQ��^�����J�F;�(���?ɼP�`� 2�9�ć<�M=��R=���=��=���=\ �=�*�=V�=V��=��g=��<����Zq���   �   �+����I�����H�þ����R��H+���<�3H�ʦK�4oG�/�;���)�bZ��n��+��"	���jH��z���T������p/<���<��*=,o6=�'=��=�/�<`6�;�_G�V��:tA�v�������������k���/���E���3O���� lϻ<�<l�=o==\�=\�=���=:��=dǞ=��r=�� = 1�k��   �   6`����f�f��Ĝ���ǾXQ�*�����"�"�%��"��A��)	�u�쾻j¾ s��~]�����ë�O��e�:���<L.=�iH=��B=R�!=���<�V�; )n�\� �Y;��&`��Q�\��|����&��t'�EL�������$���P�m��mܼ@u1;���<~�P=2��=��=Aբ=SS�=Фy=8=p��;����   �   ��n� ��o�,�y�n�ި��ʺ��.ؾ.1����#� �����h���Ҿ���p䑾�0^�����0��n9�`鿻Ͽ<��/=z�Y=��`=�G=��=Ɂ<�s���#� Y��i�b���=��]��gv�2��������~��0j�Z�K�dB&�l���%g���*��=л�C�<D==ػ|=�Y�=��=ʜy=$�4=��<�{��   �   ̸�jQ��@-���+��`��M��n���Q���m����|��)���������A���J�f��t}��2�C��n�l��<R3=�Zj=��~=�kq= 3C=�P�<@�;4���T��>2�[�+��`�XP����������H�������+-�����Ȍ��NE����J�{��䅿�ܺC�h��p�<�3=�Uj=\�~=�iq=^2C=�Q�<��;�   �   �e���#��T���
佾��P{=���]��av�񆂾*	�� �~�H*j��K��<&�X����^��H	*�`�ϻ�V�<�==~�|=�[�=���=n�y=t�4=D�<ȕ{���n���<�,�>�n�H���ͺ�2ؾ%5�E���f� �����l�/�Ҿ]���瑾F6^�d���8���9� 5�����<R�/=��Y=Z�`=��G=��=H́<�   �   @j�;�n��� ��6��FZ���I������c�&�o'��F�X��^��Ԗ��޵m�@Qܼ@52;,��<l�P=O��=k��=ע=�T�=�y=@= ��;
���b��(��R�f��Ɯ��ǾxT��+�+���"���%�` "�FD��+	����^n¾v���$]����fʫ�2Y�@m�:��<�.=�fH=<�B=��!=���<�   �   3�< O�;PLG�\H��BkA��p�����(���񆸽䠵������틽#O�d���ϻ�-�<
�=
!o=v_�=��=}��=���=^Ȟ=��r=�� =`<�ʒk��.����I�$���2�þ)�������I+���<�vH�0�K��qG���;�:�)�y\�Tr��Z������nH�L����Y�������.<���<J�*=m6=�'=,�=�   �   �4�<ls�<���;�
Q��~^�4޹�D��<�6/�p���%ɼ��`� 9�9ۇ<�W=@�R=@��=��=1��=h�=j,�=��=*��=f�g=��<�����r��A�~�v�ͯ�������?0�I;J��^�߭k�xp��Bk�r�]��XI�rb/��V��4R��=�z���$��ٿ��$-� X��8��<�3=�B%=8�%=D3=�   �   �g=8��<�հ<8��<Xe,<p��;0C�;@�m;�}�;�^"<xj�<,��<H�=fEO=&�=��=%��= ��=��=���=�E�=���=��=��Z=P��<����ʽV9�&~����ʾ����'��tH�ԕe���|����B��{n���|��)e��2H�c�'�]���̾ᓾ�/G�{󽼗z�௞�@A<�4�<�=�=�?=�   �   ��=��=�<\f�<�l�<�<��<X��<��=ք=848=�;[=���=�b�=M{�=b��=*.�=<��= ��=��=��=�,�=���=P�N=X-#<,�5�|o�4�P�B�����߾\8��7�(}[�8{��Y㑿1���7ԑ�Qቿ {��[���8�>i����D����,b���\���p����7:@v�<�0=D�=NM=�   �   .e=^=z^=$�=V�=*=��"=��1=NwE=Z�]=0�z="܍=d�=�1�=�7�=���=�(�=�>�=�[�=�g�=��=ӕ�=�ޡ=�PF= ��;�}Q��8 ��_�Xꩾ�T�^��c\B��g�`���i����������O����q��!���Q9h�:_C�Bk��&�$밾�xs���%��Z:�Pߙ�4��<p��<n=|�=�   �   `V:�`����H:��;�R<8��<���<T�'="IR=\�|=p��=�=���=&H�=v�=�v�=���=�1>��>b=>:��=��=���=�i�=��= ʲ��Rz�q��Z�̸���,վ�����"�F6;�*�N�N5[�D�_�~:[���N���;�I=#�l;�D�پ������o�g#$�S�ѽVOv�,� ��7a�����{���u���,
��   �   �p
� �� :0��;(�:<��<�5�<2=V D=<�m=&�=��=,��= m�=���= �=B;�=B>)R>�>�8�=�=��=[��=p=�M����p������U�Er����о|b���U�7���J��7W�Tq[�/5W���J���7�] �^���վy���+j����,�ʽ0�j���8�?���3��: u�9 ����   �    ��@��� Ϲ�.;���;�pS<��<(+�<^�=(~?=Zgh=v�= �='��=��=��=h%�=���=|;�=���=x�=� �=���=s�=��'= �8��U��ｾ�G�>���F�ľ����6���-�i�?�'�K�O��K�)�?���-�u���O��s�Ǿ�l��JJY��M�7���8�H������]���~";`h�; l�;�B;�   �   �w; a� 32��@� ƺ ��:q�;p,><�$�<Ԭ�<�!=N�A=�
q=t�=R��=�~�=<B�=��=�A�=�y�=<�=v;�=�=�=R
�=ʺ4=P��;@�,��ѽ42��k����i���	��+�$�.�^�9��=��K9��t.�	��ٵ�V���x���ۆ�d�>����4۔�@���,;�`_;�D,<��E<��%<���;�   �   ���;�y�����@ZB�0(s���0 ����]�X%�@����;t��<�J =R:=�2u=�!�=���=���=�;�=�g�=Ȋ�=,�=fǺ=(��=B�B=\<��UK��L)�~{b����f�ž���nw
��4���"���%��("��i�:m	��W���þ�����c��}��:ƽ,�U��W����;X�v<�<`�<��<�P5<�   �   0��;0����.���^Ӽ.]�"q*��t>�Z�F���A��-��	�J��������:<��<��B=���=��=u��=�6�=�!�=:�=^�=�o�=FmN=��<����1r������s:������^���ɾ��辂� ���rG����1���3�n�ľڠ��x�+N4��;�,���G케7�J�<���<� =���<`��<�pt<�   �   �V.;H�U�Ƚ�԰<���}�����(_���½V3Ƚ�P½Y���v ����\����x���l<��=<ic=�S�=���=怳=:�= M�=B
�=�#U=	�<�J���B5�)���?���L�Pv������x��޵Ͼ�Vܾuྶ\ھ��˾������_`y�\p<����W��`.� 4����<f�=��)=B�,=|G=���<��<�   �    �Q���ͼ�QH�*ז��ɽj�������3�ӭ%�x#%��>��{�<轮����e�� Լ &+;���<ޑF=���=E��= �=^$�=�Ň=4T=bo =p��;�ݼNÃ�ֳٽ0)���J��&x�8"��X���J"���|���c��jG��fH��`d�13��z��+��V�#���ʻ  �<.�=�SL=�|]=FU=�_6=�m=���<�   �   ��V��>-��͘��'߽*�`�4��JR�{�h�p~u���w�/+n�^Z�L�<�(s�z��n˕�j*� r��d��<j�0=z�i=N��=8ԅ=�{v=�J=j=��H<0�V��7-�8ɘ��!߽K&���4��ER��h��xu���w��%n�(Z���<�o���佶ŕ�$!� 7����<�0= �i=���=Յ=�|v=�J=&=��H<�   �   �)ݼwǃ�n�ٽ�,��J��+x�%��s����%������f��PJ���J���"d� #3��}��0��*$���ʻP��<f�=�PL=�z]=�U=B_6="n=을<��Q� �ͼ&JH�IҖ��ɽ'������\/��%��%�$:�:w�4轘����e���Ӽ�+;���<�F=��=ƨ�=.�= %�=�Ň=\3T=<m =���;�   �   �I5��-��C���L��x��ޟ���{��=�Ͼ[Zܾ��`ھ��˾����.Ś�Ndy��s<���H���4��Z�� ݜ<`�=�)=n�,=NF=��<���< x.;��U�ܲ�b�<�>�}���X��Ŀ½�+ȽI½����.����\���������l<��=�nc=V�=j��=$��=
�=\M�=
�=*"U=4�<�p���   �   v���Tw:�أ��a��vɾ���8� ����.I�K��4��66徹�ľ ܠ�$�x��P4��?��.���P케�7�$D�<���<(� =���<���<�pt<�ȡ;����0'���SӼV�rh*��j>�2�F���A�r-��	�3��@�����:<h��<��B=���=�=;��=08�=�"�=�:�=&^�=�o�=DkN=$��<D����   �   GO���+��~b����޴žϖ��x
�E6�(�"�6�%�K*"�<k�pn	��Y�{�þl�����c�{�=ƽ��U��]���Y;��v<hߧ<T�<��<hO5<���;�M���x��(KB��s�l��D���{]��� E�0W�;��<�R =�:=<9u=z$�=���=`��=,=�=�h�=l��=T,�=FǺ=���=�B=��[<8���   �   B#ѽ�2�m��������(	�-���.�ȉ9�7!=�M9��u.����������y��V܆�|�>�N��yܔ�@���3;�@�^; ?,<x�E<��%<0��; x; �`�`2���?� �ź�#�:�;�C><�1�<ܹ�<&(=��A=�q=�=���=���=�C�=B��=xB�=�z�=��=�;�=J=�=�	�=B�4=�a�;��,��   �   [����G�� ����ľg���5��,�-�{�?�4�K���O�ΈK���?�O�-����pP����ǾOm���JY�2N�������H�\����c���r";Pb�;�g�; <; ��@��� �ι H; �;�{S<l �<�2�<r�=X�?=�kh=x�=�!�=Ε�=n�=&��=`&�=P��=�;�=2��=��=~ �=<��=Kr�=2�'= �8��U��   �   4��;�U�@s����оc���7�J�J��8W��q[��5W��J���7� �l���վb��T+j�V��˩ʽ��j���h�?���3��: u�9@����m
���뺀4:p��;��:<�<D9�<*=z"D=f�m=-�=��=��=�m�=���=��=�;�=-B>9R>�>�8�=��=S��=���=0�= f���p��   �   �q��Z�_���5-վ����"��6;�X�N�h5[�D�_�h:[�r�N�D�;�=#� ;���پg�����o��"$� �ѽ6Mv�|� �h2a�	��@b���_�� #
�@L:�����I: �;�R<P��<x��<��'=jIR=��|=v��=�=���=H�=V�=hv�=���=�1>��>9=>���=�=���=�h�=��=�ܲ��Uz��   �   .����U�`r����оsb����"�7�V�J��7W��p[��4W��J���7�� �����վu���)j�*���ʽx�j������?��`3���: ��9�v���L
���� �:��;h�:<��<`;�<
=$#D=��m=e�=��=.��=�m�=���=��=�;�=4B>HR>�>�8�=��=���=��=� =�T����p��   �   q��H�G�������ľ���������-���?�G�K�ȚO�ކK��?���-�q���M����Ǿ�k���GY��K�$���$�H�d��� @��`�";���;���;`|; ���3�� �̹�{;��;��S<�$�<6�<ğ=`�?=Llh=Wx�=&"�=���=��=<��=~&�=r��=,<�=l��=��=�=���=_s�=$�'= l�8��U��   �   �ѽ2��j����!��	��*��.��9��=�]J9�ks.����������v���ن���>� ���ה����;��^_;�V,<8�E<p�%<0�;��;��_���1���?��!ź���:���;8M><L5�<���<8)=Z�A=Jq=A�=���=ր�=�C�=t��=�B�=�z�=	�=.<�=J>�=�=n�4=p��;��,��   �   �H���'�^yb�������ž��7v
�B3���"���%�'"�4h��k	��T�4�þږ��ñc��z��5ƽ�U�J�� �;��v<��<��< �<(j5<`-�;���� J���5B�s�X���
���p]����*�a�;��<xS =:=�9u=�$�=���=���=v=�=Hi�=���=*-�=zȺ=S��=�B=\<����   �   �n�����fq:�"����\��4ɾ����� �s���E���3.��00�a�ľdנ�s�x�DJ4�m5��&���6케75��V�<��<� =ؠ�<��<��t<��;�]�����LHӼ�P�d*�"g>�@�F�V~A��-��	�1��@�����:<D��<�B=���=R�=���=�8�=~#�=v;�=�_�=~q�=�pN=���<P����   �   �;5�{$��=�C�L�:t�������u����Ͼ�Sܾ��#Yھe�˾����ӿ��[y��k<��������#����<�=ě)=��,=N=X��<p��< �.;H�U� �񼎣<��}��웽�V��T�½|*Ƚ/H½��������\�L�����@�l<�=Voc=kV�=ݮ�=̂�=��=�N�=&�=�'U= �<����   �   $ݼ�����ٽ�%���J��!x����W�����1y��~`��&D��UE���d�A3��v��$��\�#��Gʻ��<f�=&ZL=&�]=�%U=�f6=~u=8��<`GQ��ͼDH��ϖ�(ɽ�������.���%�@%��9�w��3�Z��(�e���Ӽ��+;���<��F=�=j��= �=S&�=�Ǉ=�8T=�t = ݤ;�   �   ��V��.-��Ø�*߽j"���4��@R���h��ru��zw��n�V
Z�#�<�j�������.����D̸<��0=�j=���=-؅=.�v=�J=:=��H< �V��1-�|Ƙ�W߽8%��4��DR�u�h�Rxu���w�f%n��Z�|�<��n�Y�佐ŕ�� �04����<��0=�i=l��=Oօ=T�v=�J=(=p�H<�   �    ;Q�0�ͼ�?H�0̖��ɽ:���p���*��%�v%��4�>r��*����\�e�H�Ӽ�^,;о�<&�F=4�=�="�=�'�=�ȇ=^:T=bu =@פ;�ݼ����|�ٽ"(���J��%x��!�����"��i|���c��ZG��[H��Od�"3��z��+���#���ʻ4�<"�=UL=�~]=`"U=Pd6=�s= ��<�   �    �.;ȘU��񼖞<��}��盽Q��÷½@#Ƚz@½&������4|\��������l<@�=wc=�Y�=z��=턳=��=P�=�=�(U=H�<0$��\>5��&���>�ܡL��u��Ü��x����Ͼ�Vܾ`ྦྷ\ھ��˾������S`y�Mp<����4�� .�@0��`�<��=B�)=��,=(K=��<��<�   �   ���; Z�����tAӼ�K�>]*��^>�8�F�.sA���,�N	����0/���;<���<��B=n��=y�=/��=�:�=B%�=�<�=�`�=@r�=�qN=`��<ī��ap����6s:�i���K^��Wɾ���s� ���lG����1���3�j�ľڠ��x�"N4��;��+��G케�6��K�<p��<0� =���<��<0�t<�   �   $�; ���`C��x-B�8�r�����H����S]�����
����; �<P\ =^$:=Au=�'�=� �=��=�?�=k�=j��=V.�=hɺ=���=��B=\<���I���(��zb�ˡ��4�žۓ�`w
��4�}�"���%��("��i�9m	��W���þ�����c��}��:ƽ��U�W�� �;8�v<8�<��<��<`b5<�   �   `�; �_���1�@�?� �ĺ���:�ҿ;(a><�@�<��<�/=��A=�q=?�=��=E��= F�=J �=FD�=>|�=,
�="=�=?�=��=L�4=���;$�,��ѽ�2�\k�����I���	��+�!�.�^�9��=��K9��t.���ڵ�V���x���ۆ�^�>����۔�����*;��_;I,<��E<��%<p	�;�   �    ���M�� �̹��;  �;��S<X)�<<�<B�=@�?=bph=oz�=-$�=藴=X
�=��=�'�=���=D=�=b��=��=��=���=�s�=@�'= (�8h�U�y��x�G�!���0�ľ����0���-�i�?�%�K�ÛO��K�+�?���-�v���O��q�Ǿ�l��FJY��M�&�����H�H��� Z����";`p�;�w�;`b;�   �   @\
���뺀�:Й�;0�:<��<@=�<P=�$D=��m=]�=��=2��=�n�=���=|�=�<�=�B>�R>F>�9�=��=\��=���=2=0H��R�p�����U�8r����оxb���T�7���J��7W�Uq[�05W���J���7�_ �`���վx���+j����'�ʽ�j����0�?���3� ,: ��9�����   �   !��� 燽��r��fD��������Q�:D��<�P=�Y_=��=�|�=��=�Y�=�m�=���=J�>̟>

>̩>t�>���=���=4�=>�=fG=8��0n��H��<����Vh����Ѿ��<��Ym��q��p�J��6���$�Ӿ�������<�Q��"��Xս����	V���.�H�(���:�(�X��w�i燽�   �   E���,���\m��A�)�d�� Tv:�C�<W=�V=R��=PL�=b׿=�r�=(��=.��=�>�>��>��>�>�-�=J��=�|�=nI�=��=����8f��b�	e8�=U��T����;]���t����Ϟ������ϾN/��SI�� ]L�����ν^���
�J�'$�D��TM0�fN�x�m�-����   �   *�v��Ks���]�>]8�z���y�����H�c<���<�~9=u=4j�=�+�=L��=\�=B|�=2�=�`>��>�E>�\ >V��=���=J�=���=��
=p���\�O��}ؽ!�,� s��������©�>���P���O�q�����|��O¾�����{�D�<�@��ո�R$w�T]*����b� �$v��0�xP���i��   �   Q�x�T�:lH���-�(w��x��  ��]�;��<�=)?=(�u=�3�=
��=L��=4o�="��=@��=���=��=�1�=T<�=��=֥�=׋�=��= �9��.��������U�Z�z���/r��zx̾�j���V����k�FH⾀˾�`���Ꮎ��^���$�H6潒�����=������� ����
ȼ�����"��:?��   �   ��$���1���2�t;'�z_�D�(2���P� .;Al<��<�$=B�[=|ۈ=0��=�(�=&D�=���=a�=�f�=��=h��=�"�=Ī=_��=�w=0��;���e��χ�.j=�,3x�Ҕ���C�ž�|Ҿm־HѾ��þ<׮�4)��Xr���9�*#�j��Z�\z��V��IĻ������%�pj��,�ּl���   �   �\�&b�L\#��+��*��� �l������s<� 88�X<�|�<�-=��j=P��=q:�=ǿ=�k�= $�=H�=z��=-�=�[�=ey=�n=�<��ü]ŀ��Kڽ�n�"O���~�J�������N��_,���Q��*7�����J�q��@�Q�߽ƽ�)s��񼠘����;�B5<�h0<���;���@>�@S���   �   |�87���� � �?��W�&�g�*|n��cj�� Z��R<��F�d���ǻ�#:<$��<��>=Ĝ~= �=���=$0�=��=\ϸ=���=���=`&g=Y=�G<\���NH�ո��jL���&�5=L��m�k���_��*���a��h�{���\���6������ɽ��{� ���ŏ���_<�[�<PY�<k�<��<8�Y<��*;@{��   �   ��\���輺�0��Ij�����r:���H��r���ϓ����N��T冽�/C���ۼp)����< =��Y=�A�=T��=� =�8�=m�=��=�J=�= �B<�">�v��A����ZĽ�� �Z.�<�5�\H�8OR�MS���I�<|7�q�z!��3���i���׼ θL�<��=�3=8�>=�85=:�=8�<�x< I�:�   �   �N-�t����8U�������������U��H�������	�����ƽ^H����7�<����T�;��<�5=Z�d=n#~=.�=ts=�tR=R#=|��<�<(K-�|����4U�m���/����������������ښ	�g��x�ƽ�B����7�P䓼���;��<�5=��d=6'~=�/�=�s=�wR=z#=X��<��<�   �   �*>�J��:����^Ľ4� ��1���5�p#H��SR��	S���I�:�7��t��'���8���i��׼ tڸ��<�=�3=r�>=^55=�=���<�x<��:��\�t����0� Ej�a���26���C��������������G��5߆�J$C���ۼ 㞻��<Z&=�Y=�C�=G��=>Ġ=#:�=<n�=��=\�J=��=��B<�   �   ����`H�w���?Q���&��@L��m�����ua���	���c����{�h�\�7����h�ɽh�{������� �_<xS�<�Q�<�c�<��<��Y<@h*;p��,����7��R� �4�?�6�W�̱g�Jtn��Zj���Y�vH<�<<�H과 �ƻ E:<���<V�>=:�~=e�=���=�1�=4�=�и=���=���=�&g=�X=`�G<�   �   ��üXȀ��Oڽlq�dO���~�p���#��%Q���.���S��C9��l����q���@�RS�t�ƽ�/s����Щ�@��;�35<(Z0<�d�;���0!>��X��|`�6c�$\#�
+��*�v� ����Lr������R<� �X8x$X<ċ�<� .=�j=���=�<�=�ȿ=Nm�=r%�=X�=P��=�-�=�[�=�dy=�m=pz<�   �   ����h�����l=�h6x�������z�ž(ҾIo־5JѾp�þ�خ��*���r���9��$��l��,	Z���鼈�V��cĻ�·�H&�<q����ּL����$�v�1�&�2��:'��]�l�*���<���;Yl<D��<"�$=��[=ވ=���=�*�=�E�=
�=Bb�=�g�=\�=��=D#�=Ī=��=�u= �;�   �   @�.��������� [����s��Sz̾�l���7����m��I��˾�a���⎾h�^���$�8����. >�������L���ȼ�����"��=?�*Q��T�mH���-�<v�,u��p�px�;D	�<&=f-?=r�u=�5�=���=��=�p�=Z��=D��=t��=N�=�1�=�<�=��=���=I��=��= ��9�   �   ��O�=�ؽޏ,�.s��������5�Ά������P��q�"����}ᾂP¾r����{���<����ָ��%w��^*���� ��w��0�jP���i���v�$Ms�X�]�\]8����hw��`k� �c<���<N�9=�u=�k�=�,�=~��=l�=(}�=�2�=�`>��>�E>�\ >\��=r��=��=J��=��
=�����   �   j<f��d�[f8�V��/�����;�]�N�ޣ�F����(�	��2Ͼb/��TI���\L�����νL����J�L'$�����M0�0N�F�m�������� -��]m�zA��(���� �v:�E�<jX=,V=��= M�=ؿ=8s�=���=���=�>�>ʻ>��>�>�-�=���=|�=�H�=Җ= ����   �   �n�UJ��<�:���h���Ѿt��\��km��q��p�-������ӾF���Q��|�Q�="��Wս���0V���.�n�(��:���X���w�3燽⊌��懽@�r�<fD��x���@`�: ��<Q=�Y_=�=�|�=���=xY�=�m�=���=6�>��>�

>��>N�>>��=D��=��=�
�=�E=����   �   �9f��b�"e8�=U��B����;�\ﾢ�(�����e��z����Ͼj.���H���[L�v���ν���� �J��$$��� K0�:N�0�m�������+��6Zm��A�V&���� �v:�H�<�Y=V=[��=>M�=4ؿ=^s�=���=���=�>�>Ի>��>�>�-�=<��=v|�=HI�=n�=в���   �   ��O��|ؽ��,�D�r�8������ި�,������?O�Np�����?{�bN¾���u�{�B�<���Ӹ�zw�Y*�§��� ��r��0���O���i���v�^Gs���]�VX8�v���o�� 8�P�c<���<�9=u=l�=9-�=���=��=P}�=�2�=a>�>�E>�\ >���=���=��=c��=��
=�����   �   ~�.�����x����Z��q��w̾+i�	�g����i�CF⾓˾�^���ߎ��^�I�$�2������=��t����t���� ȼ�����"�@5?��	Q��T��eH���-�p��j�����;�<b=&/?=��u=6�=G��=7��=�p�=���=v��=���=��=d2�="=�=��=���=ь�=��= g�9�   �   J���b����h=��0x�L����F�ž�zҾ�j־�EѾ/�þծ�''���r���9�l �`e��(�Y��l鼈�V��Ļ�z����%�t^�� �ּb��"�$���1�(�2��2'�`V���弐���+�`�;�cl<X��<��$=�[=�ވ=Ю�=�*�=F�=B�=�b�=.h�=��=���=,$�=`Ū=٠�={=`�;�   �   h�ü����dGڽ<l�$O�H�~�N������_L���)��O���4��4����q�*�@��M�!�ƽ" s�D��{�`�;@[5<��0<��; 7���=�dC��,K��X�dR#�+���)��� �����h�xﭼXG<� ha8�*X<4��<�.=��j=1��=�<�=:ɿ=�m�=�%�=��=
��=�.�=^]�=�hy=`s=Ș<�   �   ,��� H�����F���&��9L�Ƥm�'����\�����_��}�{���\�t�6����(�ɽr�{����������_<4i�<,f�<�w�<,'�<�Y<�+;�X��ࣼ�"��~� �$�?�:�W��g��nn�Vj���Y��E<��9�糼��ƻ�H:<\��<�>=��~=��=.��='2�=��=@Ѹ=���=��=+g=|^=H�G<�   �   �>����5����TĽF� ��*�*�5��H��JR�� S���I��w7��l�{��^,��2
i�\�׼ `��l"�<֝=��3=��>=J?5=�=��<��x<�j�:X�\�|�輒�0��<j������2���@��y���Ӌ��=���F��wކ�(#C���ۼ ޞ���<�&=X�Y=!D�=���=�Ġ=�:�=9o�=F�=^�J=(�=@�B<�   �   �*-�h���\*U������|���������;�������	� ���ƽ\;����7��͓����;�<��5=l�d=t-~=�2�=�s=R~R=�#=���<��< %-�P���,U����������轪�����������j�	�����ƽAB��"�7�t㓼p��;��<��5=V�d=(~=o0�=Fs=>zR= #=���<С<�   �   8�\�����0�<:j�m����/���<��\����������@���׆��C�h~ۼ����͈</=��Y=8G�=S= Ǡ=�<�=/q�=��=j�J=��=��B<P>��������%WĽ� �-�8�5��H��NR��S�,�I��{7��p�6!��G3��Vi�T�׼ @͸(�<8�=֗3=B�>=b:5=z�=�
�<��x<��:�   �   h棼l&��� �2�?�v�W�b�g�Dhn�&Nj���Y��;<�h/��ѳ��\ƻpo:<��<Ի>=��~=��=���={4�=��=Ӹ=C��=���=�-g=^`=p�G<\����H�ǵ���I���&�2<L��m�����^�����sa��8�{�{�\���6������ɽ��{���� Ï�(�_<]�<[�<�m�<`�<��Y< �*;�g��   �   �Q�f[��S#�,+�\�)��� ����h]᭼�(<� �8@LX<|��<h	.=��j=e��=�?�=�˿=�o�=�'�=��=���=
0�=�^�=�jy=�t=P�<`�ü��=Iڽ�m�4O���~���������N��>,���Q��7�����:�q���@�Q�½ƽ�)s�T��0�����;(E5<�l0<p��;@���>�`K���   �   ��$���1��2��3'�V����������; zl<p��<��$=:�[=u�=���=[-�=RH�=>�=Dd�=�i�=4�=أ�=J%�=Xƪ=���=<|=��;����c����_i=�2x�������ž�|Ҿ�l־HѾz�þ4׮�/)��Rr���9�#��i���Z��y鼀�V�PEĻࡷ�x�%�\g����ּj���   �   4Q�̅T��gH���-�jp�@i��@��@��;��<4=X3?= �u=<8�=d��=8��=�r�=0��=���=���=��=h3�= >�=��=���=���=��= ��9��.�M�������Z�>����q��Tx̾�j���J����k�AH�~˾�`���Ꮎ��^���$�76�~���V�=��8�������	ȼ���J�"��8?��   �   X�v��Is���]��Y8����o���,���c<���<4�9=�u=qm�=�.�=$��=��=�~�=4�=�a>|�>XF>_] >���=���=`�=��=��
=���n�O��|ؽ��,���r����s������0���K���O�q�����|��O¾�����{�A�<�<��ո�4$w�"]*�h��� ��u��0�~P���i��   �   ���V,��j[m��A��&�t�� w:tI�<4Z=�V=���=�M�=�ؿ=t�=p��=T��=
>->�>�>�>Z.�=���=}�=�I�=Й= ���8f�0b��d8�(U��B����;�\���r����Ϟ������ϾM/��QI���\L�����ν\�����J��&$���M0�N��m������   �   �o-��)�����V��Jڽ���4JB�t��0�'<��=�m=·�=Zg�=�J�=l��=��>��>��>��>U�>��>� >�=��=V��=.ip=��< ?��J�:���*[���D�B�w�����~¤�A\���Y���a������c6}�z�O��$�����4U���d������P��$7��.½�b�|�
�����(��   �   �6)��%��w��~�V ֽ/6����?�`���h�<f&=��h=���=l1�=�	�=�~�=�g >��>Y
>��>w�
>��>�9�=�)�=�0�=P�=�o=��< F���5��涽�V�t�@���r����Ja������͒������\p��Dm��B7w���J� �����\����������4��4̙�JD��C����v���$��   �   �r��g��\�����ɽx���}8�����H<*�=B�X=�r�=V�=�=���=b��=�b>*~>x(>�<>y>x)�=(~�=�-�=�^�=2jj= �<�$E�H�'�a��a��>O5��Sd����>���T.��ѩ���á�V��dĆ�!�e��K;��B�j�ܽ�������ԓ`�P�f����(-��ν/����1�7��   �   $�
�����P������f���߉�@�0�H"���D�;(E�<�;=J�=(3�=C��=Fd�=xF�=z�=��=L>�t>N��=΢�=���=
>�=��=�`=ȵ�<�J�� ��͙���｡�#�(4N�/�s�ĩ���񑾩˔��퐾�Ն�@xo�j�J��m#��	���ϸ�@C��N�F���(��.���S�����'���ѽ~�*��   �   mp罕��:�۽t�Ľa���=�.��뵼`�� �<8�=� S=�ʈ=��=�p�=���=���=T��=FH�=��=��=��=@��=���=�X�=��O=�R�< n�B2 �Y[���<ѽ���P*3�?S��#l�d{�\]���w�'�d��I�j(�8!�!;ƽ�͊� 9������ü Lμ����d?�����ܣ�l!ý]�ڽ�   �   ����f������#���铽��r�Z7��M�U��{I;p�<�=~�K=�=kR�= �=q�=4��=���=���=�J�=�(�=6x�=>b�=�:~=Ҭ3=�X�<@�����X#i�ݲ��r�M���/��tC�.�N���P���H�Ff7�U�������Ž�P��Z�,�l��� w��dz�����H�M�?ɼt!��a�D���鷦��   �   Ŵ��k5��&*��#�����0Bv�VZR���'���４��@����J<���<Ė.=~i=瓎= �=��=�q�=��=.�=>z�=1�=#�=h�N=�L
=P�v<�������
5P�옽��Ƚ+>���Y����8�!�0)!�������+潖�����|�����x����:��O<4��<���<8�< ����ru����hy3�b�e��   �   j�4��Z��u�.����ʇ��n��������q��T���,�����`B�� ��lr�<v�=F�B=�v=���=��=ʞ�=ȩ�=>�=l�y=��I=X�=�ۢ< �];��a�" ���G�Q������AŽ`eܽ�?���޶轭�սa췽w��aK����P�ֻ �><��<��=�]=ns=���<��<�<0����O�� ���   �   |yڼ�#��T��b�����s��A���Lz��mr��[1��䮃��oM�r����n�`2�;�q�<N�=iG=x�e=�]q=Φj=fS=8'-=�~�<06�<@;;HKN��ڼ�#�^T��a�B����������Mv���m���,�����nfM�����ln�pk�;�~�<��= nG=(�e=,bq=b�j=S=,-=���<�?�<��; ;N��   �   H�a�� ���G����Y���DŽ�iܽ�D�[��b��+�ս���{���iK��� ׻0�><P�<�=�X=�n=���<ڭ<P�<�ƭ��Z��"��Ζ4�BZ���u�[����ɇ��l��������q���T���,�t����2�� �۸H��<Ķ=ڠB=�!v==9��=Ѡ�=ʫ�=A �=|�y=��I=<�=��<�];�   �   ��\�Ἀ7P�*��Ƚ*B���[�l��$�!�0,!���ƽ��0������|������x�@A�:�O<p��<l��<0�<@G����u�X��3�T�e�m����7���+���#������@v�6WR��'����X��`����J<��<��.=�
i=K��=C"�=��=�s�=N�=�/�=�{�=�2�=��=J�N=BO
=��v<�   �   @.��� ��&i��߲�+v��O���/��wC�7�N���P���H�i7���������Ž�S����,�p��������z��ᨻ��M�HJɼz!���a��Ď�������\i������n����铽h�r��7� H� �U���I;d%�<�=n�K=p�=�T�="�=�r�=̄�=d��= ��=L�=*�=ry�=[c�=�<~=�3=�Y�<�   �    �o��4 �t]��r?ѽ����,3��AS��&l��f{�E`�t�w���d�D�I�l(��"��=ƽ�ϊ�h9������ü�TμJ���i?��"���ߣ��$ýi�ڽMs� ��G�۽��Ľ?��N>�Z.�t赼@j�� �<ԯ=`S=�̈=��=�r�=X��=H��=���=hI�=��=
��=� �=��=w��=VY�=��O=�Q�<�   �   ����$��ϙ�~��f�#�:6N���s� ���(��̔���ֆ�zo���J�@o#���|Ѹ��D��Z�F���(���.���S�����\)��|�ѽ��w�b�
�ƴ��R��`�ོg��$����0�P ��`R�;�I�<��;=��=4�=���=te�=�G�={�=���=�>Xu>���=d��="��=j>�=��=��`=���<�   �   @FE�P�'�g������P5�ZUd����4���H/�������ġ����Ć��e�cL;�0C�m�ܽ���������`�~�f�<!���.���ν����2��7���B����i�����ɽox���}8�l����<��=�X=�s�=�V�=��=X��=��=c>g~>�(>�<>/y>�)�=X~�=�-�=�^�=~ij=p|�<�   �   @V����5�4趽�W���@���r������a��?���K�������p��ym���7w���J������,\���������5���̙��D����a���v�'�$�,7)�4%��w��~�� ֽ@6��R�?�����(�<4'=x�h=��=�1�=
�=�=�g >��>(Y
>��>��
>��>�9�=�)�=�0�=�O�=�o=��<�   �   0M��V�:�>���[�r�D���w�崒��¤�Z\���Y��wa����������5}���O�	$�����]T���c����>P���6���-½�b�n�
�ҵ���(��o-��)����vV�9Jڽp���IB�� ����'<��=D�m=ӷ�=\g�=�J�=`��=t�>��>��>��>=�>��>�� >��=���=ҍ�=�gp=��<�   �   �E���5��涽�V�J�@�Z�r�޶���`��I���P�������o���l���5w�U�J�������`Z����K����3��	˙�&C����L��^u���$��5)�%��v��}���ս�4����?�`�����<x(=z�h=~��=$2�=H
�=>�=�g >��>1Y
>��>��
>Х>�9�=�)�=1�=,P�=�o=��<�   �    E�P�'�8�����]N5��Rd�C��z���u-��ި���¡�M��^Æ�2�e��I;��@���ܽ��q�����`�h�f�
��'+���ν����Z0��5������������.�ɽ�u���x8�tP%<�=«X=ot�=bW�=4�=���=H��=c>}~>�(>�<>My>*�=�~�=(.�=T_�=�kj=H��<�   �   @ܟ�4��Q˙����#�d2N�)�s�������Rʔ�4쐾GԆ��uo��J��k#����̸�@����F���(� �.���S�κ��$��ыѽ{�Y�<�
�����L����c��܉�P�0�<���u�;dP�<,�;=� �=<5�= �=�e�=�G�=N{�=0��=�>ru>H��=̣�=���=0?�=��=��`=ػ�<�   �    i��, �/X���8ѽ��� (3��<S�!l�a{�&Z�j�w���d��|I�:g(����6ƽxɊ��9�����hü @μ���^?�R��-٣�Ký��ڽ�k�ҭ�_�۽��Ľ�����4�D	.�@۵����(�<�=�S=~͈=)�=�r�=���=���=о�=�I�=6�=l��= !�=���=i��=�Z�=��O=�[�<�   �   �L�����zi��ز��m��J���/��qC���N��P��H��b7������N�Ž�K����,� ��� [�@�y����HxM��0ɼTl!���a�����������wa�������悔�㓽��r��7��9�H�U�`J;(,�<`!=R�K=�=U�=l"�= s�=��=���=n��=�L�=�*�=2z�=jd�=�?~=�3=0d�<�   �   p������+P�瘽8�ȽD8��jV�T����!��%!�\������$潏�����|���@�x� ��:p�O<���<ृ<< ����Ru�\���o3��e�@����/��>$��������6v�dNR���'�D��d��� X���J<���<�.=�i=���=�"�=	�=�s�=��=0�=t|�=}3�=��=8�N=PS
=X�v<�   �   �za�� ���G����@���;Ž�^ܽ�8�(������ս�巽�p���UK�Ԓ���ֻ8?<�%�<��=Ld=z=���<\�<�/<@S��|<�����8�4� Z���u�˚��ć��g��[����q�<~T�z�,�����-�� ظ䂆<��=��B=�"v=2��=��= ��=,��=� �=�y=��I=�=X�<`	^;�   �   mڼ�	#��T�~V�������������o��hg��&������:ZM�4��hBn��;Џ�<��=uG=��e=thq=��j=�S=3-=ė�<�P�<@;PN�`cڼ�#�nT��U����u��,���=s��|k���*������NdM��� hn�r�;��<f�=�nG=��e=�bq=�j=�S=L--=��<E�<`�;((N��   �   
�4�Z�Z�u�ڛ��5ć�0g���}����q��wT��,�������� \Ǹ���<8�=��B=�(v=��=1��=���=���=D#�=�y=��I=�=��< Q^;la�" �t�G�%��e���=Žbܽ=����C��w�ս{뷽mv�� `K�(����ֻ��><��<h�=*^=t=`��<��<�<�����I������   �   �����2���&�����M���5v��LR���'���� ��������J<t��<��.=i=���=F%�=��=(v�=��=F2�=�~�=�5�=���=l�N=HW
=0�v<������ἰ+P��瘽��Ƚ�:��@X����`�!��(!�r������*�5��� �|�`��`�x� ��:P�O<���<x��<��< v���mu�X���v3��e��   �   ���d��������䓽��r�b7��5�ТU� MJ;�5�<�&=��K=��=�W�=�$�=Pu�=��=���=@��=LN�=h,�=�{�='f�=�B~=>�3=�i�< ������i��ٲ��o�mL���/�&tC���N��P�H�H�f7�$��h����ŽWP���,�ܱ���u�`_z�����P�M��=ɼs!���a�R��������   �   !o����۽ʏĽ*���f6��	.��ٵ� ��8.�<L�=r
S=wψ='�=�t�=���=H��=p��=0K�=��=���=�"�=.��=ҙ�=\�=�O=�_�< �g�(, ��X���9ѽ���_)3�T>S�G#l��c{�]�h�w���d��I��i(�&!�;ƽk͊��9�P���0ühKμH��d?�z��vܣ�� ýa�ڽ�   �   ��
���_O���ཊd��݉�>�0����|�;�S�<d�;=�!�=�6�=~�=<g�=(I�=�|�=h��=_>v>X��=��=Е�=I@�=��=��`=$��< �������˙�͝���#�3N���s������񑾌˔��퐾�Ն�-xo�]�J��m#��	���ϸ�1C��&�F���(���.���S�]����&����ѽ~����   �   ������"���u�ɽdv���y8�h&<��=�X=5u�=@X�=!�=���=(��=�c>�~>')>5=>�y>�*�=��=�.�=4`�=Dmj=D��<`�D�~�'���з��N5�?Sd�������<.�������á�N��]Ć��e��K;��B�d�ܽ���������`�.�f����
-���ν����p1��6��   �   �6)��%�mw�T~���սX5����?�D���8�<�(=��h=ӹ�=�2�=�
�=��=�g >�>oY
>��>ɒ
>�>T:�=|*�=�1�=�P�=No=���< :����5��嶽oV�6�@�q�r����<a������ƒ������[p��Am��?7w���J�������\����������4��(̙�>D��0��ޞ��u���$��   �   ]���i��e���ȃ�
�]���.�O=���3����� �<;��=�=�=��=v4�=!�=XF>�'>�>qS>�>��>�a>�:�=0�=�=Je�=�4b=�X�<`Jy;��ؼj�p�T廽�����޸1�.@�"E�Z;@���2��[����ݽߒ������Ky���G���E���::�Rc�JȄ�n�������   �   �6��[����M�����MY�q
+��������~�
�  S;�I=Pm~=�W�= Y�=\�="7 >�>6�
>8.>2�
>b0>L� >$K�=��=��=�ɘ=�]=���<`j;�ּ�l��X�������p�-���;�Fr@��;���-����ր�t�սج��T���̈́�L2��∪��۽����15�]������B��^����   �   X)��8���f���}r�1	L��� ��	�kߐ� ���;��=Եw=2��=#��=��=<��=��>��>ũ>+>�1>n�=�_�=�=�8�=q��=LuP=0��<�J,;l	м��a�s���A�؁���"�F/��3�h�-��� ��\����e]��aD��f�{���e���u��薽f�Ž�E���&�|SM�!zq�򞇾v����   �   �����%���yu���Z��38�^Z�?�ѽtÂ�Ȱ�@˘;8c=X�j=�ɞ=n��=�	�="��= *�=^�>�>$� >���=~��=<�=�`�=Lɣ=�O�=6�7=�f�< �9�Wͼ,�S�d��a
Խ� �L���"���f�����&o�.ɽC����%u�^bB���-�}<��9p������yݽڙ�� 4�N�U�GPq�b����   �   z�d��Fa�6�S��9=�! �D���3@���g��ʼ i�;�b�<�T=&�=A�=���="a�=���=8��=���=��=��=��=���=RS�=�Č=��X==܄<�����ؼ�2H�;����̻�l�߽����ȱ��7�̈́��9@�I������ �h�.�&��'񼸏˼����R!��Co�����6�^o2�^�K�q]��   �   �9�D�8�r�.�ԩ����*5ؽ|���D�M��B�� �:Ģ�<@�2=�z=���=.�=�E�=DN�=r��=�T�=��=���=���=�ף=|��=l�Y=�=H��<`�; 
U�ԁ���F��ޅ��줽WM��۱Ͻ�׽�Bӽ�Ľq骽%���H�M��r�����0�� ��� j�����2��[f��x��(����W�!��1��   �   �t�X��D�
�d��`�ݽē��j����@��Ҽ�2����d<Pd=fE=V	�=fۘ=z4�=�]�=�п=sN�=X�=`��=v:�=�k{=�DC=��=���< �";8�I�@!ټ�B#���U�^-������L꠽�����u�������]���Na�*�#� �ļ`� ��;@�T<��<`>m<p8�;Y��q߼TNK��(����Ľ�m�����   �   ��˽[Խ��ҽP�ǽN��[��Gڀ��XD�J��~�� ������<� =v�9=N^l=S9�=��=�@�=3̜={n�=���=��V=�=Ȃ�<���;���l��-<�į_���z�1���]���{���k��rZw�V�TB)�\�H�[�@_�:��{<���<�Y=�A=`8=��<��<�`�:ؐ��ؑ�Am����V ���   �   D�����������S��Hї�8L��|����]��i3�0��x�������8�-<�%�<*�=n�E=Z�b=��o=fk="�S=*�*=�i�< G< ���P��B!��Z�3�������q����U��`җ�dL��Y{��ķ]��e3�8�������ˇ��.<|0�<F�=N�E=�b=��o=Rk=p�S=�*=�v�<�'G<�گ�<@���9!���Z��   �   H��(<��_���z�􉆽�]��)}���m���_w�,V��H)�H�8�[����:p�{<p��<�T=�<=.3=���<��<�}�:Ԡ�����|Jm�� ��>%��j�˽S_ԽS�ҽ�ǽ�O��L��Sڀ�tWD�~��w�� @M�蒂<� =:=�bl=};�=��=C�=hΜ=�p�=��=r�V=�=��<�/�;���t෼�   �   ��I�|ټ�@#��U��-��碓�^젽Y����x��!���`a���Ua���#�l�ļ ��_�;��T<��<()m<�	�;(s���߼�VK�|-����Ľ
s���@w����\�
����ޓݽX���񋽬@��Ҽ���`�d<�g=0E=@�=Cݘ=P6�=�_�=�ҿ=PP�=`�=���=�<�=�p{=VJC=4�=|ɐ< �";�   �   �(�;�U�����ޥF��߅�z�O���ϽV׽[FӽkĽ�쪽s���L�M�jx�ğ��x������p�����*9�"cf��|��ל�c��!���1�ʼ9�Ŧ8���.����
��*7ؽ�����M��A����:0��<��2=ָz=I��=��=EG�=�O�=���=hV�=���=~��=b��=�٣=� �=��Y=�=`��<�   �   ߄<@𒻤ؼn4H�Č���λ��߽â��z���9�7���|C�@������� �h���&�,0�,�˼����W!�dIo�H�����,9��q2��K�
]�	�d��Ha�\�S�T;=��" �]����A��<
g�d�ʼ o�;�e�<�T=9�=�B�=���=@b�=܇�=`��=���=�=��=���=q��=�T�=	ƌ=L�X=:=�   �   �g�< V�9�Zͼv�S��e��Խ(� ����4$�c�����
���q��0ɽ-����(u��eB���-���<� >p�患�G|ݽ|���"4�\�U�qRq�~��������&���{u�.�Z��48�O[�~�ѽ&Ă�����͘;d=��j=�ʞ=9��=�
�=���=�*�=��>��>�� >���=p��=>�=�a�=5ʣ=�P�=D�7=�   �   ���<`;,;�м�a��t���C��� �"�:G/�3�s�-�t� ��]���^��kE��` |���e�@�u�ꖽ�Ž�F�%�&��TM��{q�����D���"*�����Bg���~r�
L�Z� ��
��ߐ�l �p�;z�=��w=���=���=���=���=��>�>�>a+>�1>�n�=J`�=��="9�=���=|uP=�   �   ��<`�i;Tּ6�l�"Z��\������)�-�<�;��r@�'�;���-� �����սOج�8U��΄��2������۽F��t25��]�
����B��Ɍ���6�������M�� ���Y��
+�e���'���r�
��S;^J=�m~=!X�=`Y�=��=>7 >�>O�
>M.>L�
>|0>^� >HK�=��=��=xɘ=��]=�   �   0V�< 4y;$�ؼ�p� 滽t���X��1�,.@�,E�D;@�ɘ2��[�Ɔ�6ݽ7���n���/�x��TG��vE���5:�Sc�LȄ�k������T���[��e���ȃ�ܞ]�Y�.�=���3��,��@�<;��=�=�=��=|4�=!�=PF>�'>�>aS>�>�>ta>�:�=��=��=�d�=t3b=�   �   Ъ�< j;�ּn�l�{X��r��������-���;��q@��~;���-������Ես�֬��S���̄�1��Ň����۽,��015�Q~]�=���B��⋛�6��ֱ��M��9��VY��	+�z������� �
�`"S;�K=�n~=�X�=�Y�=��=R7 >�>X�
>[.>T�
>�0>p� >nK�=��=��=�ɘ=��]=�   �   ���<�q,;<мΩa�wq��@�Հ�ܬ"��D/��3��-�� ��[����Z��B�� �{���e��u��施d�Ž�D���&�RM��xq��������d(��B���e���{r�}L� � ����ܐ�h����,�;8�=��w=n��=*��=��=��=��>��>�>u+>�1>�n�=�`�=��=�9�=}��=�wP=�   �   �n�< ��9�Nͼ,�S�ba��sԽM� ����� ����~������k�-+ɽ����u��\B���-�x<��4p��}��nvݽ$���4�-�U��Mq�"���L���=$��fwu� �Z�J18�?X�d�ѽ�����㼀��;�g=~�j=�˞=���=<�=\��=+�=��>��>�� >���=���=��=eb�=�ʣ=�Q�=�7=�   �   ��<@Ò��ؼ�+H������Ȼ�L�߽H�������5�5����;����&�����h�^�&�,񼼃˼ ���L!��<o�E����转4��l2���K�n
]�[�d�nCa��S��6=�> ����s;��j g���ʼP��;o�<f�T=y�=�C�=���=�b�=2��=���=���=T�= �=���=���=zU�=�ƌ=��X=�=�   �   0O�;H�T�Dq��l�F�څ��礽yH��ܬϽ�׽�=ӽ�Ľ�䪽������M� k������0���P6�X�+��Sf�t�����B�!���1���9�ʠ8��.����r��K/ؽ���d�M��0��@�:<��<��2=��z=I �=g�=�G�= P�=<��=�V�=���=���=ʷ�=^ڣ=J�=��Y=l=���<�   �   0�I� ټ�8#���U�-(��S����䠽D���Ap��U����X���Da�ҵ#��oļX���ņ; U<$��<Ym<�o�;;�,a߼
EK��#���Ľbg��� q������
�d����ݽo���zꋽ�@���ҼP魻�d<�k=�!E=<�=ޘ=�6�=�_�=�ҿ=�P�=��=���===�=�q{=�KC=2�=ϐ<�6#;�   �   ���"<���_���z�����aW��v��f��xOw�f�U� 8)���弸�[��m�:��{<T�<�`=TH=�>=l�<T��<�d�:�~������5m�������̀˽�SԽ��ҽ?�ǽ:G�����	Ԁ�<MD�N��j�� ���(��<d = :=.dl=�;�=5�=^C�=�Μ=q�=m��=2�V=��=ؒ�<�>�;X���ٷ��   �   9���|�Q����O��c̗��F���u����]��Z3��v�ؠ������ 6.<H@�<��=�E=t�b=�p=~k=�S=�+=��< JG< ���+���-!�8�Z�����V�����L��wʗ��E���u��n�]�0^3�p{�ȫ��`��� .<�3�<~�=.�E=��b=6�o=�k=�S=��*=�w�<H+G<�Я��<��27!���Z��   �   ��˽�XԽ�ҽ��ǽ�I��q���Ԁ��LD�^�\d��  p�ȣ�<z =>:=bil=�>�=��=�E�=8ќ=�s�=H��=d�V=ʍ=d��<p|�;����ɷ�0
��<��_���z�W���W���v���g�� Tw��U��>)��
��[����:��{<\��<lZ=>B=�8=��<��< r�:p���ؐ��?m�������   �   �s�j���
�y	��؍ݽ�����닽�@���Ҽ�٭���d<`o=&E=X�= ��=�8�=b�=տ=�R�=��=X��=�?�=�w{=�QC=��=(ܐ<��#;@�I��ټ�4#��U��'������1栽S���s������H\��HLa���#��~ļ��@��;�T<���<�?m<�:�;xW��p߼�MK�q(��R�Ľ�l�u���   �   ��9���8���.����:���1ؽш��0�M�t1�� 	�:���<@�2=��z=��=�=�I�=�Q�=�=�X�=Ą�=���=���=�ܣ=��=� Z=�=�ɰ<�s�;��T��k��ޚF�څ��褽J��7�Ͻ�׽ Aӽ�Ľ�誽����b�M�@r�����ؙ������g�,����2��[f�lx��ߗཡ��!���1��   �   �d�Fa���S��8=�  �����l=���g��ʼ���;�p�<�T=��=�D�=���=d�=���=��=j��=�	�=�	�=���=���=wW�=Ɍ=��X=x=��<����� ؼ�*H�Ǉ���ɻ���߽������F7�����?�����������h�ذ&�0'�L�˼����R!�^Co�Ѳ�����6�=o2�+�K�']��   �   x���`%���yu��Z��28��Y�E�ѽA���T����;Ph=n�j=f̞=̈�=$�=T��=,�=h�>&�>C� >��=��=�=�c�=�̣=S�=��7=,t�< 9�Kͼ��S��a��CԽ� ����("�w����{���n�l.ɽ���<%u�.bB���-� }<��9p�o���jyݽϙ�� 4�8�U�&Pq�J����   �   D)����tf��\}r��L�%� �`�ސ� �`'�;8�=�w=ˉ�=���=���=���==�>X�>r�>�+>g2>�o�=�a�=��=�:�=���=�yP=���<��,;�м�a�{q��x@�J����"��E/��3�9�-�b� ��\����D]��LD��J�{���e���u��薽X�Ž�E���&�lSM�zq�螇�h����   �   �6��P���{M�����Y�,
+�t���R����
�`S;�K=�n~=�X�=�Y�=�=z7 >&>��
>�.>��
>�0>�� >L�=��=��=�ʘ=J�]=��<@4j;ּV�l�!X��S������:�-�_�;�(r@��;�v�-����̀�g�սج��T���̈́�F2��ވ���۽����15�]������B��Y����   �   �
E��H����޾���
r���m��|'���ν��<� >9p=U_�={��=Ȓ�=$�=�i>��	>�a>�
>d>� ><��=H3�=L"�=�~�=_Z�=*�Y=��=��<p��� 7Ǽ�	1���t��l��.ͤ��-��0�-������V	a��MD�=�ĤU�(w�� yý� 
���=��.{����)����߾�W��h>��   �   Me����]g�˓ھ�F��6M��5�h���#��vɽ�'6����:H=�Z�=g�=Bz�=���=R�>h�>>
>�>��>XW�=�[�=T��=f�=���=eӉ=�_Q=�	=�Oo<0|����Ǽ:�.�@�o�j����k��v��k���Y�� �|�$V�v�9�DE2��pJ��T��o������8�3*u����(�����ھ�S����   �   �\��3N��tN���;XP���>���Z���u����"�@Zw;hY"=��=�ƹ=� �=�(�=�>��>xC>�>��=��=4v�=>��=2�=S;�=��w=P�7=�F�<��.<���d�̼О)��3c��I������;�����������/\�ZF6�Tg�P����)���f����n��M*�βc�.,��7�����;
��|���   �   \g�1�ܾ�~Ͼ'H���m���V���D����"򣽌c�p��;(0'=V��=���=<��=.�=���=R��=[�=,��=0��=x��=�x�=��=�=��=��F=^�
=�ٙ<�8Y;8/F�l#ܼ2�$�ZR���r������ۀ��o�
BP�^�)����Ӽ��üD�켴�.��ԇ�!�ͽ����rH����r��?����*ξ5Dܾ�   �   �@þϸ��g+���͡�o��JL`���)�i�꽚M���>̼��7<�)=���=^[�=ٿ�=���=���=xu�=�O�=���="^�=�M�=���=vr�=�m=v�5=<��<�r�<0N�;0��4���(F ��7&��8C���T�4�X���M� e5�H����ּ�U���i-�����hR�tTͼdq=�%��9C��%�._Y�(���X�������`���   �   �����+��z㕾�͆���f�8�:��G�=^��N�\�����d<�Z&=��=�T�=���=V/�=�P�=�m�=�=���=��=�e�=~:�=��E=B
=D*�<0��;��ʻ���ּ��
�@V#��P4�|�<�\�;���/�R���U� ڟ��j� �L�P7�;h<0$�;�J��`ྼ��K�ƙ��<���r+�(\X��Ѐ�S��������   �   ��~�@|��`n�84W� �8�i��%��|�-���F���o<�&="�h==��=�ɪ=���=�=�ǽ=b��=Ǹ�="R�=�HW=6�=p�<`C%;��U��ټd��bp;��]Q��d\�t}]�֦U�ΫE���-����zѼ��s� �b� ��;��<i�<�T�<��<���<�:�:5��rM�`	���x����!�x�D��a��u��   �   J=��=��w4��W$��r����&���JPv�:�������I<�{=Z�F=�}=i��=T�=r�=���=�=H�l=�r.=@��<���;�������L�[�f͊��@���w�����i���˙������/c�j�1�p���@Ç��L,�8�4<G�<�=�\+=�:=d�5=,�=$��<0 �;������7��M��Lٽr�	��e"���3��   �   $�����.�����Խ�����'���jI������7���;T�<�="�I=*�l=��=�y�=~�m=��E=�u	=h`k<P�����o�x#���ѽ(�
����1�ϷｧԽ����f)��rlI� ����7�p �;��<�=��I=��l=��=|�=d�m=��E=Z|	=�k<[�F��2o���A�ѽ1��   �   @;��or��~�������,ș�ѣ���-c��1������Ǉ��{,�xs4<�?�<�=�X+=��:=��5=�=��<���;������7��S���Rٽ�	��i"���3�2=�P=�{4��Z$�*u�&�齟���8Sv�h������J<�}=ԱF=Ϊ}=���=�=t�=պ�=��=*�l=~y.=��<�=�;X�������[��Ǌ��   �   ���bh;��VQ��_\��y]���U�H�E���-���܀Ѽ��s� c����;d�<�`�<L�<,��< ��<�r�:�C���zM�������!�\�D�4�a�8�u�֕~�Q|�Odn�r7W���8� ��(��𚽚�-�P�F�@�o< (= �h=_��=
˪=��=��=[ɽ=���=G��=U�=HOW=��=,�< �%;kU���ټ�   �   ��ʻL銼��ּ4�
�.T#�:P4�.�<�@�;�/�ș��]�(⟼`{� �]���;0�<`��;0t���쾼�K�(���v���u+��_X��Ҁ�l��� ��#����-��_啾`φ�Z�f�p�:�nI��`���\� ���P�d<f[&=�=�U�=���=�0�=4R�=*o�=��=���=4�=/h�=t=�=t�E=,
=`8�<0&�;�   �   �{�<0m�;���t���fE �8&�:C��T�N�X�\�M��h5�$��T�ּH]���x-�H��hyR��]ͼ�v=����EG�"�%�bY�Θ���Y��y����b���Bþ����1-���ϡ��p��lN`�n�)����O��B̼��7<*�)=��=�[�=���=���=���=�v�=6Q�=j��=�_�=�O�=:��=�t�=�m=��5=D��<�   �   0�
=,ޙ<`QY;�,F��#ܼ:�$��[R��r�/���i݀�J�o�VEP�� *����$Ӽ��ü���~�.�	ׇ��ͽj���tH������Ѯ���,ξ�Eܾi�� ݾW�ϾI��o��zW��t�D����i�e�p��;60'=���=��=���=��=���=(��=\�=H��=p��=���=Vz�=��=��=d	�=�F=�   �   ��7=|H�<8�.< ����̼�)�j5c��J������~�����������1\�RH6�<i�@���)�$�f�����p�O*�P�c�-��@���;B�����8^��dO���O���;#Q��3?���Z���v����"��Sw;jY"=�=ǹ=� �=>)�=R�>ȩ>�C>>��=ī�=&w�=>��=3�=N<�=J�w=�   �   �_Q=�	=No<Ё��� ȼ��.���o�*���Xl��.���k��Z����|��V��9��E2�nqJ�VU���o��~����8�+u�����������ھ�T�l���e����g�?�ھG��~M����h���#�8wɽ(6�@��:l=�Z�=��=pz�=���=l�>��>]
>�>,�>�W�=�[�=���=qf�=§=�Ӊ=�   �   N�Y=��=�<උ�$9Ǽ�
1���t�m��fͤ�	.������c����a�(MD�R=�8�U��v��yý� 
���=��.{����5�����߾�W��g>��E�qH����޾����q����m��|'�5�ν�<� �>9xp=o_�=���=В�=$�=�i>��	>�a>�
>�c>� >��=3�="�=�~�=Z�=�   �   �`Q=�	= To<ps����Ǽ��.���o������j������i��aX��Ь|��V�8�9�C2�~nJ��S��n��n����8��)u���������_�ھRS�����d�W���f��ھF���L��/�h���#�tuɽ^%6��:�=C[�=��=�z�=��=�>��>k
>�>2�>�W�=\�=ޥ�=�f�=T§=�Ӊ=�   �   t 8=�L�<��.<�����̼\�)��/c��G������I�����������+\��B6��c����r�)��f�D�l�L*�f�c�\+��B�����;���4��[���L��%M徥�;3O���=��0�Z�n��r����"���w;D\"=�=�ǹ=z�=�)�=v�>�>�C>>��=��=^w�=���=��=�<�=��w=�   �   � =d�<��Y;PF�`ܼ��$�rTR���r�ڊ���؀�b�o��<P�6�)� ��pӼ\�ü<���.�9҇�Gͽ���pH����������F)ξlBܾ�e�X�ܾ}ϾxF��pl��4U����D������]���;>4'=��=��=z��=V�=���=n��=H\�=z��=���=&��=�z�=��=U�=
�=��F=�   �   t��<���;�� ����> �@0&�>1C�T�T� �X���M�X^5����P�ּ(J���S-�X��pSR�<IͼLk=����+?�P�%�d\Y�����@V�������^���>þ����G)���ˡ��m��I`���)�w��jI���0̼�8<��)=���=>]�=w��=n��=���=�v�=|Q�=���=,`�=4P�=���=Zu�=$m=@�5=���<�   �   p�ʻ@ኼ��ּ��
��L#��G4���<���;���/�P���F＀˟�pO� h3� h�;�&<�S�;����Ҿ�4�K�V�������n+��XX��΀�)�����������n)��)ᕾ�ˆ���f���:��D��X����\�4⏼��d<�`&=��=�V�=���=81�=�R�=�o�=�=���=v�=}h�=�=�=f�E=r
=<�<�8�;�   �   l��Zd;��QQ�NY\�2r]��U���E���-�����iѼ�s��Sb��!�;"�<�u�<a�<��<l��<��:T%���hM����r����!�z�D���a�Fu�ƌ~�n|��[n��/W���8������蚽(�-��F���o<l-=��h=ƫ�=	̪=˕�=6�=�ɽ=Ն�=���=EU�=�OW=f�=�-�<`�%;�cU�Ħټ�   �   �9���p����������ę�����T$c��w1����<�����+��4<<U�<$=(c+=�:=`�5=x�=���<�=�;����n�7��G��-Eٽ��	�qa"�O�3���<��=�s4�IS$��n���f���@Dv��|�(���J<΂=��F=��}=���=��=|t�=/��=��=��l=�y.=$��<�B�;�������2�[��Ɗ��   �   ������-�Q�｟ Խ=���n#���aI�4�����6��b�;�)�<�=�I=��l=��=�~�=Z�m=��E=��	=��k<�4�8��� o������ѽ��������*�ʪ��ӽ��!���^I�`���8�6��S�;H$�<4=�I=��l=m	�=�|�=�m= �E=�|	=H�k<PY�¸�vo������ѽ;��   �   �=��=��v4��V$�pq�^�齅���JHv��~���X!J<��=<�F=��}=���=��=�v�=���=��=��l=�.=`�<���;�u��|��.�[�Y����3���j��呬�*���������!c��v1�����������+�ؑ4<M�<�=r^+=��:=�5=��=��<P�;З��j�7��M���Kٽ?�	�Ze"�e�3��   �   -�~��|��_n�Q3W���8���"㽅뚽J�-���F�H�o<j.=��h=���=tͪ=f��=�=�˽=��=(��=HX�=�VW=4�=L?�< }&;P<U���ټ���[;�rIQ�XR\��l]�t�U���E���-����nѼ�s� �b� ��;L�<�k�<�V�<��<���<@F�:|4���qM�>	���x��j�!�T�D�ؚa���u��   �   ֤���+��6㕾Z͆���f�5�:��F��[����\�x揼��d<�`&=��=�W�=ƥ�=|2�=.T�=,q�=�=��=��=Pk�= A�=j�E=
#
=�K�<0y�;�Fʻ�Ҋ�ܟּܾ
� I#�nE4�ּ<�v�;���/�l���N０ԟ�c� �G��>�;�< (�;�G���߾���K�����$����q+�\X��Ѐ�A��������   �   �@þ����7+���͡�0o���K`���)�n��vK���5̼�8<§)=��=�]�=A��=d��=��=>x�=�R�=^ �="b�=pR�=��=x�=m=f�5=���<<��< ��; ������< ��.&�B1C���T�b�X��M�Pb5�<����ּ�S��g-����gR��Sͼ:q=���"C��%�&_Y�#���X��u����`���   �   Ng��ܾ�~Ͼ�G���m��PV��t�D������F`�Щ�;�3'=��=l��= ��=�=���=b��=`]�=���=��=���=x|�=��=�
�=Y�=t�F=�=X�<��Y;�F��ܼ��$��TR�F�r�����~ڀ��o��@P�`�)�b���Ӽܹü��켄�.��ԇ��ͽ����rH����o��<����*ξ*Dܾ�   �   �\��'N��cN���;7P��h>����Z�~�&t����"��}w;�["= �=�ǹ=��=*�=��>5�>3D>�>��=��=�x�=���=�=]>�=��w=�8=�R�<p�.<����̼Ě)�"0c�XH��r���f���穏�L��/\��E6��f�����)�l�f����
n��M*�˲c�+,��4�����;��w���   �   Le����Vg󾾓ھ�F��#M���h�z�#�{vɽ�&6����:`=+[�=��=�z�=��=��>��>�
>T�>z�>vX�=�\�=���=�g�=Aç=�ԉ=�bQ=�	=�Zo<�g��T�ǼB�.���o�����	k�����j��LY��ܮ|��V�J�9�&E2�vpJ��T��o������8�/*u����'�����ھ�S����   �    ;O�F4K��x?��.-�*��k��)Qþ�d���tD�%齤:H���e;��6=>�=�'�=���=x��=v>m>��>�r>���=b��=<��=�s�=���=��=���="uS=VM$=D1�<d�<p�< ���"ѻ �"���3��$�ps�0�������z�db���a�~����j�Z�;���֠Ǿ��������Z-�z?�0,K��   �   �cK��qG���;�!�)�y9�Ӛ�h���Z����?�)��h�?��:�;&R9=ǧ�=���=���=�=oO>��>��>�z�=���=*��=���=)��=H`�=�o�=$t=F�F=��=(b�<xσ<`�; �S��ϻH��$�h��з׻P����1ٻ��X���>,V�>�������6U� ���bþb���ɧ��*���;��bG��   �   >@��<���1�ĉ ���
�	��
!������F�2�h_нT0'��1
<�@=/��=ȅ�=$��=���=q� >�>d.�=��=��=v�=n��=���=D��=@�t=�NI=��=�s�< ڝ<0'.<��P;�h-�@%Ի�y�0U��ť�@�� �T�����pV뻜詼�5�LZ�����EE��!��"��$��W��c �gd1��c<��   �   �.���+�I�!����Y��� о�9n�"���W���E��b<�YK=�f�=��=d��=� �=$��=d��=�H�= t�=_��=6�=@z�=�l�=�U=X�(=���< T�<�^< ��;��4:`\t���ջ����`yջ��t� ��9 /�;�3�;���;`�;p�#��"���������c,��u�@ꣾ
�Ͼ�n��\��!�=+��   �   ]��M��;�Y���<#ܾv����`�L�2Y���$���@��<�)V=��=^��=�D�=��=j��=��=*�=��=�{�=�C�=x�S=�Y=4=�< (_< �;��n��1�x�T���s�8Cv�P^��&,� �û >e����;�H<�f�<�̒<Yi< w;`zz�]6�LP�������M���ڲ�Ĝپɩ��j]�����   �    �����~��K�վ~E����6�i���'��,׽h�Z������<@L^=�j�=�W�=���=4X�=�i�=dJ�=�F�=|��=�]=.�=���<@�K;��@��ļ���HN�b?)�ܼ&����j��p�ͼ����"���� ;��<<�W�<(&�<��<���<���<@yT;���(	j���ѽ�� ���`��$������\�Ѿ�6�U/���   �   p:;?�ɾ�Q��̡��ƶ��7oq�ԅ9�6D���t���/:h��<R�`=]��=�\�=Y�=��=���=�n�=�z=@h1=�Ⱥ<�c\:�s���+���s��֕�lҧ��)��_1��J��y����g�&5.���㼈�R� ��:��x<$k�<�=�q(=��)=�=Ta�<���:�㼙Ն���T�'�G�`�@K��U����1��-�Ǿ�   �   �8���=��ީ���s��@b�,8�DS�=�½Z�e�֭���<��
=dO[=���=�7�=T/�=Ui�=��=q\=dV=�V:<�<y�2�.�����ǽ���2
����E�R&����mཬA������*z5�0 ��lb�<�h=��3=�T=*�_=�JS=�5,=!�<�4�:@^�ԉ�'�ཌྷ���kL���u��݋�gK���   �   ��_�~B^�%�R���>� 6$��j���ɽSሽ+��Y��&i<�E=2dL=��x=`�=T��=�Xv=>_C=��<��;pӼ�t��Ľ2����'�*KC�deV��_��G^���R���>��9$�~m���ɽc䈽�.�@b��#i<`F=�eL=��x=��=��=(]v=�dC=d-�<�c�;`�ҼT�t�7	Ľ��#�'�FC�$`V��   �   Z�~A�x"������'=��N݈��u5��跼���Lb�<�g=��3=�T=��_=�FS=�0,=��<�C�: q�Jډ�&�ི���pL���u�����[N���;���@������v��Ib�v!8��U���½d�e�Dܭ���<F�
=(P[=[��=�8�=�0�=Pk�=C��=8w\=�]=@{:<Py�L	2����ǽ[���
��   �   f˧��"��I+��������
g�F0.����X�R����:��x<�g�<|
= o(=@�)=�=$W�<��:�㼃چ��	��'���`��M��,���5��\�Ǿ�=;V�ɾ�T��]��������rq���9�OF����4"� /:���<��`=爔=v]�=VZ�=n�=���=qq�=X�z=�o1=�ں< _:�[���+��s��ϕ��   �   2��D�@6)���&�8z����$�ͼh	������� ;��<<�S�<@!�<@��<���<���<�)T;8���j���ѽ�!�r�`��&������9�Ѿ�9꾋2��� �Υ��d���վ�G������i�.�'��/׽|�Z�H�����<L^=k�=�X�=���=�Y�=<k�=~L�=pI�=��=*�]=��=l��<��L;�t@�(�ļ�   �    A�;�kn�����T�h�s�7v�^� $,� �û >f� ��;��G<,b�<Tǒ<hLi<`�v;��z��b6��S�������M�����*ܲ�)�پu����^���������m<�����Q%ܾ.��P���n�L��Z�
�� �����<4)V=	�=Ԑ�=^E�=��=���=���=,�=J�=p~�=�F�=��S=�a=PM�<�H_<�   �   D��<�]�<��^<��;�A5:�@t�@�ջ�����~ջ�u� �9� �;@#�;���;`�;��#��&�ꮃ�����e,�\u��룾��Ͼ�p��0]��!�K>+�E�.�6�+�j�!�����Z��"о����:n�`��oY���G�@	b<�YK=�f�=:��=��=B�=��=���=.J�=�u�=`��={�=�|�=do�=��U=�(=�   �   �QI=R�=�x�<�ݝ<0,.<��P;�f-�0(Ի�|�P]�pϥ���� hV��┺�d��쩼f5�\����4GE��"��>��w���jd �Je1��d<� ?@���<�f�1�z� �v�
����!��>����2��`н�1'��.
<��@=<��=���=|��= ��=�� >�>R/�=��=B�=��= ��=���=���=��t=�   �   Pt=J�F=F�=c�<�σ<��; �S���ϻ���$������׻����7ٻ��X��⼜-V�*�������7U�� ��{cþ!���5��b*�y�;�cG�ydK�rG���;�z�)��9�H���h��7[����?�����?��9�;.R9=ԧ�=���=���=:�=�O>��>ޫ>t{�= ��=���=X��=܎�= a�=Wp�=�   �   D��=xtS=�L$=�/�<��<��< 铹 &ѻ8�"�H�3��$��r�@�㻠����z��a����a�+~������Z�R����Ǿ��������Z-�!z?�2,K��:O�=4K��x?��.-���k��Qþ�d��ZtD��$��9H�`�e;�6=3>�=(�=���=|��=zv>j>��>�r>���=H��=��=�s�=���=͟�=�   �   �t=�F=8�=xe�<�҃<p"�; TS���ϻ0
��$���Ъ׻�����$ٻ@�X��⼢*V�^���d��T6U����hbþج��w���*���;�bG��cK�qG��;���)�9����g��dZ����?�����?��I�;�S9=\��=O��=��=f�=�O>�>�>�{�=0��=���=p��=���=,a�=�p�=�   �   �RI=��=|�<D�<�6.< 
Q;�.-��	Իxl��;�@����S� R��V��@@��⩼�5��X�����DE�� ��2���澭��b ��c1�	c<�&=@�)�<���1�� ��
�������������2��\нH,'��>
<��@=>��=���=���=Z��=�� >�>r/�=�=d�= �=.��=㌦=H��=t�t=�   �   p��<�a�<�^<���;�*6:`�s� �ջ�e���Qջ��t� �9pP�;0S�;`��;�,;�p#���$������b,��u��裾p�Ͼ�l���Z�`!��;+���.���+�
�!�w���V���оY���n6n����UT��l@�`b<�]K=#h�=8��=���=��=f��=���=XJ�=�u�=���=��=}�=�o�=��U=�(=�   �   �O�;�Fn�����T��s��"v�(�]��
,���û H_� 	�;xH<�p�<֒<(ki<�Lw;�ez�:W6��L������M�R���'ز���پ:���\����������9������ ܾG���D�L��V����ȩ����< .V=�
�=��=.F�=|��=��=���=>,�=z�=�~�=�F�="�S=\b=dO�< N_<�   �   0���A�3)��&�~u�*����ͼ����0����l;��<<�c�<,1�<t��<���<,̞<��T;����pj��ѽ�� �4�`��"��������Ѿ�3�,��e �c���O��P�վ�B�����%�i���'�5'׽<�Z�`m�4��<`Q^=�l�=�Y�=���=&Z�=�k�=�L�=�I�=��=��]=�=���<@�L;0p@�D�ļ�   �   mʧ��!���)�� ���|��Rg�*.������R����:x�x<x�<�=xw(=�)=�#=8m�< ��:����І������'��`��H�������.����Ǿ7;��ɾ�N��ʞ�����ejq���9��@�:y���� �1:���<��`=Պ�=�^�=C[�=	�=��=�q�=Ҏz=Xp1=�ۺ<�#_:�Z��+��s��Ε��   �   � ��@��!�����ཌྷ:��Rڈ�o5��ڷ�`%��q�<�o=��3="T=��_=,PS=�;,=p.�< /�:�K��Ή�K��}��gL�P�u��ڋ�LH��z5��|:��Ϧ���p��b��8�9O�S�½��e��­��<|�
=\U[=3��=�9�=�1�=�k�=���=�w\=b^=�|:<�y��2�����T�ǽ���x
��   �   O�_�B^���R���>�$5$��i�	�ɽUވ��$�x>��Bi<"M=�kL=�x=j�=ȿ�=�bv=,kC=4<�<Щ�;P�Ҽ��t��Ľ���T�'��@C��ZV��_��<^���R�y�>�N1$�\f��ɽ�ڈ���3��Gi<�L=JjL=��x=��=꽇=:^v=�eC=x.�<�f�;��Ҽ�t�	Ľچ� �'��EC��_V��   �   �8��u=������^s��jb�.8�R���½��e�Hʭ�X<��
=�U[=���=%;�=V3�=�m�=&��=�}\=�e=Р:<��x�L�1�|���P~ǽ;���
�`���<������.�c5��^ֈ�fi5�tӷ���$r�<�n=��3=z
T=8�_=LS=�6,=X"�<�B�:�]�Zԉ��ཀ���kL���u��݋�LK���   �   W:;�ɾ�Q������o���jnq��9�)C��|������0:(��<��`=H��=�_�=�\�=���=,��=Wt�=&�z= x1=��<��a:�B����*�؜s�qǕ�ç����#�����w��>�f��#.���㼰�R�@��:X�x<�t�<>=nt(=\�)= =�b�<���:8�uՆ���H�'�<�`�:K��M����1���Ǿ�   �    �����_���վ>E�����{�i�+�'��*׽z�Z��z����<�P^=m�=�Z�=� �=~[�=cm�=�N�=HL�=��=��]=��=�¡<�:M;C@��ļ���n6��()��&��m�(����ͼh���@���`k;8�<<�_�<�+�<���<8��<\Þ<��T;���j���ѽ�� ���`��$������X�Ѿ�6�K/���   �   X��D��	;�9���#ܾ?����ıL��X����������<-V=�
�=f��=�F�=���=p��=���=J.�=���=���=DJ�=��S=�j=�`�<�q_<�;@�m����ȫT�Pks�Xv�X�]��,���û �_�p��;�H<$k�<�ϒ<�\i<�w;�xz��\6�7P�������M�뤋�ڲ�Üپɩ��j]�����   �    �.���+�C�!�����X��~ о�����8n�����V���C�hb<�\K=h�=h��=��=t�=Z��=��=�K�=�w�=���=�=��=�r�=܎U=|�(=8��<�m�<`�^<p��; ,7:��s�Љջp^���Qջ��t� �9�?�;�?�;���;��;�~#��"�r�������c,��u�?ꣾ�Ͼ�n��\��!�=+��   �   >@��<���1��� ���
����� ��������2��^н�.'�8
<��@=��=���=8��=���=*� >^>p0�=H�=� �=�!�=���=ߎ�=[��=��t=$WI=��=���<��<�A.<�)Q;�-�`Ի�l�PA�ඥ��m� T� ����R��穼~5�BZ�����EE��!�� ��#��X��c �gd1��c<��   �   �cK��qG���;��)�w9�ɚ�h���Z��m�?�ھ⽸�?��@�;�R9=1��=H��=2��=��=�O>"�>+�>|�=��=���=a��=��=Nb�=�q�=J
t=^�F=d�=\i�< փ<�,�; S��ϻ�	�0$������׻ ��� /ٻ��X���&,V�7�������6U� ���bþb���ʧ��*���;��bG��   �   �U������g����{��(\��X8�db���߾���*,O�tV�x�+��S<�&]=\�=p�=�l�=4A�=3� >a�=0��=a�=X>�=���=\�=���=2	�=x��=��e=�zM=&�8=�\'=�2= K=:�=z�=��=�t=�= ��< �z<0����U��ģ�P@d�x����侢���F9�K�\�[,|�I���Ï���   �   ������������w��0X�U�4���</۾�����JJ�$���"�hzi<4�_=���=X_�=��=,��=��=:��=�<�=د�=���=���=~�=�і=4ׅ=�-m=tkR=�};=Γ(=H�=�N=~$	=�5=�=N�="�=��=���<�A�<������国s`�a�^�rƢ�}�߾��X�5���X�B�w���������   �   J��?������πj�y�L��+��y�^ξ�	��n/<��̽������<�Ag=%�=���=��=��=n��=��="�=@`�=5�=���=al�=|�p=�KM=�/=��=�?=���<X�<�4�<�{�<���<���<P�=�2=�=��<<L�<��Q;\"μ%-��w���*9N����kҾ|�	�:�+�z�L��Zj�怿�q���   �   @G~�ٟy�W�k��#V�P�:�;������w��j���*`&�zî�T ü��<��q=L�=�7�=R�=$��=��=�#�=X�=�=� �=pi=�6==d��<�܆<x3<<��<�<q<pH<���<B�<(��<�� =66=67=�}=��<ؕ=<Pi�B�W��Eٽ�4�^��\ȼ�=�������D:���U�&Wk� Xy��   �   ��_�h�[�h�O��?<�R�#�C�$�׾�o���9`�"��1��P�C����<��|=���=ފ�=B��=���=�S�=��="/�=�sm=
�)=��<��<������x��﷼�ռ��ּ�������s ��)T���<D�<���<�J=�J"=�[$=R�=���< V¹p��"���@0�md�!ġ�� ׾�y�:�"��Q;���N��`[��   �   �y=��:��/��
��	
���侟D������V6���ٽV�?��iU:hP=�=�ݦ=�&�=���=��=p��=,�=H==���<@�W;C��2��$�d�\/��{q��x��_���_���`�r�&�T�̼@]� �;�l�<p�=�^(=nZ8=d,0=:�	=��y<(�`��*`�U�޽�4�HY��k;�����b����f.��{9��   �   Q�����n�G� ���޾i����Џ��DR�����$����ۼ0 X<D�2=v,�=՟=p�=��=SÓ=B�i=��=�)@<�u���:����Ίν;*��c��{��p����&����Qֽ1է�rOl�Z 	�`�+��'<�<�'=�H=��O=p9="� =��<9ּ�P������G���&h����پ������@A��   �   ���)�S�ܾERǾb竾o����Z�A��Pǽ.�H���	�(��<�E=+�=r�=�=a��=j�T=�7�<��:;�$���R��Y�ؽzH��6�]S�`g��p�s�m�T`���I��,�8
��̽�4��~	��I���=�<�= vP=Bj=��e=�Z@=4��<�~;��G���
��/H�L����Ǥ�����c�ؾJ'��   �   0̮��D��r���c���^{��cL����	�׽R��\hʼ  �;��=��O=�(}=ׅ=lFz=:�G=��< .���h�T~���;�*�5�+6h�F[��	����Ϯ��H��ru���f���c{�BhL� ��m�׽8���rʼ�;�=v�O=*}=F؅=Jz=@�G= �< ǃ�x]�?w��T7��5�:0h��ꊾ~W��J����   �   t�o�N�m�VN`���I�T,��
�>�̽0��*���(��XB�<ȸ=�uP=�j=ʰe=�V@=x�<@;�������
�w4H�,����ʤ�d���k�ؾ+�% ��-�.�ܾ�UǾg꫾�����Z�D�RUǽr�H� �	�ė�<L�E=x�=X�=��=���=@�T=G�<�#;;���@K����ؽnC�H�6�WS�
g��   �   �v��k�f�������JֽTϧ�<Fl�r�� �+�x!'< �<�'=� H=̣O=m9=ғ = �<�Hּ�U����*�G����:k��[�پ���"��}C����!�
q�"� ���޾  ���ҏ��GR�m�� (����ۼ��W< �2=�,�=�՟=Jq�=��=�œ=��i=��=hR@<P]��~{:��y����νk ���]��   �   �i��sp��R����X��>�`���&���̼(I�P/�;�p�<4�=�^(=2Y8=8*0=�	=P�y<��`�^2`�m�޽8�4�a[��>��Ղᾛd������.��}9��{=��:��/���E
�����F��đ��KY6�?�ٽ�?���T: O=��=ަ=�'�=���=��=��={�=t
== ��< �X;)�����ނd�q'���   �   �ط���ռ�ּ��������Y � �R���<��<���<K=J"=�Z$=4�=���< \Ĺ� ������2�pd�ơ�U׾M{���"��S;���N��b[���_�l�[�L�O��A<���#�TD�(�׾mq��4<`���+4��8�C����<,�|=ࢪ=���=\��=D��=�U�=�=D2�=2{m=��)=X�<�<P����ix��   �   ��<XR<<��< <�<pH<��<pF�<���<v� =6=t6=�|=@��<X�=<�]i��W��Hٽ��4�c_��ʼ�S�����hF:�E�U��Xk��Yy��H~���y���k�%V���:�D������$y��`����a&�MŮ��ü<�<0�q=p�=8�=�R�=<��=,�=�%�=��=���=��=pi=<"6==Ȟ�<�   �   �"/=b�=�C=H��<�
�<�9�<(�<���<$��<r�=�2=>�=��<tI�<��Q;\'μ�.�������:N�����ҾC�	�(�+���L��[j��怿�r�����ن�����΁j�V�L��+�Zz��^ξZ
��X0<�H�̽������<�Ag=<�=���=l��=ė�=`��=<��=�#�=�a�=2�=�=�n�=��p=QM=�   �   �/m=~mR=�;=R�(=r�=�O=%	=R6=2�=6�=�=|�=���<@@�< �$���曽a�J�^�Ǣ�>�߾H���5�0�X��w���������������k�w�A1X���4�Z���/۾��KJ���ང�"��yi<2�_=���=�_�=,��=���=\��=���=@=�=���=���=���=��=�Җ=^؅=�   �   B��=|�e=jzM=��8=f\'=:2=�J=޳=.�=l�=�t=�=��<(�z<���6�(V����~@d�1x����侷��G9�a�\�m,|�O���ŏ���U������_�����{��(\��X8�Ib�V�߾����+O�V�Ȗ+� �S<']=%\�=��=�l�=:A�=2� >a�=&��=a�=P>�=���=:�=���=	�=�   �   P0m=�mR=8�;=�(=R�=�P=>&	=�7=��=��=x�=&�=��<D�<���n���䛽`�ښ^�Ƣ��߾����5�*�X���w�G��f���h���j��]��I�w�?0X���4����v.۾	����IJ���ོ�"���i<��_=��=�_�=b��=���=x��=���=P=�=���=���=���=��=�Җ=~؅=�   �   |#/=H�=E=$��<��<�=�<���<Ⱥ�<L��<:�=�5=Z�=���<�P�<�R;�μ�+�������7N�/��lҾ܅	�x�+���L��Yj��倿Mq���������^���j�j�L��+��x��\ξ����-<���̽������<,Dg=&�=���=܀�=��=���=`��=�#�=b�=I�=��=�n�=��p=�QM=�   �   ��<PW<<8�<�<��< *H<��<`M�<���<V� =(:=�:=R�=���<x�=<�@i�ڵW��Bٽ,�4��\���Ƽ�n�������C:�=�U��Uk�HVy�|E~��y���k�"V��:��������v������]&�!�����¼�$�<��q=�	�=�8�=XS�=���=n�=�%�=��=���=�=�i=�"6=�=,��<�   �   dַ�бռ|�ּ���P���L ��R��
<`�<8 �<�O=RO"=0`$=j�=��< 	��������.�Djd�`¡���־�x���"��O;���N��^[���_�Q�[�e�O��=<���#��A���׾�m���6`����-��P�C�t��<��|=j��=���=��=���=4V�=R�=q2�=v{m=��)=��<P
<Д��Pfx��   �    i���o��\����W��J�`��&���̼�7�@U�;�z�<��=@d(=b_8=10=��	=��y<أ`�*#`���޽�4�\W��9���|� a�Η�L}.�Uy9�Bw=�|:��/����
�����A������CS6�'�ٽ��?��%W:
V=e�=�ߦ=�(�=���=�=e��=��=�
==���<��X;h(��r��D�d�
'���   �   lv�@k�������Iֽ�ͧ�<Bl����o+�6'< �<�'=BH=ܪO=*u9=�� =@�<�)ּ�K��z��G����=e��d�پ}�����?������l�=� ��޾:����͏�(@R�Z�����L�ۼ�X<H�2=/�=wן=zr�=Q�=KƓ=f�i=N�=�S@<�\��>{:��y���ν$ ���]��   �   7�o���m��M`� �I��,��
�V�̽�-������ �� M�<n�=�{P=�j≠e=X`@=���<`�;���R��.
�+H�����XĤ����a�ؾ
#辌�p%�-�ܾiNǾ�㫾g���cZ��<��IǽށH�h�	���<@�E=��=�=��=N��=:�T=TH�<�*;;���K��z�ؽ`C�5�6��VS��	g��   �   ̮��D���q��tc���]{�cL��#�׽;��X_ʼ�F�;��=N�O=N/}=�څ=tOz=b�G=�.�< �~�pR�mp��'3��5�k*h��犾�S��{���HȮ� A��Mn��7`��GX{�P^L�ރ��׽����Rʼ�f�;��=��O=�.}=�م=Lz=��G=�!�< ���]�"w��H7���5�20h��ꊾtW��<����   �   �)�1�ܾRǾ"竾"����Z�5@�OǽD�H���	�H��<�E=�=��=�=\��=ԪT=W�<��;;�����C����ؽo>���6��PS��g���o���m��G`���I��	,��
�݅̽�(��<��0ٟ��R�<��=�{P=,j=D�e=�\@=|��<��;���#���
��/H�H����Ǥ�����[�ؾ>'��   �   M�����n�6� ���޾/���@Џ��CR�7���"����ۼ�X<��2=�.�=�ן=�s�=�=�ȓ=��i=>�=({@<�D��m:��q��cxνJ���X�0q� f�������kAֽ-ǧ��7l�&��(Y+��D'< $�<*'=�H=�O=Fr9=�� =P�<�7ּtP������G���$h����پ������>A��   �   �y=��:��/��
��	
����hD��Џ��9V6�s�ٽ��?��1V:�S=	�=�ߦ=�)�=��=�=�=��=�==���<@ZY;������rd�����`���g��Р���P��\�`�,�&���̼��pv�;��<��=4d(=B^8=/0=��	=0�y<h�`�4*`�3�޽ݷ4�DY��j;�����b����f.��{9��   �   ��_�g�[�d�O��?<�H�#�C���׾�o��x9`����0����C����<��|=z��= ��=��=3��=,X�=��=�5�=�m=��)=�+�<H6<�6��@5x�����ęռЛּ����t(/ ���P��<$�<\�<~P=�N"=�^$=R�=T��< ����������70��ld� ġ�� ׾�y�;�"��Q;���N��`[��   �   BG~�ڟy�W�k��#V�J�:�3�������w��D����_&��®���¼� �<��q=�	�=H9�=T�=���=��=�'�=��=vĨ=6�=�&i=~*6==���<D �<�y<<�< 2<ب<0?H<\��<,S�<ج�<F� =8:=$:=�=���<��=<�Mi��W�nEٽ�4�
^��\ȼ�=�������D:���U�(Wk�Xy��   �   K��?������̀j�w�L��+��y��]ξ�	��9/<���̽h����<>Cg=�=���=B��=���=���=���=$%�=�c�=\�=_��={q�=l�p=LWM=D)/=��=^J=���<`�<\D�<��<���<���<��=�5=²=���<N�<��Q;�!μ	-��h���&9N����kҾ|�	�;�+�|�L��Zj�怿�q���   �   ������������w��0X�S�4���3/۾�����JJ��ཊ�"��|i<��_=ꘫ=�_�=���= ��=���=v��=>�=���=���=���=��=IԖ=�م=P3m=�pR=�;=��(=��=�R=�'	=�8=D�=��=p�=��=ԫ�<�B�<������国n`�`�^�rƢ�|�߾��X�5���X�B�w���������   �   �̿�rȿ�轿%p��4���ހ���P�t� �q�꾐��.E�Q�Ƚ�+ּ��<g��=��=H��=8��=�Q�=T��=u�=��=r��=���=0�=>��=.�u=�/`=ƜQ=�I=��G=�RK=��R=�g]=��h=N�r=R�w=Lyr=�a\=�S-=,V�<�q���e�����VX��\���w��"��R�d��aԘ�C����콿cmȿ�   �   ٞȿ�ſ����J����啿�8}�(�L�>���K澵���2b@�l½��ż��<P��=2�=P��=�y�=Z��=��=*^�=q>�=���=za�=��=�w=FNZ=��D=��6=�0=v�0=R<7=:�A=h�O=.X^=xrk=�s=�Np=��\=X�/=xZ�<`2��0�Z�-���R�"���{�뾖���1N�9 ~�"%��ۓ������iſ�   �   ����$C��gg��D�H��p���A��&���ؾ����?x2���������k�<s��=��=���=��=\��=��=���=Ld�=���=X�|=��N=��&=��=��<���<�2�<l��<�'�<.�=�X%=*�==�T=H>d=(5i=ֲ\=|�6=(��<@m�ʪ:���۽2'C�阾ZGݾë���B���p��W���ݡ�B���'���   �   ��嫿LϢ����YS��%|[���0��z���þ�\����������p�={�=��=\��=4��=�=�<�=��=$$�=�E=n�=@�<P�; ���{�ȴ"�hn	���s� bc;�K<,��<,�=ֺ*=�YI=�d[=D�Z=�Z@=`W=@��; ���#��Ȗ*��*��0Ǿ�c�_(1��p[�:"��n;������-����   �   �����D���&��\��uf��4A�F ��I�xl����_����R�\�@o�:��(=҇�=�+�=���=z2�=�K�=^��=��S= �=�w:<h��<p伈�1���_���x���{�z�i���D�br�`��� ~��h�<<d=�<~�=D=�&T=�NI=x=8b�<41��8D��p���e�i骾0�쾱����@��(e�*ڂ�絏�F���   �   B<�����u�l�_��_C��r#�*q�Tž����J�4�fLƽ�
��NU<��>=�,�=�o�=��=�K�=�w=��'=�ӊ<��$���������Ȼ�Z"�^��������*r����߽�涽�z��(�*��!���o�;�2�<��=*�E=6�N=�4=���< ^K��a1���нz66�(C����þ&S�""�l�A��>^���t�>����   �   ��X�"U�OXI�H�6��,�����Ҿo-��2�Z���;����k����<�P=Z��=
�=[�=�]=��= Q�;�������ҽ #�d)3��O�V�b�Yk���g���Y�)�B�X$��(�n��ld�(7¼ X�;��<3,=�M=�J=�=�ɉ<�����������T�$����ξl�!��5���G�YUT��   �   �1*��>'������������+;���#m�q �����<�� ;��="%\= �=f�z=F]M=���< 
94x�����~v�bv;��bo�����z��?��������Z��L��������N�>���ս�v��O��8W<:�=�DB=��X=`G=�	=��;8e �����*�Ka�/���#PǾ��V��SH��j&��   �   cl��� ���뾙�Ծ����֔����h�
'�Dֽ�\�@�F�l��<,�,=�'_=�h=
�F=�8�< �z:lJ�b������hSX��鎾�ﰾ2�Ͼ��8<���q���%�������Ծh���������h�!'�Jֽt�\���F����<��,=4(_=�h=�G=�D�<��|:?����0���MX�:掾�밾��Ͼ��7���   �   䆳������V������H����N��
� �ս�|v��A���i<��=rEB=��X=�G=l�	= ��;|n �󴨽4.�VPa�m���	TǾh�����K��m&�f4*��A'�A���������j/;�
��[(m�� �z���̪����; �=�$\=� �=��z=bbM=��< �9zk������q��p;�.\o�D�����v���   �   Mk��g�o�Y�T|B�E�#�J$�g��Xad�('¼���;��<�4,=�M=tJ=�=��<���������\�T�񟙾ξ,n�|#�45�cH�YXT���X�U�[I���6�/�����Ҿ�/��ȉZ����?����k���<v�P=ԭ�=_�=v!�=�]=��=`��;g����X�ҽ��6#3�F}O�`�b��   �   o��|��<h����߽�޶��s����*�x�����;�:�<:�=6�E=��N=Z�4=@��<��L�i1�r�н�96�]E��t�þ�T�8"���A��A^���t������=��g���V�u��_��aC��t#��r�eVž|����4��OƽP�PDU<��>=-�=|p�=���=DN�= w=j�'=��<�$����E�������������   �   ��x�N�{�،i�<�D��f�ܞ���>����<<@F�<n�=�D=N'T=�MI=�	=�[�<�:���G��Vr���e�~몾ڗ�T��t�@��*e�fۂ�9������'���F��((��1]��wf��6A����K�n���_�X����\���:��(=臋=~,�=¼�=R4�=FN�=���=��S=غ= �:<h��|S��1���_��   �   �N�h�"��E	��s���c; �K<�<P�=ν*=|[I=�e[=b�Z=�Y@=�U=���;���&��ʘ*�+,���Ǿ�d��)1��r[�,#��x<�����S�����%櫿WТ�����-T���}[���0��{�I�þ�]��b������@����=�=��=9��=���=��=@?�=��=�'�=�E=�=���<�q�; !��   �   ��<h��<@?�<���<�1�<R�=\%=��==<T=X?d=�5i=��\=��6=p��<����:���۽�(C�꘾�Hݾ�����B�0�p�zX��gޡ��B���(��t����C��#h���󡿱H��p���A�Q'���ؾL���"y2�����<���j�<y��=��=r��=��=���=���=���=�f�=@��=2�|=�N=ο&=�=�   �   ��D=�7=ޓ0= �0=�>7=�A=ҥO=DY^=$sk=:s=Op=��\=��/=�X�<�<���Z�h.��R�è��K����62N�� ~��%��G�������ſH�ȿ)ſ�������敿d9}���L����L�󟜾�b@�ul½@�żX�<Z��=f�=���=\z�=���=��=_�=�?�=���=�b�=#�=�w=�QZ=�   �   �/`=t�Q=��I=��G=VRK=<�R=:g]=��h=�r=�w=$yr=�a\=rS-=�U�<`s�F�e�X���MVX��\��"x���"��R�d��oԘ�M����콿fmȿ�̿�rȿ�轿p��&����݀���P�T� �9��b���-E���Ƚp*ּ!�<���=.��=^��=D��=�Q�=Z��= u�=��=h��=���=�/�=(��=��u=�   �   6�D=,7=<�0=x�0=
?7=��A=��O=Z^=tk=8s=8Pp=Ҝ\=^�/=\\�<*��
�Z�Z,�Z�R�Ч����M��91N��~��$������2����ſi�ȿNſE������a啿?8}���L�����J����4a@��j½(�ż��<���=��=��=�z�=��=��=$_�=�?�=̬�=�b�=/�=w=�QZ=�   �   ��<���<�@�<t��<�3�<��=�]%=<�==T=NAd=�7i=.�\=��6=`��<`I��:��۽&C�T蘾YFݾ���B��p�/W���ܡ�AA���&��͛��PB���f����mG���p���A��%�D�ؾ�����v2�(���l
��dq�<���=��=���=��=���=ҿ�=���=�f�=N��=L�|=�N=��&=�=�   �   �L���"�B	���r�@�c;�K<��<��=>�*=0^I=�h[=��Z=�]@=~Z=P��; ��o!��"�*��)���
Ǿ�b�,'1��o[�b!��x:���������㫿3΢����jR��~z[�%�0�xy��þ}[�����̰���}�B�=��=�=���=
��=5�=p?�=��=�'�=,�E=�=���<�s�;���   �   �x�~�{�֋i�ھD�e�ܚ��0,��P�<<L�<��=DD=r+T=�RI=�=�j�<,'��A���m��e��窾ߒ�>����@�&e�ق������ ��g���MC���%���Z��<f��2A����G�Zj��z�_�;��Љ\��'�:j�(=߉�=�-�=���=�4�=�N�=ڥ�=��S=�=Х:<��0S���1�P�_��   �   F��H���g���߽�ݶ��r���*�����;�A�<2�=��E=$�N=��4=���<��I��Z1��нz36�/A���þ�Q�6"�,�A�U<^��t�ǜ���:��t큿��u���_�@]C��p#�fo�#Qžk����|4�Gƽ���hU<��>=3/�=�q�=���=�N�=�w=ޑ'=��<��$�x��.���辻�������   �   -k���g�+�Y��{B���#��#��e��z^d�� ¼0��;�%�<\9,=JM=!J=f�=�Չ<����V��������T�����Vξ(j���� 5���G�_RT���X�U�kUI���6�k*���Ҿ�*����Z�| �s6��`�k����<ܣP=
��=��=d"�=]=r�= ��;hf��E�ҽ��0#3�:}O�J�b��   �   ֆ�������V����������N�X
���ս�yv��:��y<0�=�JB=�X=�G=�	=�;�[ �����B&�0Fa�!���uLǾ�������E��g&��.*��;'������'����';���em�	 ��𺽀����;��=6+\=�"�=t�z=2dM=d��< z9k������q�|p;�*\o�B����zv���   �   [l��� �����y�Ծ|��������h�p'��Bֽޝ\�X�F�|��<��,=�-_=6h=�G=�R�< �~:4� ������ HX��⎾�簾P�Ͼ�2��-g��m������Ծ����@�����h�'�<ֽ,�\���F�؜�< �,=�-_=�h=�G=�G�<��|:�>�؟��$���MX�:掾�밾��Ͼ��7���   �   �1*��>'������������+;���]#m�� �\���:��pބ;8�=l*\=p#�=8�z=�hM=���< �94_������l��j;��Uo�����顾*r��r���V����R������2��X�N���M�ս�nv��*����<f�=�KB=��X=�	G=(�	=0��;^d �r���*�Ka�-���$PǾ��X��TH��j&��   �   ��X� U�MXI�?�6��,���bҾ<-����Z����:����k���<��P==��=��=J$�=�]= =���;(M�-�����ҽ+�3��vO�J�b�
�j���g���Y��uB�n�#�*�M^���Rd��¼pԆ;X.�<�;,=�M=" J=ތ=p͉<������������T�!����ξl�!��5���G�ZUT��   �   C<�����u�h�_��_C��r#�q��Sž�����4�gKƽX�PZU<H�>=*/�=�r�=��=Q�=w=�'=���<x�$�����燽`���|�j��������X]��{�߽�ն��k��4~*�H�����;�K�<4�=*�E=4�N=��4=L��<  K�a1�A�нh66�$C����þ'S�$"�m�A��>^���t�@����   �   �����D���&��\��sf��4A�> ��I�Wl��l�_�U����\����:��(=���=A.�=���=�6�=�P�=�=��S=��=��:<HL�h6�D�1� �_���x�B�{�^|i���D��X�x����哻�<<tV�<&�=fD=<,T=rRI==�e�< /���C���o���e�f骾1�쾲����@��(e�,ڂ�鵏�I���   �   ��	嫿MϢ����YS��!|[���0��z���þ�\�����R��������=��=F�=���=:��=��=�A�=��=&+�=D�E=�=`�<`��;�b����X"�h	��^r���d;0�K<x�<f�=��*=�`I=0j[=*�Z=B]@=:Y= ��;D���#����*��*��/Ǿ�c�_(1��p[�<"��o;������/����   �   ����%C��hg��E�H��p���A��&���ؾ����x2�#������Xn�<S��=��=\��=��=ֱ�=H��=���=�h�==@�|=��N=�&=D	=�,�<P��<�N�<h��<d?�<x�=�a%=p�==^T=�Bd=�8i=Z�\=8�6=���<�`�X�:���۽*'C�阾ZGݾī���B���p��W���ݡ�B���'���   �   ۞ȿ�ſ����J����啿�8}�(�L�<���K澬���b@��k½x�ż��<���=��=��=�z�=���=L�=`�=�@�=��=^d�=��=�w=hUZ=��D=�7=֗0=�1=B7=JB=��O=�[^=Puk=s=�Pp=�\=,�/=�[�< /����Z�-���R�"���{�뾗���1N�9 ~�"%��ۓ������kſ�   �   �~�(�z���
��Fɿ����΋� yZ��B"��㾑쒾�U(�l���]��V`0=���=N��=��=��=��=���=��=�=���=dxq=�O=�
6=�%&=b =�n$=J21=��D=�<]=Pow=1'�=ʑ=���=�p�=�5�=̝:=l:�<�޼.���x�8�NᙾT����$�g�\�����ի��ɿt��j���t%��   �   �D��� ������߿��ſ�;��ag����V��:��޾ո��c�#��ލ� CC���2=�#�=C�=��=?�=-�=��=���= ��=�A}=0dR=H9.=^>=�=h��<ʭ==�*=rF=r2d=�y�=��=��=�=�~=L�;=���<�ͼ\(���3��i��U,��!��X�B��qި�D+ƿ~�ǡ��2� ��   �   #���m`��G��|տE$���㟿3f���;K��j�TiѾ�l��~f�D�{� u�:h9=�g�=mp�=���=t8�=z�=�H�=�f�=r`=,H'=�X�<\��<�!< l�;P�;P��;�Z<�P�<�M�<@)=`�Q=BNt=�c�=m�=n�x=bR?=<Э< ��"����%��[��XF־�h��L�o����@��MA�� տ��迨8���   �   �����|9ֿ�Ŀ$���Ò�V�n��p9�A������{�o������I��'<J0B=#��=��=���=>ȫ=���=rq=~9*=ǻ< ��;؆H���Լ���¡%���$��y�l�ռ�_��{w:<��<�F =I6=��^=&�s=8'm=�B=��<hQ&�*���� ��iy������	�]:��@o����� ���S�ÿ��տT��   �   >̿|�ȿ׍�� O��
���G끿A�R���"�q/���K��ֽ:��G�<FsJ=��=n��=��=G�=/D=��<@�;�¼�oI�ԯ���ɹ���ӽ��߽d�ܽ�U˽H���D����3�����
�:Ը�<$N=��I=�X=AC=Hc�< �n:�)=�Z��4�Q�	C��q���"��LR����� 󘿤����񽿷yȿ�   �   �g���}��P���j��MH��Mb]��2�"		�~�ƾޅ�}�!��Ȟ�O�����<�O=��=�w�=6�d=�=��[<LI����R��A��ێ���\���8��CJ�D�Q�zON���@�**�����׽T8������s�p��<�=�69=��===HtQ<�/ּE����\%�����{Xƾ&q�1�1��[�vm������tԢ�����   �   N��������xZv�߽W�-5�m�Y�ܾH�����O�^���L�������=�%M=�+c=Z�H=^=o�;)���-���c��Ң.���`�`����Ř�p���1|��K���fy����vn�Z�>��3� ��n�H���V�0�u<"=p�.=�C#=t��<���T�U�0��4pM�;Л���پ�X��3�Q�U��Ut�2S��"4���   �   �Df��]b�V���B�f�)�e�����]�P�l�����ǝ�H�ü�>d<VH=NB=�16=�t�<�Q	;r��<����t�}BT�Ǚ��GW����̾���R���
������={�0�Ѿ�o��:~����b�\v!��̽��L�p+(���<F=�K*=�m=��[<��������S��N/e������9ܾ���H'�`v@�(wT�za��   �   ʈ.�c�+���!����j���*�Ҿ�D��Jbs�}$������k(���?��j�<x%'=܃,=���<�V�;����*��͎�j�g�D��?�̾|���l�L ���*�&�.���+���!�˽�b���a�ҾH���gs��$������s(� <A��e�<Z%'=��,=���< ��;y��#����T�g�U@����̾<	���i��H �E�*��   �   P��:����u�_�ѾOk���z����b��q!��̽��L�@(��<�=vK*=�j=��[<�ƴ�t���T���4e�b���4>ܾ{��K'��y@��zT��}a��Hf��ab�� V���B�+�)����r��d���l�Ԟ�̝�ļ82d<�G=�B=�56=���< �	;.��'���qo�<T�򕌾�R����̾,�侦����   �   �w����u��&���n��~>��.�����H��cV�ؠu<4=^�.=rB#=��<`:���U�f��{tM�ӛ�O�پ[��3�i�U�PYt�
U��6��=������|!���]v���W��5�s���ܾ�����O�H��L��	����=�&M=�.c=Z�H=�&=�;x���%���Y����.�M}`�U���D���ط���   �   �Q�vHN�$�@�$*�w���w׽�0�����P����<�
=�89=�==~=fQ<T;ּ�����_%�䅆�\[ƾ�r�v�1���[� o��\���F֢�o��}i���������k���I���d]��2��
	��ƾ�߅���!��˞��V�����< O=��=�y�=�d=�=��[<�.����R�8�������V��8��<J��   �   �߽�ܽ4L˽d���q���t3��� !�:�Ŵ<�R=��I=V�X=�@C=�_�<  n:�/=����0�Q�E���sﾎ�"��NR�0���l���5�����u{ȿ�?̿0�ȿp����P��T���a쁿�R�p�"��1�M��K��ֽ�
��D�<>sJ=O��=ᷜ=O��=\�=27D=d��< H;��¼0_I���������,�ӽ�   �   �%���$��l���ռh�^���y:��<�L =�M6=��^=��s=�'m=��B=	�<X^&�������fly�������	��^:��Bo���5�����ÿ��տʀ�_��2���:ֿĿ/����Ò���n��q9�%������J�o�����I�h"<0B=���=��=V��=xʫ=���=Zyq=TB*=�ۻ<@��;�RH���Լ���   �   P��;�5�;���;P'Z<T^�<|Y�<�D)=�Q=Qt=�d�=�m�=��x=�Q?=\ͭ<%�����%��\���G־�i�.�L����^A��1B��տ��迹9��1���ra��9��Qտ %��`䟿�f���<K�9k�2jѾ"m��Cg��{��X�:�g9=Qh�= q�=���=�9�=^�=�J�=�i�=�`=�O'=i�< ��<��!<�   �   h�=���<��=�=�*=F=�4d=�z�=��=�=C�=�~=��;=���<h�ͼ�)����3�2j��*-�o�!�ȨX��B���ި��+ƿ�W���|� �4E��� �i���]�߿4�ſ"<���g���V��:�m�޾�����#��ލ�`FC���2=�#�=��=^�=�?�=�=;��=��=���=�E}=hR=�=.=�B=�   �   �%&=�a =2n$=21=��D=h<]=�nw='�=�ɑ=���=tp�=�5�=v�:=�9�<�޼������8�{ᙾ����$���\�����)ի���ɿ���t���v%��~� (�m������3ɿ����΋��xZ�cB"�M�_쒾qU(��k��pX���`0=֢�=f��=4��=���=��=���=��=�=���=Lxq=�O=Z
6=�   �   ��=��<�=�=J*=~F=5d=�z�=h��=h�=��=*�~=8�;=P��<8�ͼ�'����3�Ni���+価�!���X��A��$ި��*ƿ�K����� ��D�X� �a���l�߿^�ſh;���f���V�:�B�޾6���x�#�Iݍ��"C�2�2=n$�=��=��=�?�=5�=@��=$��=���=�E}= hR=�=.=�B=�   �    ��;�7�;���;@)Z<�_�<[�<�E)=*�Q=FRt=Ze�=on�=��x=�T?=�ԭ<D�������%�<[��gE־!h�7�L������?���@��Cտ��迡7�����^_��A�迅տe#���⟿�e���:K��i��gѾ�k���d���{���:�j9=Ci�=�q�=��=$:�=��=K�=�i�=`=�O'=i�<��<��!<�   �   Ԓ%�0�$��k�H�ռ��^��z: �<N =BO6=�^=l�s=�*m=>�B=,�<�B&�摃�l���gy�|�����	��[:�2?o�������ÿ0�տ�}�s��S��8ֿ�Ŀ����������n�,o9�������o������I�0:<4B=���=��=潴=�ʫ=ñ�=�yq=vB*=�ۻ<���;�RH�X�Լ���   �   ��߽ܘܽ�K˽���򆆽< 3���X�:�ɴ<$U=��I=�Y=lEC=�k�<�p:$=���轪�Q�OA���n�S�"��JR�Ј����,���@�xȿD<̿��ȿ-����M������ꁿ(�R�F�"��,���K�d�սL ��R�<xJ=��=鸜=�=��=�7D=��< J;��¼._I��������� �ӽ�   �   �Q�^HN� �@��#*�0��Fw׽/0��8���G�(��<�=�<9=��=== �Q<l"ּ
����Y%�ҁ���Uƾ�o�$1���[�l������Ң�����e��|��}���Rh���F���_]���2�L	���ƾ�ۅ�(�!��Þ��?��x��<x"O=���=�z�=��d=ԯ=x�[<.��x�R��7�������V��8��<J��   �   �w������u����Wn�:~>�e.������H� YV���u<$=x�.=8I#=X��<�Խ���U�_��PlM��͛�T�پ�V�h
3�d�U��Rt�gQ��>2��]��-������Wv�ºW�x	5�'���ܾ`����O��｀�L�������=4,M=H2c=��H=$(=pƜ;x��\%���Y����.�M}`�X���D���ط���   �   L��2����u�H�Ѿ0k��~z��d�b�Rq!��̽&�L�8(���<�=R*=�s=�[<����������h*e�Ω��6ܾ��F'�:s@��sT�bva�1Af�=Zb��V�=�B�p�)�ԓ�K���쨾�zl�D��
��� �ü0_d<RO=�B=�86=P��<��	;f��󌮽eo�<T�򕌾�R����̾.�侨����   �   ̈.�a�+���!���P����ҾrD���as��|$������h(��?��s�<�+'="�,=p��<PҰ;�n���������g��<��n�̾6���f��E ���*�l�.��+�Z�!���������Ҿ�@�� \s�	x$�ݴ���_(� �=��z�<x,'=Ȋ,=���<���;�w�Y#�����M�g�U@����̾B	���i��H �H�*��   �   �Df��]b�|V���B�]�)�Y��x��4��l���bƝ�h�ü�Nd<�M=�B=�;6=��< v
;(��o����j�6T�F����N����̾�������������xp�I�Ѿ�f���v��$�b�Xl!�"̽��L���'����<`=FR*=�q=�[<0���$���2��B/e������9ܾ���H'�cv@�*wT�za��   �   P��������tZv�ٽW�$5�b�:�ܾ"���&�O�o�N�L��,��t�=0,M=f4c=��H=�.=`�;����[���O����.�Nv`�`���𼘾B����r������p����0n�x>�T)����r�H��4V���u<�=�.=�H#=|��<�����U����pM�8Л���پ�X��3�T�U��Ut�4S��$4���   �   �g���}��P���j��KH��Hb]��2�		�a�ƾ�݅��!��Ǟ��I��\��<�!O=t�=�|�=ʩd=N�=(�[<���ƳR��.���x��lP�4�8�n5J�ʝQ�<AN�1�@��*�����m׽F(������ �d��<�=n?9=��==T=�Q< ,ּĤ��n\%�����yXƾ&q�3�1��[�xm������uԢ�����   �   >̿�ȿٍ�� O��	���F끿<�R���"�]/���K�Aֽ4��M�<BwJ=M�=��=�=���=H?D=P��<�	;`�¼�NI�T���������ӽ<�߽I�ܽ�A˽�����~����2�ר� ��:�ش<nZ=,�I=�Y=�EC=�i�<�ko:�(=����Q�C��q���"��LR�򉁿󘿥����񽿺yȿ�   �   �����~9ֿ�Ŀ$���Ò�Q�n��p9�9��z���G�o����8�I�0<&3B=#��=��=D��=�̫=���=��q=�J*=��<�T�;�H�H}Լ"��΃%�h�$��]�@fռ �^���|:��<�T =�T6=��^=ܯs=2,m=p�B=<�<`K&������ ��iy������	�]:��@o��������U�ÿ��տW��   �   $���p`��I��|տE$���㟿2f���;K��j�GiѾxl��Rf�P�{�@��:�i9=Di�=*r�=���=q;�=F�=EM�=xl�=�`=W'=�y�< ʏ<��!<P�;`��;� �;�JZ<�n�<�g�<:K)=��Q=�Ut=�f�=<o�=��x=�T?=Pӭ<0�������%��[��WF־�h��L�o����@��NA��!տ��迪8���   �   �D��� ������߿��ſ�;��`g����V��:��޾θ��J�#�aލ��9C�|�2=\$�= �=��=�@�=�=X��=~��=S��=,I}=2lR=�A.=`G=:=d��<f�==*=�F=�7d=|�=M��=�=*�=��~=N�;=씓<D�ͼ<(���3��i��T,��!��X�B��pި�D+ƿ~�ȡ��2� ��   �   :)��&&��Q�H��%O��Y0ٿ����s	���CT�(0��sɾ�t�kA��:�!����<�l=��=��=���=�`�=��=��=���=BT=4A'=�k=���<H��<�۶<���<�� =��!=�G=v_o=�ډ=���=�<�=�=��=��$=��A;�{\��e�w��VFϾH�$W�!t������Gڿ�����j`�(%&��   �   xM&�FP#�`����4����տ�¯����UwP�aT��Zž� o�T��@��Z�<*l=$��=���=�=�
�=�	�=�"�=Zg=�1=�=�z�<H�u<Ѐ><h�A<�~<0��<�t�<j*=��V=z�=�ʏ=槗=�v�=�|=|%=��;��R��i���z�(�ʾR�z'S�틿𰿄�ֿ������v���F#��   �   F���*��v��aHn˿�&��闃�iE���Pu��/�^��F����۴<X�h=�]�=<��=���=t��=U�=N=B�
=Q�< f;;���x!������d\���y��;˻`��;�<�%=�B=bp=*��=�f�=�3r=f&=��;H�6�W���zzi��Q��9P���G�t���������˿|��� �����   �   ����i��2����ۿ�P�������q��4�^���⦾��E�f/��h���4s�<��a=yG�=��=�Ì=~f=�N=�2�<�{����޼�A�Vu��ɫ��U��'ɝ����0�d������@� ;xױ<ȩ=��Q=j�i=��^=U%=�F<D���\Խ�eN�M���K� �S�5��,r��陿cV��?Jۿˢ�����x��   �   �%����pZ��Hݿ��ÿ����$���T����� ݾ�X���%�r"��8�J��G�<��S=$�x=�"m=��9=�#�< B��h~��Ā��R��[�����~#��\)�&�g��j�Tpֽ暽8':�T`����<�`�<"]/=?=��=4��<Q��7��tO,���޾ǐ�$�T�����p����¿Wܿlz�B����   �   t�޿�ۿ�пϤ��yL���Ԏ��Xh� \4����������i��>��X�������<<�;= ?@=�=H�a<(�����`�}�ǽ���z�>��
g�����q��ۣ����I�����o� LI�6
���j��̐�� ؖ9p��<�d=P�=��<�	�@gn��E�J]l��H������3�D5g�i����0���t��Ͽukڿ�   �   =���G�����WJ���R���lk��P>����lվK���;3�o���t5���&<���<�=p��<0��;��ܼ`!��2��^�<���|�N���3���;оC߾߰�ʣ�PӾV��Wʢ�[��~�H����(:��X��c�H��<���<p;�<�Ŏ;Ժ�<���>63��W����Ӿ�I��<�u+i����� �����t����   �   �R��B鑿LP���b|�0:]���9�)���\���`�W�wm���Cl��7�,�<��<��<���;Lg�\~��.2���X��o��\��K		�XA�6"�r�%�\#�����L�j8�Ǿ͇����c�r%��{��ε� ���<t1�<Ьz< �<�r�g��.��X|S�#���y߾���WH7���Z�4�y�GO��O[���   �   -fc���_���S�hS@���'�W��&�ݾty����h�Bk���߼p��;���<�4�<�^<8��,y��)����`������ؾ�	��%�=�=�R�Q��^�^jc�Ɲ_��S��V@�!�'�����ݾ�|����h�o�<���<#߼�t�;̿�<|9�<t<�&���r�������`���U�ؾ�	�� %���=�X�Q��^��   �   ��%��#�i���I�3�Ǿ����zc�� �)u��֬��\�����<�0�<��z<�=�N�g�6��\�S�~���d}߾?���K7�X�Z�E�y�vQ���]���T���둿nR���f|��=]�z�9�����Q¢���W�ls���Kl��.7���<���<���<`�;�Q��v��$-�.�X�땾�j�����%	��=��2"��   �   ����ྟJӾY����Ţ����e�H�����2������b���<��<�9�<0��;�������:3�wZ��i�ӾL���<��.i�u
����H���Ѱ��g?��J��,
��^L���T���ok�?S>����oվ����>3������>��p<H��<4�=X��<@�;ğܼ'���'��ԉ<��x|��������v5оr߾�   �   L���I��������o�ZEI�n���⽎b���y�� ��9���<h=�=�	�<��	�bnn��H�<al�SK�����8�3�8g����s2���v��O	Ͽ�mڿϓ޿�ۿ�пʦ��;N��%֎�[h�^4�s��8�����i��@��X�@e�����<��;=�C@=�=��a<,���.�`�N�ǽ���h�>��g�E����l���   �   8V)��&�5��Td�Rfֽ~ݚ�:��I����<Tm�<*a/=*?=�=�}�<`Y�����R,���K�޾}��N�T�������z�¿Yܿ�|�m���'����j\�JݿN�ÿ���:%���T�����ݾkZ����%��$����J�dG�<.�S=��x=(m=�9=P7�<@����_��	���qH���������#��   �   �K�����s���z�d�0�����`;;@�<ί=T�Q=�i=,�^=�T%=(F<���_ԽhN�񵪾j� �́5��.r��ꙿ�W���Kۿq������y���Ҭ��i�+4��A�ۿ�Q��t���rq��4����㦾~�E�D1�����xr�<��a=�H�={�=Yƌ=�f=�W=�H�<���x�޼d�@��l�������   �   �����E��8�y���ʻ���;�<�+=ԲB=�ep=~��=lg�=:4r=�&=���;P�6�����@|i�8S��Q�ߔG�'���}���}�˿7}�|�����p�����+������HI�ro˿1'��h����iE��v��.�^�,H�L���۴<�h=�^�=���=h��=���=,�=�#N=\�
=�c�< 	<;�T��
���   �   ��><�B<�%~<dǵ< }�<�m*=��V=��=�ˏ=r��=�v�=$�|=�%=0	�;��R��j���z���ʾ��&(S�t틿���ֿT���F��԰�G#��M&��P#����Z�/5���տï�8����wP��T�=[ž� o����\@��Z�<�l=���=H��=���=��=F�=Y$�=Rg=l�1=~=l��<8�u<�   �   ���<@۶<`��<�� =h�!=��G="_o=�ډ=���=�<�=�
�=��=4�$=@�A;�|\�f�9w���FϾn�;$W�9t������Gڿ����p`�*%&�:)��&&��Q�<��O��?0ٿu���[	��kCT�0�ysɾ��t��@��j�!����<r�l=��=>��=���=�`�=*��=��=���=VT=*A'=�k=h��<�   �   �><�B<0&~<�ǵ<l}�<�m*=�V= �=�ˏ=¨�=]w�=4�|=h%= �;��R��i�6�z���ʾ�&'S��싿�ﰿ&�ֿA������(��hF#�M&��O#����~�%4���տ^¯������vP��S�,Zžno�����=��^�<�l=���=���=ʙ�=��=I�=`$�=Xg=j�1=z=`��< �u<�   �   �����E����y���ʻ��;ࢠ<P,=��B=�fp=��=*h�=>6r=�
&=p�;��6�����Fyi�Q���O���G�𓄿������˿-{�V��d������.*�x�ܯ�MGm˿�%��;����gE���t��V�^�KD���t�<X�h=L_�=���=���=⨞=F�=$N=d�
=�c�<�<;�T��
���   �   �K�����U����d���������H;P�<�=��Q=<�i=�^=�X%=8)F< ��ZԽ�cN����k� �&5�l+r��虿BU���HۿK�����w����:h�1���ۿ�O��s���+q�4�#��"ᦾ��E��+������@|�<޳a=�I�= ��=�ƌ=f=�W=�H�<�����޼z�@��l�������   �   8V)�~&�(��:d�fֽݚ� :�dG����<,q�<�c/=�?=��=���<hF�����1M,�s푾��޾V��G�T��������¿GUܿnx�$����$����_X��Fݿ��ÿ)����"���T����>�ܾW��@�%�G���J�S�< �S=�x=�)m=��9=L8�<�����_�����}H���������#��   �   K���F������Նo�0EI�:�
���a���v�� 	�9 ��<�k=@�=4�<|	��_n�XC��Yl�8F��Z����3��2g����.���r���Ͽ*iڿ�޿Nۿ�
п�����J���Ҏ��Uh��Y4���6���l�i��;��X�@3�����<��;=hF@=�=x�a<,�����`�B�ǽ���n�>��g�I����l���   �   ����྘JӾL����Ţ����"�H�j��2���� ~b�P�<h��<<H�<@��;��������23�[U����Ӿ�G�O�<�W(i����������������:��RE�����5H���P��cik��M>����iվ����73�C���p"���F<X��<~�=���<��;�ܼ���y'��щ<��x|�Ć�����{5оv߾�   �   ��%��#�h���I��2�lǾ샛�Hzc�� �,t��@���괺���<$?�<�z<0�<��g��'���wS��u߾��ZE7�8�Z�N�y�'M��Y��FP���摿N��~^|��6]�K�9�x
��򻢾%�W��e���7l���6�x&�<��<���< ��;�N�bv��
-�"�X�땾�j�����)	��=��2"��   �   0fc���_���S�dS@��'�L���ݾTy��1�h��j��흽\߼д�;�ͺ<�G�<��<��kl�����B�`�d��ؾ7	���$��=�y�Q�ɘ^��ac���_���S��O@���'�r��P�ݾ�u��\�h��f��睽H�޼���;Ѻ<E�<��<"��r�������`���X�ؾ�	�� %���=�^�Q��^��   �   �R��C鑿LP���b|�*:]�y�9� ���;����W�yl��Al��7��!�<��<X��<`*�;;�to��b(��X�6畾Cf��Y��	��:�/"�5�%�:#�����F�L-�Ǿ����sc����l��������$��<�@�<�z<0�<�x�g�>.��6|S����y߾���ZH7���Z�:�y�IO��Q[���   �   =���G�����UJ���R���lk��P>�߉��lվ(��>;3�J����.��8:<���<Μ=��<`T�;�ܼ<�������<�Rq|�\������0о��޾��(��EӾ'���N��������H�6���)�������a���<���<@H�<��;.��x���	63��W����Ӿ�I��<�x+i����� �����v����   �   y�޿�ۿ�пФ��yL���Ԏ��Xh�\4����ݵ��8�i�>�$X�@������<@<=:J@=�=��a<�g��N�`���ǽʳ���>���f�
���h�������돾�����~o�>I�&���}��Y��t]�� ��9�<�o=��=4�<��	�,en��E�&]l��H������3�H5g�j����0���t��Ͽwkڿ�   �   �%����rZ��Hݿ��ÿ����$���T����� ݾ�X����%�p!��0�J��P�<��S=��x=B.m=��9=�J�<�/��`B��A���J>��=t��p��D
#�vO)��	&�Ȣ�X^��[ֽԚ� 	:��.���<(�<zh/=h?=��=��<�K��s��AO,����޾Ȑ�&�T�����q����¿Wܿnz�E����   �   ����i��2����ۿ�P�������q��4�N���⦾��E��.�� ����y�<�a=�J�=���=*Ɍ=�f=4`=|]�<������޼b�@��c��p���\B��ȶ��w�����d����Lܘ���;���<ܷ=��Q=��i=��^=JY%=&F<r��@\Խ�eN�E���J� �T�5��,r��陿eV��@JۿϢ�����x��   �   H���*� �v��bHn˿�&��藃�iE���Bu���^��F�����ߴ<H�h=�_�=���==��=���=��=�*N=:�
=�u�<�<;�(�p��l��D.���]y� �ʻ�M�;$��<03=2�B=,kp=���=Ni�=�7r="&=P�;$�6����dzi��Q��8P���G�u���������˿|��������   �   vM&�FP#�`����4����տ�¯����UwP�`T��Zž� o���v?��\�<�l= ��=�=���=��=��=�%�=
g=��1=d= ��<��u<ح><�+B<8<~<�ѵ<���<�q*=b�V= �=͏=���=�w�=��|=�%=��;�R��i���z�'�ʾS�{'S�틿𰿄�ֿ������x���F#��   �   �#R�@�M��-B��0��z�B���ۿ'���d��[!?�#������5��㛽��ƻv/$=�r�=���=ʩ�=n*�=ޖ=T�{=��C=h�=Dױ<��?<�f�;@��:@K<;`��;�-�<��<� =D,R=_D�=�x�=��=
�=�i=4N�<
��E����r?�"#�����0B�7�����ܿ8x��:�0��HB���M��   �   �/N��*J�ʶ>���-������˕׿tF������;�}�������281������٤��g#=�È=H��=�`�=�f�=[y�=�|]=D�=�I�<��,< /�� ���$3�й�������;L�<���<$44=�*h=���=���=�K�=�vd=Xl�<�cs���3�:�y{��<��ۈ>�b����묿t,ٿ=��e�(�-��>�dJ��   �   6�B�.[?� �4�|�$�f��Z����QͿ�ࢿ��v���1�t��Q���dX$�W�����c =Af�=���=�!�=���=�&I=�� =�H<��ۻ��¼,���(?���N�f�G�.*��{�H�g��Ma;ؘ�<<�=�U=*�x=�^|=� V==�<�c9�	Ù�q�,��晾�o����3��gy�����hο���R����$� �4�@2?��   �   �?2��!/���%�J��h5�y忊%��J���B�a��!�9پ\����z�B�c����:T=��b=�ht=�{Y=�J=D/�<�L ��:x�C���ҽ�-�7r������۽~9��RN��޽0������;���<f�.=K=4�;=7�<�̻9�����}����ܾrd#�N�c��T�������Z��\�6w%��.��   �   � ��h�؈��B�*��޷̿kS������RG��r��� �d�h｠�-����;�I
=�#5=��&=̄�< �:(H��	@��Hս�����2��MN��b`��ig�t�b���R��=9�)z����9���:�"������<dT=N|=�K�<��B���F�����+�i�+^��}n���G�����*&���̿k�������P��   �   ���0���|�������ο�W���h��g2b�y�(�}$��z��*�8�ܸ���PN<�>�<��<P�n<h�A��yH�V���8���AM�2ҁ�.F��׭�ܯ��-���%��#[����������lV�"9�ڹԽ�+m�(n���B�;�D�<|E�<pۀ;��ȧ����;�/���ȶ�s(��a�>���E���[Ϳ]��;���s��   �   ���
x߿�oԿ#�¿�(��A���-n��!9�@������T�s����!��h��(,<��<`5�; ���L)w�{���:7�����׹��7�;������j��2h��(����}mҾ�����\C@�����[���Tfռ���: M< `�;<!��@L��C����s����$��e�7��4l��됿W���>0���ӿ��޿�   �   w۶�n�����l��M���O�h��<������Ҿ�����2���������X����<�F;���(�~������H��ؑ��ľ׽�������-��E@��EL��P�H9M��	B�10�R�����vɾ�#��4�O���؉��˼ N7� ��;�"˻����<����0�����\pо��%�9���e�{#���⚿w���=M���   �   �k��#���ჿa�p�9�R���0�����#׾`����&K�����Ti���� V#;@	D;ĺ��_���TBF�v���d+Ӿ�&��
.�6�O��m�MԂ�����[n���%��䃿��p��R�*�0�B��A(׾�����+K�U��.]i�\���H#; 2D;����_�8���<F�׎���&Ӿ�#�w.�8�O���m��т�#����   �   ��P��4M��B�V-0��N�����fqɾ ����O����҉�H�˼ 4�0��;�>˻����B��V�0����rtоY�`�9���e��%��.嚿����O��6޶� ��v�>o��d����h��<�3��M�Ҿd�����2�n������pf��0�<�gF;Ԑ��8�~�������H��ԑ�*�ľ��������-��A@�1AL��   �   ����d�)%�n ��hҾ��������d=@��{��Ţ��@Tռ�0�:�(M<@X�;�)��QP��}��X�s�&��U��0�7�8l��퐿�����2���ӿt�޿g���z߿GrԿ��¿�*���B���0n�;$9�(��u���A�s�<��$�����,<,�< m�;ܝ��fw����p47����������;�𾋬�T���   �   ���������U��弝������eV�L3���Խ~m��Y���z�;�L�<�G�< ΀;��������;�������Hu(���a�𿏿G���]Ϳ������,u�> ����m��\���ο�Y��j���4b�Y�(�B'��|����8�߸����`N<D�<���<h�n<x�A�@jH�^���
��T:M��́�XA���ѭ�W����   �   \ag�f�b�!�R��69�t�c�潊x��Z�"��
�蘃<xY=
=`L�< fC�Z�F�Ź��Z�i�v`��p���G������'��~ ̿���0��.���	��Nj����C���}�̿�T��ʛ��G�t����V�d��j�f�-����;�K
=�'5=�&=x��<���:,*���6��OսU����2��EN��Z`��   �   �f���z�m۽�/���E��8�0�|뎼�\�;���<��.=�K=�;=�6�<p�̻R;��Ľ�����ܾ�e#��c��U��u������@��]�Vx%�@�.��@2��"/���%�4��26�Uz忡&��*�����a��!��پN���
|���c����:�=Z�b=Pmt=�Y=.S=�D�< �����w�j��q�ҽ�"��   �   ��N���G�*�)��c�Џg���a;��<T�=��U=v�x=�`|=�V=0<�<hk9��ę���,��百Cq����3��hy�\���iοD��� ��R�$�ަ4�*3?� �B�
\?���4�&�$����E����RͿ\ᢿ��v���1�e��𖕾"Y$�������c =3g�=2��=�#�=���=P-I=,� =ЭH<0sۻ��¼���?��   �   0
3����獻���;P �< ��<�74=�-h=���=[��=L�=�vd=8k�<(is���!�:�(|�������>�ʮ��o쬿	-ٿf=�Df���-�b�>��J� 0N�P+J�.�>��-�*��&�� �׿�F�����.�;�֍��ٜ��n81�����Pؤ��h#=wĈ=��=�a�='h�={�=Ā]=��=�T�<-< ������   �    ��:�H<;П�;d-�<���<n =�+R=7D�=�x�=뙘=���=hi=(M�<t��ɛ���r?�]#����>0B�S����*�ܿHx� �F�0��HB���M��#R�:�M��-B���0��z�2���ۿ�&���d��,!?����H����5�㛽��ƻ�/$=�r�=���=婰=�*�=1ޖ=t�{=��C=��=Lױ<��?<pf�;�   �   H
3� ���獻0��;� �<|��<�74=�-h=���=���=nL�=xd=hn�<�_s��֫:�7{��
����>�/����묿,ٿ�<��e���-�~�>��J�"/N�Z*J�R�>�R�-�������:�׿�E��>��K�;�����򛟾671���� Ǥ��i#=�Ĉ=S��=�a�=Ah�={�=Ԁ]=�=�T�< -< �������   �   ��N���G�"�)��c��g���a;訰<��=f�U=��x=`b|=�V=DB�<�Y9�����n�,�晾�n����3��fy����hο#��������$�8�4�d1?�N�B�HZ?�H�4���$����7����PͿ�ߢ���v���1����5����V$��	�����~f =h�=���=N$�=Ә�=~-I=4� =ȭH<psۻD�¼���$?��   �   �f���z�e۽�/���E��ʮ0�<ꎼ�b�;���<>�.=�K=ʵ;=4?�<�^̻�6��`���|��o�ܾcc#��c��S������Ć忌��[�&v%���.��>2�` /���%�J���4�}w�=$��6�����a���!�8پ�����x��~c� * ;>=��b=�nt=��Y=�S=�D�<� �����w�z����ҽ�"��   �   hag�l�b� �R��69��s�)��3x����"�`�
�@��<�[=x�=PV�<��A�Z�F�����x�i�F\��0m���G�y����$���̿������� �H���g����hA����̿�Q��l���EG�3q������d�$c��-�p!�;2P
=�*5=��&=���< ��:�)���6��Xս`����2��EN��Z`��   �   ���������U��޼�������eV�3��Խ6m��U��`��;DT�<�R�<��;���H�����;������(q(�p�a�����5C���YͿ��翟��^r�b�����z��|�鿸�ο�U���f���/b�G�(�&!�fx����8��ָ��鼈l<�M�< ��< �n<H�A��iH�>�����^:M��́�bA���ѭ�_����   �   ����d�)%�g ��hҾu���炅�)=@�{��ߡ�� Oռ ��:(?M<��;���zG��!��V�s�����0����7��1l��鐿1����-��Cӿت޿���5u߿�lԿ��¿f&��?��E*n��9���P���_�s�������~��8,<4 �<���;���Rw�H��b47����������;�𾐬�Z���   �   ��P��4M��B�R-0��N�����Pqɾ ��T�O�Q�Nщ��˼ �.�p�;��ʻ$���6����0������lоQ�$�9��e�g!��j�����J���ض�����J쪿rj�����r�h�V<�-����Ҿ����L�2������������<`�F;܊��x�~����߃H��ԑ�-�ľ���������-��A@�6AL��   �   �k��!#���ჿ_�p�4�R���0�����#׾@����&K���ｌQi������#;��D;�����^����7F�|���b"Ӿ&!�2.�m�O�[�m��ς�����Qi��� ��X߃��p�0�R�`�0����3׾����N!K�%�ｘGi�h�����#;��D;d���� _�v�轾<F�ώ���&Ӿ�#�}.�?�O���m��т�&����   �   {۶�o�����l��K���J�h��<������Ҿ������2�I���f��&��(< �F;|��ڎ~���:~H�<ё���ľQ���G���-��=@��<L�W�P��0M�}B�v)0�EK�����`lɾ��@�O����ʉ���˼ 2*�`'�;p�ʻ����;����0�����Vpо��'�9���e�#���⚿{���@M���   �   ���
x߿�oԿ#�¿�(��A���-n��!9�5��������s���\�� ���6,<|%�<@��;<����w���_.7�ӹ��y���J�;��9��Ҙ�5��a��!���nbҾ�����~���6@� q������l:ռ�{�:XLM<@��;h���J�����g�s����#��h�7��4l��됿Z���B0���ӿ��޿�   �   ���0���|�������ο�W���h��b2b�q�(�g$�z����8��ڸ���鼘g<Q�<���<��n<`A�0[H�ղ��%��83M��Ɂ��<���̭�᤺����� ����P����������1^V��,�!�Խ�m��>��0��;L^�<lW�<��;������4�;�������s(��a�@���	E���[Ϳa��?���s��   �   � � i�ڈ��B�*��޷̿iS������LG��r������d�g�f�-���;�P
=�-5=�&=Ĩ�<��:���
.����Խ5����2�D>N��R`�$Yg�H�b�V�R�n/9��m����n����"���
����<�a="�=\Y�< �A���F�������i�^��}n���G�����-&���̿o�������T��   �   �?2��!/���%�J��j5�y忉%��I���=�a��!�&پ>����z���c�@ ;x=��b=�rt=v�Y=b[=�X�< ��������w�����ҽ�콙[��wo��ڽ�%���<��`�0�HЎ����;\��<n�.=�
K=\�;=A�<e̻
8������}���ܾrd#�O�c��T�����"��Z��\�8w%��.��   �   8�B�0[?� �4�|�$�h��[����QͿ�ࢿ��v��1�f��?���&X$����@��Jf =�h�=ߋ�=&�=P��=�3I=� =(�H<Pۻ�¼�w�:?���N��rG���)��J��ag� �b;p��<��=��U=��x=6e|=XV=�C�<h[9�[�@�,��晾�o����3��gy�����hο���T����$��4�B2?��   �   �/N��*J�ʶ>���-������ʕ׿qF������;�v�������81�8����Ф��i#=ň=Բ�=�b�=di�=�|�=��]=r�=�^�<X,-< ܳ� �����2����в���;�+�<4��<<4=j1h=?��=���=5M�=yd=po�<�_s�U��:�u{��;��܈>�b����묿s,ٿ=��e�(�-��>�fJ��   �   cC����z��k��S���8����@|�ܟο�>����f�P��X�˾h"m��N��i��(��<ea=�*�=�\�=ޒ=�;|=x�C=�=���<`�<;�s��b���������3���m��|E<���<V�*=��a=�!�=��=g�=KF=p�<���e���t�rZо�!��j��(���п���~ ���9��gT��>k���z��   �   >/{�6�u��yf��P�b�5�~k�����I˿̖��رb����ʺǾ\�g�V/���6�<�i[=t��=��=X��=^�_=j� =�9�< ��; %�����D�����	�<5���̼xd� �9�Ǉ<��=�(E=Ht=7N�=D�}=¯@=���<0�����[Po��̾�l���e��]��cAͿ�k ��M�$q6��[P�2�f���u��   �   t*l�VUg��zY���D���,�p����3���Kד�(�V��3�zɻ��rX���ν`AԼ,h�<b�H=v�v=�Os=��J=�h=��U<`������b.M��w������ʣ�]���O����]�����o��W�;���<�/=|pX=Zb\=�/=$��<����8۽�4_�����?c��VY�
@��^ÿ7��F����,���D�0<Y��g��   �   HV�*R�H/F�FZ4���������5������'+D�B���6����@�����pH��X^�<�	'=�:=�X=��<�{q�<@�t�������� ������Z �U�%�"����� �Auʽ卽�)���&�Eh<�y= �!=�5=��m<�M׼�뾽NlF�5?��6P���E�Y�����i�࿊������3���E�D�Q��   �   �)<��8�#/��  ����U/��ǿ�p��}�o�$X,����pϑ�>#�"����)��8��<�_�<�<�<��;�m���o��ͽ^Y���@���h�p���뎾�ᒾ�ꏾ~P���n���F����`۽F���J� �9��<�]�<�9<𛥼����'�)����뾍X-��p�$�����ǿ�x����M��V.��l8��   �   � �Hl��y�d
�����-ѿ;!�������L�sR��9¾�do����x�c���<���<��#<��Ȼȏ�꺤��5	��KG��T���T��>��ؾ�羴��-B�-Qھ�'ľ�᧾2���N�� �w���.� �7���;pj�;�Mx���p�^����q��<þ���& L�+g��`����Ͽ���	�~������   �   ����6��.���Q̿�C�������u_��x&�f�ZG����9��Ľ�$��7!� �
���n�28:��O��.� �e�n��:���<ѾW'��1��4#�Υ-�%�1�3p.�4�$���7�(�վ�B����u���&��ʽ��L�(]��Pҭ�L�Ɓ,�,�ǽ9�:��L��8��z�%�^�F���B���rʿR����������   �   S�ؿ5cտD�ʿ���U���}���b��0�Z��{˳��g���%���޼��?����\�=���½*(�2k��(U���`���ud7��xR���g�7�u�]{���v��i���T�}�9�v�z���1���r���,��CʽXwI��S���X����H����v���e��Z��"~ �Q.��u`���ҏ��{F��jɿŎԿ�   �   d���V���~���7���H}�̑U�T(,�-�`���ځ�s�!�ӣ���(��;��xn��l�#��䮽���̬�<����3�c�)�A�R�E2z�C����_��UU��Q���4���9������M}���U��+,���C����܁�\�!�ʨ���(�>���h��J�#��ޮ�v��s������41���)�2�R��-z������\��pR���   �   >{���v�G�i�k�T���9� |��������Ko��<�,�=ʽoI�L���X���异���.z�f�<^���� �$T.�cy`���_���LI��%mɿ�Կ��ؿUfտ<�ʿ���UX�������b��0�����γ���g����(��<�޼(�?��u��N�=��½�$(��g��~P���Z���p`7�\tR���g�(�u��   �   �1�	l.�A�$�
��3���վC>��y�u�J�&�(ʽ�L�8P��0��� L���,��ǽ �:�SO�����%�L^�B��������tʿE��'���,��`����9����]T̿�E������x_�${&�mi꾯I����9���Ľ�$�85!���
��ln��+:�=G��Z� �ڲn��5��7Ѿ� ��_-��0#���-��   �   �쾰;�Kھ;"ľ�ܧ��	���N�N��n��ĥ.��7��(�; v�;�Tx��p�ھ���q��?þ���L��h���a����ϿK��	�������� ��m��{��	
����0/ѿ�"�� ���L�T��;¾�go�����c���<���<@$<бȻ:��ӱ���/	�\DG��P��jO�������׾I ��   �   �ܒ�1揾�K��L n�t�F�T���U۽�=���1� ��9�#�<Dd�< 9<l���Ϡ����'����{�jZ-�V�p�����ȭǿ�z�����N�.X.�nn8�`+<���8��$/�P" �җ�81�J�ǿ�q��x�o��Y,�����Б��?#�γ���*��D��<�h�<@K�<�h�;�R����o�R�ͽ�R�<�@���h��k��&玾�   �   ��%��"����E �8kʽp܍�^��d&��gh<0�=�!=�7=@�m<�R׼�xnF��@��dQ�B�E�c���`�����x�������3��E�άQ��V��R��0F�j[4����l��@� 6��h���Y,D����7���@�����I��a�<�'=*�:=�_=%�<�p�,1�~���0���0�����T ��   �   ����P���vG��v�]�����}o� ��;,��<|�/=ttX=�d\=�/=8��<����:۽�6_����)d��WY��@��WÿB8�������,���D�N=Y�� g��+l�zVg��{Y���D�B�,���z������ד���V��4�8ʻ��sX�z�ν(BԼ�i�<~�H=�v=�Ts=��J=Xp=@�U<8�������M��o��vx���   �   ��	��-�|�̼�c� �9�ч<��=H,E=�	t=O�=D�}=�@=X��<���[��vQo�[̾!m���e�r^���AͿ.l �dN��q6��\P�ֆf�<�u��/{���u�>zf�P���5��k�r���<J˿���(�b�����Ǿ��g��/ཐ�8�<�j[=[��=(�=ﰇ=N�_= � =�D�<P˩;X%�Ќ�������   �   (��ر��X3� �m��{E<`��< �*=��a=�!�=��=�f�=�JF= �<��Tf��t�t��Zо�!��j��(��=�п���� ���9��gT��>k� �z�cC����z��k��S���8����.|���ο�>����f�&���˾"m�JN潀h��L��<�ea=�*�=]�=.ޒ=�;|=��C=�= ��< �<;`s��b���   �   ��	��-���̼��c� �9 ҇<�=�,E=&
t=VO�=�}=(�@=Ь�<&��W���Oo�?̾Vl���e��]��AͿ�k ��M��p6��[P���f��u��.{���u�yf�P���5�k�h���bI˿U����b�����Ǿ4�g��-ཐ�P;�<�k[=���=]�=���=d�_=*� =�D�< ˩;�%� ��������   �   ����Z���~G��|�]�|���|o����;��<$�/=xuX=Nf\=�/=���<Ļ�7۽�3_�璿��b��UY�}?���ÿ.6�����&�,���D�&;Y��g�>)l�$Tg��yY���D�Ķ,��
�{��B����֓���V�3�,Ȼ��pX�֜ν�8Լp�<l�H=�v=bUs=Z�J=�p=0�U<X��$���$ M��o���x���   �   ��%��"����B �"kʽM܍���8b&��kh<��=0�!=�:=��m<�D׼;龽�jF��=��PO�j�E��������࿾����n�3�P�E�ƩQ��V��R��-F�Y4�������z��3�������)D���5��J�@�����<���i�<�'=��:=�`=&�<@�p�1�����C���M�����T ��   �   �ܒ�9揾 L��M n�i�F�B���U۽�=���/� y�9�(�<�k�<19<ȏ������ӕ'�������W-��p�؜��[�ǿ�v���4L�U.�k8��'<�l�8�~!/�� �v��7-���ǿo���o�NV,���v͑�4;#����� �����<o�<$O�<pq�;�Q��V�o�Q�ͽ�R�J�@���h��k��4玾�   �   �쾷;�Kھ9"ľ�ܧ��	����N�� n��
�.���7�PH�;P��;�0x�h�p�ȹ�I�q�@:þD����K��e��D^��k�Ͽ3��8
	���>��^� ��j�Vx��
�����*ѿG�����PL�{P��6¾O`o�����xc�`|<���< $<��Ȼ�������/	�[DG��P��sO�������׾U ��   �   �1�l.�C�$�	��3���վ2>��H�u��&�Mʽj}L�HH������X�K��x,���ǽ��:�	J�����/�%�^�v�������oʿ������ޑ��\��3��9��1O̿=A�������r_�Nv&�.b�tD��~�9��yĽ^�#��!� Z
��^n��):��F��6� �̲n��5��	7Ѿ� ��e-��0#���-��   �   D{���v�I�i�k�T���9�|��������*o����,��;ʽTkI��@���oX�`��Ѐ��)s�(�e�XW���{ �<N.�r`�����k����C��0gɿ��Կ%�ؿ`տ:�ʿ@��VS��z{��E�b��
0����ǳ���g���U����޼H�?��j�� �=��½l$(��g��{P���Z���u`7�dtR���g�/�u��   �   h���X������8���H}�ʑU�M(,�#�F����ف��!����L(��+��\V��̪#�1خ���~������.���)�`�R�1)z�2���!Z���O��z���r�����������C}���U��$,�b����ց�t�!�=�����'��&��DY��`�#�Vݮ�
��;��춼�51���)�9�R��-z������\��sR���   �   U�ؿ7cտE�ʿ���U���}���b��0�N��V˳���g�J�d#����޼��?�Pb��z�=�c�½�(�4d��L��GU�����\7�pR���g�,�u�${���v�j�i���T���9��x�������k����,�\4ʽ�aI��5��(jX�X��-���v���e��Z�� ~ �Q.��u`���׏��F��#jɿɎԿ�   �   ����6��/���Q̿�C�������u_��x&��e�.G��*�9� ~Ľ��#��!� +
��Cn��:��>���} ���n�z1���1Ѿu���)��,#�}�-��|1��g.�>�$�R��0��~վt9����u�)�&���ɽHqL��8���l����K�6|,�s�ǽ��:�lL��.��{�%�
^�H���F���rʿW����������   �   � �Fl��y�d
�����-ѿ9!�������L�iR��9¾do����}c�@�<���<8&$<p]Ȼ�t����n*	�n=G�iL���J�������׾���~��(5��Dھsľ�ק������N�;�	e����.���7��w�;@��; 2x��p����v�q��<þ��( L�-g��
`����Ͽ���	��������   �   �)<��8�#/��  ����U/��ǿ}p��y�o�X,����Eϑ��=#�e��� ����<�u�<�[�<��; 8���o��ͽ�L��@�Z�h�g��m⎾�ג�i᏾eG����m���F�����J۽�4��p� ��97�<@t�<p89<L���X�����'�����뾎X-��p�&�����ǿ�x����M��V.��l8��   �   LV�,R�H/F�FZ4���������5������$+D�:���6��\�@�u����@���i�<�'=�:=hg=8�<��o��"�꤁�6����	��t���M ��%���!�y��k ��`ʽ=Ӎ����0&���h<ڈ=8�!=�==0�m<$F׼�꾽�kF�?��1P���E�[�����l�࿌������3���E�F�Q��   �   t*l�XUg��zY���D���,�p����1���Iד�%�V��3�iɻ��rX�Ξν�<Լ�o�<��H=��v=nYs=�J=�w=xV<c�����M�+h��hp������"|���?��؇]�T���No����;���<t0=(zX=�i\=�/=x��<<��8۽�4_�����>c��VY�@��_ÿ7��H����,���D�0<Y��g��   �   @/{�8�u��yf��P�b�5�~k�����I˿˖��ױb����úǾ>�g��.�p�P:�<Rl[=5��=L�=Q��=��_=v� =�N�<���;��$�L~��\�����	��%�L�̼��c� C�9T݇<��=�0E=Zt=�P�=��}=\�@=(��< �����DPo��̾�l���e��]��dAͿ�k ��M�$q6��[P�2�f���u��   �   �Ș��,��P���lx�|V�6[4�t��h쿝嵿/����9�˺�@I��bw���Y����;�21=6|=�V�= �}=��O=��=쪔< ��:�5j��Zټތ�<�X��L�H≼ <��p<�w=.�?=�m=:C�=6�k=�� = �B;�l����0j�� ���5@<��6���߷�Q��VT�6�5��tW�vy�R!��1���   �   p\��!��h��ws���R��M1�|����O沿;M��BT6���b8��i��V�S�P��;0�*=T�o=�,~="�d=8�/=�@�<���;PME���ԧ-��Q���_���U��^5�7��@y��jR;��<��=D�T=�n=6�_=8�=��<;H�e�z���<�����@�8��̈́�����U��<��
U2��SS���s�����ۑ��   �   ���e���.v�xve��]G�:�(���
�Y�ݿ*(��!y��m,�YD߾�`�����x1C� �;n�=�oI=LE=>K=��< �n�����W�6��_�����ҽ^�۽�սjͿ��Ᵹ�e��V�P���7u<��=�b5=r�9=�f=`�;Z�S��q����R�⾾t.���{�����Q0߿��@#)�~�G��ge�D.��{���   �   (&{�r�u���f���P���6�* �&	 ��I̿�a����c������ɾ~�m����BL+����;l��<��=�O�<@̛;(<����a�2��������-��'7��zG���M���H���9��!�z�������is�x,ܼ �(:|-�<L��<<�< �J:�%:�#���X�q�j�̾5v���e��N��!(ͿfX �
1�>H6��&P�bJf�ԇu��   �   rjZ��^V��JJ�
8��"�8`
�_��E��A���q�H��C	�P���K�&�˽��� b'9x]< I<(N9��I1��5��SU�M�:�ǆm��y��V����o��NЯ�I���.��ݖ��ar��@�/U�������B��ty��Ѣ;k&<�ED����#:ҽ��N�᰾;
���I�a���2���w�&�	��b!��"7�]I�b�U��   �   �9�F6���,�
�����)��_ſ�j����l��*�y3�`��DH&�ǵ��,k��0~���ۻ4ͼ��u��߽�g.�I-u��ޟ�XľW�H!����o.�]��5� �S���bǾ��(�z��3��2��������X���I'����Zq���(����~羪T*�իl���� �Ŀ���2�
������+� l5��   �   |_���L��������=�ǿ�5���J���B�3�	��g����d�-� �*��X�鼠^��:���ꍽ�����H�(���7þN���v��P,��u>��?J�S�N��K���?��.�Yh�*���|�ƾH��z�M���pd������x!�������ދe� i����	�(QA�ҝ��W��]'ƿ��翎�����2r��   �   ,������ �� տɉ��Y����-�� �L�
�3`վGE��Qx*�S���^kC�Hj��(��O����Z ��8Q��r���ھK[��3���U� #t��+�����9吿J���f���}v���W�Y5�x\��\ݾ����_	U�)6�<����!��| ���E����)�#���}Ծ����&K�Q���f������!ӿ�o濇��   �   �o��)m��
봿̳�����|Bw�0RH�.��i��y(���\H�U8���������~��f�5 F�y��,$���F�t����2������߾���r��cp������c���Fw��UH���ۚ⾸+��8aH�>������`�$�~�`�F�fu��J�����F�,|t�ބ��)/��o��������   �   U␿t�������xv��W�NU5�UY��Wݾ���U�b2�[7��$�!��| ��E�����)�����Ծz��J*K�t������뷺��$ӿXs��˰�����#��տ���������/��Q�L����cվ�G���{*������mC��f��ܼ�����zV �y2Q��n��Cھ�W�� 3��~U�t��(��� ���   �   ��N���J�<�?��.��d����_�ƾ<���S�M����Q^������촼�#�����v�,�e�Kl���	�TA���������)ƿ���<����� t�pa������H����鿫�ǿ�7��,L��TB��	�Ej���d�6� �������LU��@���㍽�����H�����2þչ��Ur��L,�dq>�$;J��   �   �*������ ����<]Ǿ��8�z���3�3)����輠���B'����nt��ފ(�!�����V*�®l����Y�ĿX���
�t����+�,n5��9�J	6���,����(��_+��aſMl��$�l�q*�6� ��\J&������k���c����ڻ��̼H�u���߽�`.��$u��ٟ�FRľ��,����   �   �ʯ��C��f)��$����Xr���?�UO�6�����B�PKy���;z&<@;D�
��G=ҽ��N�;㰾�<
���I����Y4���y�b�	�d!�:$7��^I�z�U��lZ��`V�rLJ��8��"�Na
�#�俱��_���"�H��D	�����K��˽h�� �)9h]<i<0 9�r:1��+��0O���:�9~m��t�����j���   �   ��M�C�H���9���!����ڜ���Ys�|ܼ�r+:�;�<Ч�<��< �J:h(:������q�K�̾�w�~�e��O���)ͿHY �2��I6�b(P�2Lf�ȉu�$({�V�u�l�f��P���6�!��	 ��J̿sb����c�����ɾ�m�]��M+�`��;���<j�=�_�<#�;� ����a�.���'�� 7�sG��   �   ��۽i�Խ�Ŀ��❽he��J�P���0Xu<�= g5=:�9=h=@�;��S��r����ɏ��u.��{�s���i1߿���$)���G�$ie��/�w|��Է��!���xw��we��^G�܋(�(�
�!�ݿ�(��"y�:n,�4E߾Ga��|���1C�`�;��=�sI=��E=$R=�ϛ<�n�dx��V���������ҽ�   �   ��_��U�|V5��/� &y� �R;L�<j�=�T=�
n=X�_=��= �<;
�e�F��>=������8�)΄�5�����꿢���U2�pTS�@�s����7ܑ��\���������ws�F�R��M1����9�迍沿hM���T6�f�쾌8�����<�S�@��;~�*=T�o=t/~=��d=��/=tK�<P)�;�0E����^�-�8�Q��   �   "<�r�M輨≼`@��p<:w=��?=��m=C�=��k=h� = �B;�l���jj��P���i@<��6���߷�x��lT�L�5��tW��y�Z!��1���Ș��,��G���lx�dV� [4�`��h�{嵿����9���I��w���Y���;j31=�|=�V�=F�}=��O=0�=\��< ��:`5j��Zټڌ��   �   Й_� �U��V5��/��%y�`�R;��<��=p�T=0n=�_=��= =;�e�&��d<��_����8��̈́�i������ ���T2�fSS���s�3��bۑ� \����� ��Xvs�H�R�M1���C���岿�L���S6�,�쾺7��v��p�S����;��*=�o=�/~=��d=��/=�K�<)�;(1E���|�-�Z�Q��   �   �۽|�Խ�Ŀ��❽\e�dJ�`����Yu<��=�g5=Ĭ9=pj=�);4�S��p���b��t.���{�򙫿�/߿d���")���G��fe��,��z��D��������t�Bue��\G�l�(��
�L�ݿO'���y��l,��B߾�_��h���,C��+�;� =uI=X�E=�R=Л<�n�hx�,�V���������ҽ�   �   �M�R�H���9���!��������<Ys�hܼ �+:�>�<��<��< L:� :�#���T�q���̾2u�E�e��M���&Ϳ�W �0�G6�`%P��Hf��u�*${�~�u���f��P�<�6��J �lH̿j`����c�R����ɾ�}m����E+����;p��<N�=b�<p'�;���n�a�G��� '�� 7�!sG��   �   �ʯ��C��n)��)����Xr���?�>O�㢶���B� Ey���;��&<`�C����>6ҽb�N�O߰��9
���I�<��11��v��	�Ba!�� 7�0[I�X�U�PhZ��\V��HJ�X8�"�_
�Z�俙 ��騊�]�H�)B	���֍K�=�˽��� F/9�&]<�q<P9��91��+��0O���:�M~m�u��*���j���   �   �*������ ����9]Ǿ���z�p�3��(�.񂽌�輠���('�����l��(�(�������R*�K�l�0��%�Ŀ[����
���Ċ+�j5��9�<6���,�R��>��i&￙]ſ�h����l�Y*�+0�����D&�R��� X�� 2�� �ڻ��̼��u�z�߽�`.��$u��ٟ�PRľ��<����   �   ��N���J�A�?��.��d����R�ƾ(����M�-���\��b~�`ߴ�\���������e�Df����	��NA�*���N���$ƿР������Np��]���v�������鿜�ǿc3���H���B���	�Ld����d��� �Y��Pt鼤H��^���⍽z�����H�����2þ޹��[r��L,�mq>�.;J��   �   Z␿w�������xv��W�KU5�PY��Wݾ��xU��1�V5����!�0s �b�E��輽��)�g����Ծ=���#K�X��� ��X���uӿ�l� 󿑩�����[�翑�Կ膼�Ў���+����L�D	��[վ*B���s*�@����_C��S��Ҷ������U �22Q��n��@ھ�W�� 3��~U�t� )��� ���   �   �o��-m��봿ͳ�����{Bw�,RH�'��Q��N(��1\H��6�C�����H�n�~��X�F�r�������;F��wt�`���_,��e���l���Rl���i���紿߰��7���=w�HNH���o�⾴$��WH��/�a�������~�o^齞F�Ku��B�����F�2|t�ℐ�./��s��������   �   1������ �� տɉ��W����-���L��`վE���w*�孼��cC�(S����� R ��,Q��j��Gھ�T�9�2��zU�%t�Q&��*���vߐ���������sv�~�W�MQ5��U�oRݾ|d�T�z-��/����!��q �$�E��켽4�)�����iԾ����&K�T���i������!ӿ�o濋��   �   ~_���L��������;�ǿ�5���J���B�'�	�kg�� �d�.� ����v�4B�����e܍������H����x-þ�����n��H,��l>�u6J���N�	�J���?�P.��`�c���ƾ����c�M�@��V���u�Pִ�L�������X�e��h����	�)QA�՝��[��`'ƿ��習�����4r��   �   �9�H6���,�
������(��_ſ�j����l��*�X3�$��|G&�A����[���"��@�ڻ �̼��u���߽�Z.�u�!՟��Lľu�>��Y��&���$� �S��YWǾ�袾��z���3�J�~邽���l�('�����n��P�(����g羨T*�ثl����$�Ŀ���4�
������+�"l5��   �   tjZ��^V��JJ�
8��"�8`
�^��D��?���k�H��C	�$����K�D�˽��� 096]<��<��8��+1�Q"��\I���:� vm�Lp������d��;ů�>��-$��P���Pr�N�?�I�𘶽0�B��y� ]�;x�&<`�C����B8ҽj�N��ా;
���I�b���2���w�(�	��b!��"7�
]I�d�U��   �   (&{�r�u���f���P���6�* �&	 ��I̿�a����c������ɾ�m�i��H+�@��;t��<�=�p�<�w�;���F�a�N䷽ۥ��� ��7��kG�c�M���H�l�9���!������� Hs�x�ۼ�c.:O�<d��<h%�< tL:�!:�������q�T�̾1v���e��N��$(ͿhX �
1�@H6��&P�fJf�҇u��   �   ���e���.v�zve��]G�8�(���
�[�ݿ*(��!y��m,�ID߾�`������.C��(�;<=�wI=�E=�X=|��<@|m�`� �V�����w��p�ҽ�w۽'�Խֻ���ڝ�� e�x=�@f��P}u<��=Pm5=��9=�l=`9;��S�Tq����E�⾼t.���{�����R0߿��B#)���G��ge�D.��{���   �   o\�� ��h��ws�ގR��M1�|����N沿;M��@T6���R8��6���S����;�*=:�o=�1~=��d=��/= U�<�V�;`E����(�-���Q�ؐ_�,�U��M5��'��y��,S;X �<�=�T=�n=$�_=�=`=;��e�E���<�����?�8��̈́�����V��<��U2��SS���s�����ۑ��   �   �E��-��X����-��"�q��I��
$�Ĵ���ɿ;ϔ�hBP�M��O꥾i72��d������Њ	=�[=��q=&*]=X@+=,,�<p��;��C�8��~�*�&�M��Z��]P�`�/�p����c�`g�;0»<��!=h�S=tfh=`�Q=4* =��	�d;��6�5�">��]W
�+VR�!.���V˿f���9%�KJ��~r� {��������   �   @���"���k���,����l��E�dV!�N� ��Kƿ�D��2L�U)�>����M.�2����ƻTq=�M=dq]=��A=�u=�q<`���Hy׼�6��r��S���x�������0w�8�=��*輈T��8K<���<�8= @T=p�D=$F�<`>�����l�1�߿�����wN������ǿ����c"�:�F�d�m�b���w��c���   �   B˟�����`���ji_�Y;����
�������܊�0�A����J��� #������Oݻ(X�<�*$=��=�C�<���;�����l5��Ȑ��:����罂f �X ��4�?��DŽm���Ѝ?�����P��;X��<�w=�=�,�<8��� ��V?&�^������u9C�tꋿ�����x��4A�@�;�Ҵ_������=������   �   �Ɏ�祋����sj���K�R�+������옭�fr~�wr0��n徱����(�r�� �$�<xG�<8/S<�	�����D���8����";��qV��4h��n��6i�VOX��=����i5��.���(��3��f,<��<(�l<xS2��|�J���.���s�7�1�>��lg����⿆��(�+��FK���i��<��sk���   �   �v��2q���b�F>M�:�3����q���K�ɿ�-��x�`�ٱ�(�Ǿ�fm����XV� �V���:�~��H�ӼX�y�q�ٽ�t"�cK[��}���z��\b���Rþ�ȾN�þ(���|��TQ���_�� &��-�ꒂ��D��λ�q)� �v�0)^�Q	����o��ɾtw��ma�����A�ɿ)o������3��TL���a��p��   �    �N��J���?���.��r���`5ڿ|}���샿i�>��+��\��RD��9Ͻt?�\ɮ������&�b?��ʼ�l�M�2׍�� ��O;߾ՠ�a��p<�������f��&��a��sa�����g]Q��������/�ܟ������tE�]`ҽ�E�#������>��ჿ�/��sٿ�i�`����-���>�HJ��   �   ��)�#'��������� ��ܿ굿�ˏ�T�X��@�բѾa����������J4�lE�<�N��������j�����޾�
��8(�,TA��3U��b�ǵf�|�b�f_V���B���)�������x쨾l7n�n����<�U������8�7x��/^� ����Ѿo��JX��4��I𴿞Hۿ~	 ����V���&��   �   V��~��d �84뿖jп᱿�ˑ� �d�l�*�Fn�����vH�h��誄���;�j�^�T ���K��s��&���U��u�!���H�[�n�����I���ϝ��栿`C���������p�b�J��+#�L������J�v�>Z�|����b��^>��s��]��T�G�8��eb��)�[4c��Ð�;���^�ο��鿃����?��   �   ��տ�ҿ�!ȿ�z��_��ǀ��(�_��-����;$��`�h�&&��q��t�X�EX�rX����*g�&Ұ�K���9,���]�^R��\���h'���ǿB�ѿ=�տj�ҿ�$ȿ~��!	��+���$�_�R�-������'��T�h�N)�u���X��AX�T��&��g�&ΰ������,�|�]��O��}���:$���ǿ��ѿ�   �   �㠿G@��������B�p�6�J�h(#�����o��7{v�V�F
����b��^>�v����轤�G�I;���f��)�38c�#Ɛ�������οu��I����A�V��t��> ��7뿕mп�㱿�͑���d�"�*�Fr�Ġ�H�v��Q���ΐ;���^�(���F�S�s�"���O��΃!�8�H�X�n�����F���̝��   �   ~�f�K�b�xZV�4�B���)�M������稾�0n����Y��� �U�r����8�6{�� a�`���k�Ѿ��)NX��6����~Kۿ% ����d��>�&���)�0%'����^��l� �*�ܿT쵿^͏�'�X��B�˥Ѿc��������:J4�T@�z�N�����e����j�5��� ޾��4(��OA��.U��	b��   �   x�������������\�����zVQ����k���T�/�����䗼�BvE��cҽ �E�|%��ք�p�>�yヿ�1��ށٿRk�����-��>�rJJ�t�N�`�J���?�l�.�>t��	��7ڿ9��-y�>�b-��^���D�*<Ͻ�?�H®� ��л&��6�� ���M��ҍ�*����4߾7��u��U8��   �   y�ǾH�þs���F���L����^�@�%��#�����-�P�ͻ�h(��v��+^������o��ɾ&y��oa�1����ɿnq����6 3��VL�>�a���p�vv�5q���b�"@M���3�"��c���ڃɿ�.��R�`�.���Ǿ�hm�6���$V���V�@̵:�8����Ӽt�y���ٽ n"�?C[�y��;u���\��vLþ�   �   ��n��.i��GX��=�C���*��%���(�@�2���,<8*�<��l<�S2��!|���70���u羲�1�<���h��V�⿂��b�+�^HK�j�i�>���l���ʎ��������juj��K�Z�+�ʀ�B��虭��s~��s0�[p従������r�������<�S�<�RS<������,;��U-彚��z;��iV�7,h��   �   *���/����F;Ž�x��x�?�`��� ��;���<x|=�=`/�<8��'���@&�q��������:C�7닿����z���A�6�;�
�_�����v>�����2̟�����a������hj_��Y;�������a���{݊��A�}��ܯ���#������Gݻ@]�<�.$=6�=S�<�"�;�⎼�^5������1����ca ��   �   �s��䲍��'w��=�T�h;��MK<���<�8=<BT=��D=�F�<xA�����M�1�����6���wN�)�����ǿ��bd"�̌F��m�xb��^x������@��t#��>l���,��B�l�:�E��V!�~� �%Lƿ�D��uL��)�q����M.���0�ƻ�r=(�M=Ht]=f�A=�z=�3q<�����i׼d�6���q��N���   �   "�Z�^P���/������c� e�;���<:�!=�S=fh=��Q=�) =��	��;����5�c>���W
�dVR�C.���V˿|��:%�8KJ��~r�-{��������E��'��M���t-���q��I��
$����[�ɿϔ�2BP�#��꥾72�7d��`���\�	=.[=�q=z*]=�@+=�,�<���;��C����d�*�"�M��   �   �s��𲍽�'w���=�\�(;� NK<(��<T�8=�BT=��D=`I�<H9�"����1���������vN������ǿx���c"�܋F��m��a��uw������?��y"��Zk��),���l�T�E��U!��� �OKƿ+D���~L��(������L.��
���ƻt=ڢM=�t]=��A=�z=�3q<І���i׼��6���q��N���   �   <���/����X;Ž�x��f�?�������;��<j}=n=X4�<��"���M>&���������8C��鋿����w���@�|�;�γ_�S����<�����Tʟ����`��2���:h_� X;�X���	��ɲ��?܊��A�������J#���� *ݻ�a�<*0$=�=�S�<�$�;�⎼ _5������1����va ��   �   ʧn��.i��GX���=�F���*��%��(���2� �,<|.�<(m<0>2�B|�����-��r��1����kf��u�⿴���+�zEK���i��;��Nj��^Ȏ�����ߐ���qj��K� �+��s�῭���sp~��p0��l�*���� ��r����$�<�W�<XWS<����� ;��^-彩���;�jV�P,h��   �   ��ǾV�þ����N���L����^�0�%�X#ཛ����*��ͻ d'���v��!^���)�o�� ɾv��ka�t�����ɿ.m��z��3�SL���a���p�Vv�0q�J�b�J<M���3����6���y�ɿ>,��/�`�%����Ǿcm�����dV���V� I�: &��h�Ӽʏy�n�ٽn"�JC[�y��Gu���\���Lþ�   �   ������������!��\�����TVQ����������/��������|kE�w[ҽܓE�� �������>�|����-��H}ٿ�h�΍��-���>��EJ���N���J�H�?���.��p�:��2ڿ�{��9냿��>�*�6Z��{�C�4Ͻ�>�ȴ��|��H�&�A6�����M��ҍ�2����4߾>��~��^8��   �   ��f�T�b��ZV�9�B���)�M������稾e0n���������U�r����8��r���Z�����ȘѾG�HX��2���Eۿ� ���Z���&�b�)�� '�����4� ���ܿ�絿�ɏ� �X�7>�3�Ѿx^��Ҕ�T}���?4��9�<�N�D�������j�.���"޾��4(��OA��.U��	b��   �   �㠿K@��������D�p�6�J�d(#�����S���zv�nU�1��&�b�>T>�n������G�5��G^���)��0c��������h�ο��ݬ���=�V������ ��0�qgпSޱ�fɑ�F�d�`�*��i�Z���dH��~�w�����;���^�(��dF��s�"���O��у!�=�H�`�n�����F���̝��   �   ��տ�ҿ�!ȿ�z��`��Ȁ��&�_��-�����$����h�7%��n���X��6X��M���g�lʰ������,���]�|M��ª��-!��9ǿ3�ѿ�տU�ҿ2ȿ�w��|��A~���_���-����� ��0�h��!�xj����X�P8X�%Q��B�g�ΰ������,���]��O������@$���ǿ��ѿ�   �   X�����f �;4뿘jп᱿�ˑ��d�b�*�%n�����H�Ӄ�Ҧ��@�;�ؘ^����3B��s����[J��a�!��H���n����C��}ɝ�k࠿*=�����+��9�p�ӴJ��$#��������tv��P���`�b�\R>��o��ܜ轖�G��7��Ob��)�^4c��Ð�?���c�ο��鿉����?��   �   ��)�
#'��������� ���ܿ굿�ˏ�N�X��@���Ѿ�`�����?����@4�6��N�������ˏj������޾���0(�KA��)U��b�=�f��b�{UV���B���)������$㨾)n����]���U�p��D�8��t��)]�����ǛѾh��JX��4��M𴿢Hۿ�	 ����Z���&��   �   �N��J���?���.��r���_5ڿ{}���샿b�>��+��\��~D�J7Ͻ�>�Ȱ��t����&��.������M�>΍������.߾������I4�U�������������ᾈV�������NQ����!�����/�8|������kE��]ҽ;�E��"������>��ჿ�/��wٿ�i�b����-���>�HJ��   �   �v��2q���b�F>M�:�3����p���K�ɿ�-��s�`�α���Ǿfm����V���V��Ͷ:�脻��Ӽ �y�6�ٽ�g"�~;[��t��p���V���Fþb�ǾD�þ��������G����^�`�%�c������@jͻ�&�@�v��"^�S��`�o�eɾmw��ma�����C�ɿ-o������3��TL���a��p��   �   �Ɏ�祋����sj���K�R�+�����옭�cr~�pr0��n�}���\���r������<4b�<wS<x��>��C2���"�^��n;�7bV�$h�^�n�W&i��?X���=����J�Z����'��2���,<�:�<�m<882�.|�����.���s�4�1�A��og��ü⿈��*�+��FK���i��<��tk���   �   D˟�����`��ﳁ�ji_�Y;����
�������܊�-�A�z��)����#�M���0-ݻ�d�<T3$=�=�a�<`l�;�̎��Q5�����(��d��`\ ����*���H2Ž�p��Dr?�$k���O�;���<,�=�=|9�<���h����>&�?���	���t9C�uꋿ�����x��8A�B�;�Դ_������=������   �   @���"���k���,����l��E�dV!�N� ��Kƿ�D��1L�Q)�1���ZM.�|��@�ƻht=,�M=�v]=�B=�~=�Hq<�T��<[׼0�6���q� J��o�����Nw�@�=��輠��eK<���<@�8=�ET=��D=`L�<�5����6�1�ҿ�����wN������ǿ����c"�:�F�d�m�b���w��c���   �   �߿��L��h��x@��?3���X�R�/�@���׿�����s`��F�_�����F�����y��H�<�zC=�>[= �E=�+=x��< �����`U���V��={��)��8�|�\�Y��"����`[=�L1�<��=�WA=T�V=@B?=��<���j�����H�ᶾ�7���a�������ؿN��j�0��Y���z���2��UQ���   �   Y������"'��wؖ������T�f�,�ނ	�Z4Կ�����m\�"u��᱾��B��m����{��Y�<D5=2F=Z)=P��<P�;�Mu�Dr��Bd�*V��N~�������I��͒��+h�X��tK����;��<\|$=�A=�1=d��<(���qO���D�}+���Z�E�]��ӝ�5Jտ�,
�&�-�N�U��Ȁ�z ���0���	���   �   ����RԪ�����7����q�oI��V$�`����ɿ����P��K	��V����6�X��h������<�	=��=d��<������߼ld��u����޽������~��E����+�Z����i�<�꼠&#�ۗ<\ =�4=���<Ա�����g8��y���
�+�Q��ŕ��ʿ�o���$��I���q��3���ɞ�ռ���   �   x����j���"���~��N[�vH8��9��m��ڹ������o>��9������b$�뒽����<(�s<�;������J�@ٲ�����+��O���l��� ��3����m��fQ�B.-���_,���Q�|�����k;��a<P��;����3I����%�e��<j��2?��$���a�����~k�dS8�f[���}���r?���   �   %����؂�(Hu��]�8�@�@~#�2���R׿?.��ؑq�#,'�;Dپ�܂�I0��u���T�� k�V�|��Ŗ�ٮ��R�5�v�r��������#�ƾ7cԾuAپ�Ծ�|ǾB������L�t��8��f�����Z� Zi�Ц�����w��,P��mھa�'��r��c���k׿,��<#��S@��l\���t�o����   �   ڶ^�,{Z�>N��k;�
 %�������m�������9aM�_��䝵��RY�T���m�����p'��l�T��p��Ƈ���c������Ǿ��*x���z|%�,�(�b�%��7�E,�����)ɾ���9Hf�2h�u����Y��� �hM�X�p��Dｼ%Z�����zM��u���K���c�
n��^$�"�:�$]M�vZ��   �   �6���2���)�I��	�	g뿏O¿�����i�
�'����3�� �,�������a�||9��K~���ӽ{�+�}x���<��%t񾓬�R�5��`P�cne���r�+�w��hs��4f��\Q���6����-� �������Q-��Aֽ/���w<���c���½�G-��J������['���h�O���O���j꿂��V����(��2��   �   j�x����������I޿������Uu���7�p���Q��^$]��������@�h��'����ӽ��,� 0���{þ}-�(�.��kX�U��r���������2��Q�����ƒ������Y�
�/����ľ}��4 .��ս�P���j�zޝ����3�\���M�L97��`t��O��H���)ݿ}������k��   �   kq俇��+�տm�ÿM$���-��:�o���:��:
�N���׼��0�,���&s��t<���M��ފ���~�^���;�	�A�9�&�n��c���=��4�¿U�Կ�X�@u�G�࿻�տ��ÿ;'��j0��v�o���:��=
�%���'��84�� ���s���:��I����|�~����\�	���9���n��`���:����¿��Կ)U��   �   ]/���M������0Ò���3�Y�]�/����ľ?���.�]{ս�M���j�᝽�����\�1���{O��<7�et�=R��2��Q-ݿ6������m������|��l���M޿�������Yu��7�����T��;(]������:�h��#���ӽ��,�i,��wþY*�C�.�4gX�XR��}��k	�������   �   ��w�&cs�X/f��WQ���6�T��'�9�������K-��:ֽ���6t<���c���½K-�MM��D��\^'���h�t������#m�H��\��$�(�N�2�*6�F�2�)��J�\�	��i��Q¿u����i�I�'����5����,������a�w9�vA~���ӽ��+��t���7���m�¨��5�\P�ie�4�r��   �   ��(��%��3�}(�M���#ɾ�
���@f��b��l���Y��� �VK���p�.H�)Z��
��!�3}M��w���M��)f返o�|`$�L�:��_M�$Z���^��}Z��N�n;��%�6�����G�������jcM��������JUY����4�m�$�������T��g�������c������Ǿ%��Mt���x%��   �   �:پ��Ծ�vǾ���������t��
8��[���홽L�8:i�8����;y�� R������ھ.�'�+r��e��~m׿d���=#��U@� o\�z�t�ۣ������ڂ��Ju��]���@��#�>���T׿�/��ԓq��-'�#Fپނ�q1�;v���O���<�V�*�����D����5�Ɍr�{�T�����ƾ�\Ծ�   �   ������d�m�V_Q��'-�N���"����P�Hz�� +l;��a<`��;�����J��{�%����nl���3?��%���b��a��l��T8�![���}�>���@��� ���k���#���~�FP[��I8��:��n��۹�Ȯ���p>�5;������c$��뒽�����<x�s<�_�;�q����J�@ϲ����y+�>�O��l�D���   �   �x�@���������x�i����@�"�|�<,a =.8=���<ܲ��M��yh8��z��]
�`�Q�fƕ��ʿ�p���$��I���q��4���ʞ�ݽ������Nժ�����8����q��oI�hW$����k�ɿ<����P�9L	�tW��,�6�PX��8��� ��<@�	=��=x��<@W����߼4]d��l���޽ԣ�X���   �   f����D��=Ȓ��"h����>�� /�;X"�<�$=2�A=�1=��<����zP��٤D�9,��n[��]�Aԝ��Jտ-
���-��U�ɀ�� ��-1���
��戻�W���'���ؖ�Z����T���,��	��4Կ����n\�Ou��᱾��B��m���{�]�<jF5=H	F=b)=���<�M�;�0u��i��9d�4Q��y���   �   �)��L�|���Y�*"������_=��0�<,�=~WA=��V=�A?=؎�<��������H�Tᶾ8���a�������ؿf����0�,�Y������z���2��[Q���߿��L��\��h@��/3����X�8�/�*����׿p���Vs`�pF����(�F�7���y� J�<{C=4?[=\�E=6,=��< �纤���6U�l�V��={��   �   |����D��GȒ��"h����>���/�;�"�<�$=��A=�1=���<|����N����D�=+���Z���]��ӝ��Iտ�,
�ޡ-��U�ZȀ� ��+0��y	��̇��C���&���ז�����T���,�~�	��3Կ ���m\��t�᱾��B��k����{��_�<<G5=�	F=�)=��<�M�;�0u�
j��9d�CQ��5y���   �   y�0@���������r�i�h��@�"���<.b =�9=���<Ԫ���� f8��x���
�f�Q�ŕ�L�ʿzo�&�$�(�I�v�q�3���Ȟ�ٻ������LӪ����"7��\�q�
nI� V$������ɿ�����P��J	��U����6�3U��L�����<	=��=|��< O����߼F]d�m��&�޽��j���   �   ������z�m�b_Q��'-�L���"��V�P��x�� Al;p�a<p�;x���TF���%�; ���h���0?�$��v`��U��j�<R8��[���}����'>�����^i��}!���~�M[�$G8��8��k�ٹ�����n>�e7��+��~`$�6璽| ����<(�s<�i�;Dp��6�J�8ϲ����y+�S�O�*�l�]���   �   �:پ��Ծ�vǾ���������t��
8��[��T홽���/i��������s���M�s���Xھ�'��r��b���i׿ ���:#�R@��j\�d�t��������>ׂ��Eu�F]�d�@��|#���
Q׿�,��n�q�R*'��Aپ�ڂ�m-�q���B�� �V������������5�ӌr���a���
�ƾ�\Ծ�   �   ��(��%��3��(�U���#ɾ�
���@f�Wb�l��,�Y�� �D�@�p�p?�`"Z����~�^xM�yt�� J��Ha迢l��\$��:��ZM��Z��^�~xZ��N��i;�6�$�F����T�������^M�p������NY�����m�Ď�����6�T�g�������c������Ǿ0��Vt����$x%��   �   ��w�0cs�b/f��WQ���6�U��'�+�������`K-�,9ֽ�	���l<�`�c��½hD-�`H��4��|Y'���h�d������Ag����j����(���2�J6���2�X�)�G��}	��c��L¿i����i�m�'���1����,�������a��o9��<~�D�ӽX�+�|t���7���m�ƨ��5�\P�ie�?�r��   �   c/���M�����4Ò���4�Y�\�/��s�ľ��.�9yսzJ���j��؝�F����\����J�a67�9]t�wM��� ���&ݿ������i�D�Z��~������F޿�ｿN ���Qu�]�7����@N���]�����|��`�h�q ����ӽ�,�?,��
wþW*�E�.�7gX�[R�����p	�������   �   qq俌��0�տs�ÿQ$���-��:�o���:��:
�(���H���/����=n���4��bB�������~������	�,�9�h�n�V^���7����¿/�ԿrQ࿟m�þ࿌�տ�ÿA!��6+����o�߸:�8
����G���+�s���tl���5���E������~�����V�	���9���n��`���:����¿��Կ0U��   �   l�|����������I޿������Uu���7�`���Q���#]����J��"�h����e�ӽ��,��(���rþj'���.��bX��O�����S��V���
,���J��ґ��<���o����Y�s�/������ľx��.��rս�F���	j�5ڝ�u��k�\���M�G97��`t��O��K�� *ݿ�������k��   �   �6���2���)�I��	�g뿏O¿�����i� �'���㾔3���,�������a�4l9�N4~��ӽ�+��p���2���g�#����5�JWP��ce���r���w��]s�*f��RQ�F�6����� ��������E-�1ֽ`���g<���c��½�F-�zJ��e���['���h�Q���R���j꿄��X����(��2��   �   ޶^�.{Z�@N��k;�
 %�������m�������2aM�Q�������QY����&�m�������@�T��^���{�H�c�o�����Ǿ���p�أ��s%�V�(���%��/��$�l��ɾ����8f�D\�%c����Y�,� �h@���p��A��$Z������zM��u���K���c�n��^$�$�:�(]M�zZ��   �   '����؂�(Hu��]�:�@�B~#�2���R׿>.��֑q�,'�Dپ�܂�:/�vr���@�� ��0�V����n���;���<�5�|�r��Ն����ƾbVԾg4پ/�Ծ�pǾ
������9�t�\8��O��G䙽X��@
i�Xm��	��vt��!O�����GھZ�'��r��c���k׿.��<#��S@��l\���t�p����   �   x����j���"���~��N[�vH8��9��m��ڹ������o>��9�����'b$��蒽d ���< �s<���;Y���J��Ų����\r+���O���l���� ��i���m��WQ�� -�P������P�\_�� �l;�b<�/�;L����F���%�1��$j��2?��$���a�����k�fS8�h[���}���r?���   �   ����RԪ�����7����q�oI��V$�b����ɿ����P��K	��V���6��V��4������<�	=��=�Ρ<�!����߼Od��d��Ĝ޽Ş� ���s��:�n~�B��v��v�i�<�꼠�!����<Bh =$>=�<����f���f8��y��|
�+�Q��ŕ��ʿ�o���$��I���q��3���ɞ�ռ���   �   Y������"'��wؖ������T�f�,�ނ	�[4Կ�����m\�u��᱾��B��l����{�``�<�H5="F=�)=���<�y�;@u�Db�1d�pL��t��;����?��NÒ��h�H���/���`�;�,�<�$=�A=1=��<�����N����D�n+���Z�D�]��ӝ�7Jտ�,
�&�-�N�U��Ȁ�{ ���0���	���   �   ���s���׵����t����Ga�t6�:�B߿S�� �h��;�������Q�2������K�<X�6=RoO=xv9=�x=0�f<��ƻ8/ռ@�3��,m�����w��9���m�i4��׼�cλ(Vc<�=p�8=��N=��6=��<�,������a�Q��Խ�3d��i������U߿T���V6�V�a��Ո�J'��ߵ��t���   �   خ����������v��օ���\�l�2�,!��`ۿ����d��O�๾�mM�羹�H����<�c(="�9=��=,$�<�0;,����*�^�{�鰝��"���?���R��o����|���+��%�� � ;0s�<�<=�(9=�(=@��<H3���׹���M�����t���d�}���]�ۿO��'3�t.]�y��Y�����j���   �   �����\���إ�=6��Rb{�<�P���)��G���пV���X�����﮾��@�	?���p���.z<<��<̀�<Xc�< 񷻖���|��4������k
����(�����T�Թ��~��9����d��<tP�<�;�<by<ফ��R���A�7��f���X�|����пh�6*��P��p{��3���ϥ��T���   �   �բ����j������mc�>�>��*�C����Z}����E������z�-��7��L컼}�;K3<�h:ɹ���b��/���F��5���Z�;x��������ƾ��W�x�8�Z�<�5�^�������Bd� 综 p�9A1<�2�;84��wF��>�-��'������E�����-��a���5��>�\c�l�������   �   �8���!��$�~�� e��]G�"�(�6��6޿N����z���-�%G������u��ȫ�h�@�ꑼ^�*�WF��'(��@��~�띾�L���Ͼ��ܾr�ᾶݾ�7ϾΒ��27��9�b�@���������+��P��h�B� �q ��r��"���U�N�-�h*z�!����4޿����(��4G���d�|�~�t���   �   �g�(sb�;U�:�A��/*��/�(�?o��0A��#�T�\��X���.d��>��uՂ� ���}��l�;	ͽ�#���o�袾�Iо����C�T�!�ң+��/���+���!��6�������оWE��;p�9$���ͽ��m����� ₽:��X'd�=S��W�W�T�5��}V�������)�J\A��U��Pb��   �   3<���8�R�.�f
 �X��1z�Mȿ��,�p�0�-���s���]+6���ϽB�x�4�O��^��,���L5�]����H��)v��H��џ<�X��m�
w{�� ��E�{���m��ZX��<���������������5�T�����` P���x�A�ϽG6������u�.�-��p�a̞��ȿq)��k�"����.�d�8��   �   ����+�R����h��۶ÿ>꠿tk}��=>����������g��������U�P9��B_�"`6�L���s�˾b��fQ5��v`�y��5������]���Wʱ�Է������wi���)����`��5�@���?̾Fʌ�<�6����v{����D橽#��Tag�VU��&f��>��}�T���lÿ5�俈� �����   �   �뿞�翡ܿ��ɿ
p���ʗ�زw��A�m:�Hɾ�}���'�Zν�֎�������ͽRT'�:N��(ɾ���@��Rw�쎗�,��`�ɿ��ۿ3��
��z��Iܿ@�ɿs��[͗�2�w�%A� =�Lɾ����~�'�νl׎�ﾎ��ͽ:P'� K����Ⱦ'��@�FNw�,����(���ɿ�ۿL���   �   �Ʊ�u���Q����f��-'����`�H�5�:���:̾�ƌ���6���⽩x��B��詽���fg��X���h�
>��}�᳠�oÿ���t� ���N���.�\��� ���俪�ÿ�젿Io}��@>�Ќ�Ї����g�2��J����S��5���X��Z6�����r�˾#��aM5�(r`����2���}�������   �   �����{�]�m�VX���<�N���������

��<�5��L�e�����O���x�z�Ͻ|6�V����y�؇-���p��Ξ�`ȿ�,��m�<���.��8��5<�:�8���.�j ���}�Pȿ��Eq���-�M�쾚����-6���Ͻ��x���O�SY��ޯ��F5�S���YC���o��X��E�<��X�z�m�Uq{��   �   /�0�+���!��2������о�@��r3p�J3$�c�ͽV|m�l�j��$ソ�=���*d��U���X��T��6���X��y�ￜ� �)��^A�(U��Sb��g��ub��=U�d�A��1*�81���(q���B��g�T��]��Z��$1d�A���Ղ�*���u���l� ͽȺ#���o��⢾�Cо����I ��!�N�+��   �   ���ݾ�1Ͼ���'2���0�K�@�����>�+�@��pwB�h��!��S���#��gX�'�-��,z�����7޿�0�(��6G��d�>�~����3:��J#����~��"e��_G���(�N�~8޿�����z���-�!I�:��������Ħ���@��֑���*�=��,"�@��~��坾	G��m�ξC�ܾ�   �   &���<����}x�c�Z�P�5�u��.���3d�Xϻ� ��9�W1<�I�;@4��	H����-�$)�������E�1���1/���b���6�x�>��]c����S��y��ע�_ ��������6oc�r�>��+��D��%��,~��՗E�������|�-�Z8��黼 ��;f3<��: ���J�b�8%���@�j5���Z�V2x������   �   7��
#�D��?K˹���}��-��ʿ�(Ѐ<[�<hB�<�gy<觫�T��
A�b��H��L�X��|���п�h�*�0�P�,r{��4���Х��U�������]���٥�7���c{��P���)�TH�S�п�V��ފX�e����Z�@�]?��@n��:z<$�<,��<�s�<����� ���|��+��;��V�����   �   7:���M��}���|���+����� ;|�<@=+9=$(=���<�4���ع���M�����u�c�d�������ۿrO�|(3�/]����ނ���������i���g������w��\օ�.�\���2�`!�9aۿO���8�d��O�=๾�mM�ؾ��x����<0f(=^�9= �=�.�<�u0;8���*��{�Ϋ��p���   �   �w��9��2�m�Li4� ׼�eλ�Tc<��=�8=N�N=x�6=��<0.�������Q��Խ�dd��i�݈���U߿l���V6�v�a��Ո�Y'��ߵ�u�����s���׵����c����Ga�X6�$�߿�R����h��;�s�����Q��~�����<L�<��6=�oO=�v9=Zy=x�f<p�ƻ�.ռ�3��,m�����   �   G:���M������|���+���`� ;d|�<B@=�+9=�(=���<�0��3׹�H�M�~���t�T�d�G����ۿ�N��'3�.]�-������x������I���K����(v���Յ��\���2�� �N`ۿ����)�d�O�;߹�nlM�$���(���p�<g(=ا9=8�=�.�< v0;H��0�*��{�߫������   �   K��#�X��^K˹���}��-�@ȿ�Dр<]�<�E�<pry<�����P���A�r�����F�X�z{��;�п�g��*�2�P��o{�*3���Υ��S������p[���ץ�Z5���`{�$�P�$�)�4G���п7U��وX�������@�+<��f��xDz<\	�<(��<u�<����� ���|�,��Y��f�����   �   3���I����}x�t�Z�\�5�u������2d��ͻ� l�9�`1<Pf�;�(���C��{�-�w&�������E�K����,���_���4�ޚ>�~Zc�f��������4Ԣ�����������kc�ښ>��)�cA�����H|���E������� �-��3���ݻ����;o3<�*:������b�%%���@�x5���Z�r2x������   �   ���*ݾ�1Ͼ#���/2���0�F�@�j���򤽴�+��:��hfB��⼋��*��� ���S�΋-�[(z�ǵ��G3޿��@�(�
3G���d�؉~����7��P ��f�~�6e��[G���(����4޿����2z��-�nD�����������س@��ё��*��<��"�
@���~��坾G��~�ξW�ܾ�   �   /�;�+���!�3�����!�о�@��X3p�3$���ͽ�ym��	����W݂��4���#d��P��XU��T��3���T��x�ￎ	�L�)�&ZA� U��Mb��g�Vpb�h8U���A��-*�..���m��u?��v�T� Z��U��W*d�
8���ς�����p�(�l�5�̽��#�x�o��⢾�Cо����O ��!�Z�+��   �   �����{�g�m�VX���<�P����������	��׷5�RK����*�O�0�x�~�Ͻ�6�G���yr�ӂ-���p�gʞ�Jȿ�&�Bj�"��v�.��8�z0<�B�8���.�P ����w��JȿZ��p���-��쾌���'6���Ͻښx�8�O��V��z�⽖F5�;���OC���o��[��K�<��X���m�bq{��   �   �Ʊ�{���V����f��0'�� �`�I�5�7���:̾�ƌ���6����$u��*t�K੽�~��\g�R���c��>��}�����>iÿ��俲� �����l���)�>������ܳÿ�砿Bg}�s:>�������*�g���������H�2��QV�LZ6�l���]�˾ ��aM5�,r`����2���}�������   �    �뿥�翧ܿ��ɿp���ʗ�ڲw��A�d:��Gɾ�}��
�'�/ν�ю�����ͽ�K'�H����Ⱦj���@��Iw������%����ɿw�ۿy��/�뿿���ܿp�ɿ�l��ȗ�1�w��A�n7��Cɾhz���'�oν�ώ�޹����ͽ@O'��J����Ⱦ��@�HNw�/����(���ɿ�ۿT���   �   ����+�V����l��ܶÿ>꠿sk}��=>���������g����]���rH�B/���P⽶U6�����˾���I5��m`��/��mz������{ñ�������}c��q$��7�`�E�5�����5̾Ì�̲6����jq��r��᩽Ā��`g�U��f��>��}�U���lÿ9�俋� ������   �   3<���8�T�.�j
 �Z��5z�Mȿ��)�p�'�-�ۗ� ���C*6��Ͻ�x�x�O��R�� ��)A5�~���c>��fi������<�	X�$�m��k{�����{���m��PX�$�<�`��)���У������5��B㽽�����O�r�x���Ͻ)6�l����u�'�-��p�b̞��ȿt)��k�$����.�f�8��   �   �g�,sb�;U�<�A��/*��/�,�Ao��0A���T��[��X���-d��;���Ђ����hj��yl���̽ƴ#�ڐo�)ޢ��=о�}��m��͖!�ޚ+�}/���+�X�!�/������оq;��=+p��,$�V�ͽ�lm���.���݂�17��x&d� S���V�R�T�5��}V�������)�L\A��U��Pb��   �   �8���!��(�~�� e��]G�$�(�8��6޿M����z�|�-��F⾴�������d��ء@�0�����*�4��x��@�X�~�����[A��:�ξ��ܾ���{	ݾd+ϾC����,���'�Ҕ@�l��a餽��+��'���NB�����`���!���U�F�-�g*z�!���5޿����(��4G���d�~�~�u���   �   �բ����k������mc�@�>��*�C����Z}����E�ܲ�r����-�n5���ݻ�pљ;p�3<�P:����`�b�o���:��5��}Z��)x�����󈾸���ux�l�Z�4{5�M�������!d�賻� E�9�{1<���;�%��D���-�r'������E�����-��a���5��>�\c�l�������   �   �����\���إ�=6��Rb{�>�P���)��G���пV���X�����﮾;�@��=��g��`Jz<�<̙�<�<�L��r���|�q#�������N�����~����nA¹���}�� ��s����<�i�<�N�<X}y<p���&Q��)A���_���X�|����пh�8*��P��p{��3���ϥ��T���   �   خ����������v��օ���\�l�2�,!��`ۿ����d��O��߹�]mM�*�������$�<dh(=D�9=��=8�<��0;����0�*�ڕ{�䦝�A���4��wH��k����z|�L�+�$	��@c!;���<�D=�.9=\(=转<�.��׹�n�M�����t���d�}���^�ۿO��'3�v.]�z��Y�������i���   �   �3���������j���C��F�`�f�5�~N���޿M ��:�h��vv��e�Q�Qz��H����P�<Nh6=��N=P�8=�=�7f<�
ƻ�NԼ޷2��k�����1��e���Zj�N�0���ϼ0���@
q<��=��;=��Q=f�9= �<����Ÿ����O��b���\�ªg�#����޿����V5�NG`�|��mL��m���,����   �   �����+���߰��ɜ��\���c\���2����ۿ�M���Yd�}����@M�*�������x�<b�'=`9=�s=@{�< $.;�à�`f*���z�ꜽ���H׷�ޢ���%��Ԕx���'��p����Z;>�<�k=r;<=
?+=���<l���+����K�5����t���c�	ɡ��uڿ؍��52��\��6��)����ٰ��,���   �   9۵��y�� �����pgz�&P�p�)���eп���#1X�Š�̱���@�e$��@«���x<,#�<<��<��<@e������[|�%Ǹ�L�&�0R������ٲ
�.��_���Yy�v��� ����<��<���<�<lQ�������+?�ҿ���
�jxW����x�Ͽf��>A)�:�O��Fz�������H����   �   2��?.��-Q���p��tqb���=�R����������0��0E�8s�R͝��-�����㻼p$�;`[2<�,:x���4�b�W����� �4�@ Z�zrw��$��V��U���p�v��<Y���3�)
�v2���g_�Xp�����:�F?<�;�2��]ɝ�TM,������� ���D�ތ��J���P������=�N�b������m��_B���   �   �����q���g}���c��mF�
(��
�z�ݿ4���ny�'-�ӹ� ʈ�p���Ï��&�Py@�PǑ���*�A!����B�?��@~�����฾�kξ@4ܾ��ྣ�۾�ξ�]�����P}��>�L�C[��؊'�������3��nڼ�����q�n(��� �^�,��y����fݿt�
�+(���F�x>d���}�����   �   �$f��^a�> T�P�@��W)�$���ￕ���Q�����S�
�������{c��q��_������,l��̽ �#�ENo�������ϾP��'���2!��+��p.���*��� �\[�'W��;Ͼ���b'n�P�"��˽�+i��G��I�〽W���ޔb�7G������S�,��������E�:���)���@� tT�,�a��   �   ^�;���7��.�n6�\���H�o^ǿV=����o�*�,�����	��k5�i�ν2\w�`�N��ۊ�� � �4�򃇾���L��o�N<�1�W��m�Ƕz�KR�'�z� �l�*W���;����A��JP�������4�+�ི����xL�THu�:�ͽV�4�0Ȗ��t뾘�,�p��b����ǿz��v0�t���g.�F(8��   �   �4�����
�*u �1�㿈�¿��3%|��M=�>��u���'kf���
�jި���}�f���w���5��/��}v˾W�45�^`�������"���#���,�������ߤ������h��%�_�o�4�~�
���ʾ�͋�rL5�|���ő��u|�3Z���
��Hf���� ��J�=���|�xd���ÿ:俾� ��F�����   �   ���߿�
ۿ��ȿlw��A�Ov��@��j��Ⱦ����Ol&��n̽䇍�@�����̽I�&�$ۄ��rȾ����o@��v�T��k豿�6ɿ<iۿ��濰�꿵�濦ۿ7�ȿhz������bSv�P@��m��!ȾF����o&�?r̽̈��o���ې̽<�&�؄�7nȾ����k@�m�v�CQ��H屿�3ɿ�eۿ����   �   >)�������ܤ�����Qf���_���4�|�
�'�ʾ�ʋ��G5����Ñ�Ju|��\����
��Mf����������=��|�g���ÿ�=俪� ��H�ڲ��6�ҏ���w �q��W�¿b��)|��P=�s������,of���
�਽��}�db��qὼ�5�E,��~q˾�S�25��`�Ի���얿���6 ���   �   �L��{z�Įl�2%W�>�;�Q���;��dK������)4����E����tL�xIu�o�ͽ��4��ʖ��x�=�,�}p�e��)�ǿ���J2�����i.��*8��;�H�7�.�n8����K��`ǿN?����o�z�,������m5���ν�[w��N�?֊�@��4�����������-k�zI<� �W�'m��z��   �   Sl.�Z�*��� �~W�QP��:5Ͼ����n���"��˽L i�LA��G�%䀽����6�b��I��֨���S�籑��¾�_H�и���)���@��vT���a��'f��aa��"T�v�@��Y)����Y����ӽ��� T���� ļ�n~c�Zt��6_��"����dl���̽�#�.Fo�樢���Ͼ8��.���.!�W+��   �   ����۾�ξX���	���}�
�>����R��r~'�t���p�3� mڼ⍽�s�*��p�3�,�wy�����hݿ��
��,(���F��@d�H�}�����#����r��~j}���c��oF�l(��
�4�ݿs5���py��-�л�Tˈ����<ď��!� b@�@�����*�������?��7~�c���(ڸ�=eξ�-ܾ�   �   xQ��������v��4Y���3�.#
��(��X_��X��@��:�\?<���;�2���ʝ�O,�]��� �@�D� ߌ�AL���R����J�=��b�����Fo���C������/��eR���q��sb��=�<�����Ԥ���1��71E�t�NΝ�$�-���@໼`E�;�v2<��:�⹼��b�����
���4�?�Y��iw� ���   �   �������
����W��bKy�b���u��\�<� �<p��<쾃<�R�����-?��������yW�Ҧ����Ͽ��B)�R�O��Gz�������X���Jܵ��z����Ɉ���hz��&P��)���vfп*���1X�M��s�����@��$�� �����x<�+�<���<�ǁ< ����:L|�M���l�?!��L��   �   �ѷ�����!��΋x���'�8c��`3[;G�<�n=�=<=j@+=x��<����2��~�K������u�E�c��ɡ�wvڿ>��J62��\��6������Kڰ�m-������V,��[��Eʜ�2]���c\��2���jۿ�M��BZd���:���6@M����������<��'=� 9=�w=���<��.;�����]*��z��䜽5���   �   �1��p���4Zj�r�0�l�ϼ����	q<T�=�;=R�Q=��9=�
�<h���X����O�
c��"]���g�H����޿
���V5�lG`����~L��z���3����3���������j���C��&�`�J�5�fN���޿( ����h���2v����Q��y�������Q�<�h6=��N=��8==�8f<`ƻ$NԼ��2���k�����   �   �ѷ�����!���x���'�4c�� 4[;XG�<>o=R><=@A+=$³<�������,�K�󝸾�t�8�c��ȡ��uڿ����52�|\�:6��ų��Bٰ�R,��b���;+��P߰�\ɜ�x\���b\�:�2����~ۿM��3Yd���5����>M�g�������d"�<��'=!9=
x=��<��.;����]*�,�z�圽L���   �   ������
����W��hKy�F��`s��p��<��<���<ă<\J��⟬��*?����+
��wW�x�����Ͽ���@)�Z�O�REz�솒�"��C���'ڵ��x���� ���fz��$P���)�h��dп����/X�ߟ�����6�@�v!������ �x<4/�<���<�ȁ<P�����:L|�Z�����P!��L��   �   �Q��������v��4Y���3�4#
��(���W_�@W���ǩ:�e?< س;�'��rƝ��K,������ �v�D�>݌��I��lO������=���b������l��A������,���O��o���ob�p�=�>��ʤ��_����/��j.E�r��˝���-�����Ի��b�;�2< �:Ṽ&�b������
��4�P�Y��iw� ���   �   ����۾�ξ#X���	���}��>���QR���|'�`�����3��_ڼ�܍��o��&�����ߧ,��y�����dݿb�
��)(��F�F<d��}��������
p��$e}�,�c�lF��(�Ș
�z�ݿ~2��ly�J-���+Ȉ����߾���ἘP@�讑�l�*���������?��7~�l���5ڸ�Meξ�-ܾ�   �   ]l.�d�*��� ��W�\P��A5Ͼ����n�X�"��˽�i��<�L@�aހ����o�b��D��<����S�������eC�ȵ�N�)�`�@��qT�j�a��!f� \a��T��@��U)����\�o���������S�������wc�\k��eY�������tl��̽�#�Fo�ᨢ���Ͼ@��5���.!�b+��   �   �L��{z�Ѯl�<%W�E�;�T���;��[K�������4�s�������mL��=u�|�ͽ��4��Ŗ�Fq�@�,��p��`���ǿ���.�t��Fe.��%8��;�X�7�n.�Z4�����E��[ǿ';��/�o�|�,�ơ�����f5���ν�Ow�b~N��ӊ��⽩�4�����������-k�I<�(�W�2m�!�z��   �   E)�������ܤ�����Vf���_���4�{�
��ʾlʋ�:G5���མ���Dj|�:T��E�
�Df�Ġ�����I�=��|�b���ÿ�6�� ��D����r2�z��|�Ds �˰㿏�¿~��!|�oJ=���������ef�v�
�sר�~�}��^���n��5�,��eq˾�S�15��`�׻���얿���= ���   �   �����
ۿ��ȿqw��D�Ov��@��j��ȾG���Zk&�fk̽悍������̽ȑ&�	Մ�jȾ٫�|h@��v��N��KⱿ10ɿ�aۿ)�������Rۿq�ȿRt���nJv�	 @��g�$Ⱦ-���Cg&��f̽���\�����̽<�&��ׄ�nȾ����k@�n�v�EQ��K屿�3ɿ�eۿ���   �   �4�����
�.u �5�㿌�¿	��3%|��M=�0��?���[jf�N�
�ڨ�T�}�\��*i�|�5��(���l˾�P�k�4�`�5����閿_������%��7���J٤������c���z_��4�B�
��ʾ�Ƌ�
B5�ߡ�ٻ��$h|��U��~�
��Gf�ԣ����B�=�݈|�xd���ÿ :��� ��F�����   �   b�;���7��.�r6�^���H�r^ǿW=����o�!�,���뾊	���i5���νQw��zN�vϊ�~�B�4�|���񽾍��mg�E<�:�W��	m�}�z��F��uz�_�l�/ W���;�l��C5��!F�������4�$�ཨ���hL� =u���ͽ6�4��ǖ��t뾎�,� p��b����ǿ{��v0�v���g.�J(8��   �   �$f��^a�B T�T�@��W)�&���￘���R�����S���������zc�o���Z����r��F�k���̽�y#�y>o������Ͼd
��T��[*!��+��g.���*�^� ��S�JI��./Ͼ����n��"���ʽ�i��4�z<��ހ�s�����b��F��ئ���S�-��������E�:���)���@�tT�0�a��   �   �����q���g}���c� nF�(��
�}�ݿ4���ny� -�����Ɉ�`��W���L��>@�p����*� ��L����?�/~�_���~Ը�_ξ'ܾ��u�۾D�;LR������
}���>����I��Po'�Hq���3��Zڼ3ݍ��p�(��� �U�,��y����fݿv�
�+(���F�z>d���}�����   �   4��?.��-Q���p��vqb���=�T�����������0��0E�,s�͝�b�-����Ի��x�;(�2<�
:(ɹ���b�A������4�}�Y�Raw�����L��Q�P�v��,Y���3�
�u��&G_�`=�����:Ѐ?<0��;P$���Ɲ��L,������� ���D�ތ��J���P������=�N�b������m��_B���   �   8۵��y�� �����rgz�&P�p�)���eп���"1X����������@��"��ȸ�� �x<6�<\��<�ׁ< �������=|�Ե������G�R��n�R�
����;N��<y�x������ �<�<x��<�Ƀ<H��)���&+?������
�hxW����y�Ͽf��>A)�:�O��Fz�������H����   �   �����+���߰��ɜ��\���c\���2����ۿ�M���Yd�|������?M�e������#�<��'=x#9=z{=��< �.;`����U*� �z�������̷�f������~�x�:�'�pT��`�[;�Q�<ps=�A<=�C+=Xų<М��e��R�K�%����t���c�	ɡ��uڿڍ��52��\��6��)����ٰ��,���   �   h0��!��������Y��f����FW�0�.�`,�W�ֿb��!�_�A���봾�}F���� w~�l��<(jA=~*Y=�C=�=�ؐ<�<�x櫼���<�R�p�u��s��̳s�VO��'���� ̃�t�<L_=p�J=`&`=D�H=���<PxY�X����	C�<����D��]��ߝ�e`տ�F
���-�4IV�w��n�����e����   �   ����r��ȧ�����O~��/S�t�+�
��hJӿwQ��m{[�����<���@B��d����� ��<P3=�D=<M'=d��<���;�ht���f�a�w!��>[��u����W���?���k\�f� {Z��<t��<F2.=�K=��:=���<��[������>�����{�$�Y�f1��'�ѿ �2�*��UR�T�}�����ӻ��"v���   �   �����O��l����N��,o�ڝG�l.#�/�c�ȿ�Q����O�������D6��!��\��<Ǚ< �=FR=t��<���%༪uc��K��w�ܽ�$�H��������
���ٽ�ަ�J(\�MѼ e�94b�<t
=@,=�<�<Йg�����3������k��&N��a����ǿ��<�"�G���n��P��x����h���   �   }ҙ��!��_����iz�p�X�zZ6�������F���Zȇ�r<=�ܾ���E��
�#��o��({��hw<�o<���;�����J�4[��FG�rx*��PN��j���|�X<��B�{�,i��uL��[(�N �
����B�$J���3�;��<��)<ॄ��T� ��������E<�����ַ�{��x���C6���X���z�l;���P���   �   ������x�q���Y��/>��!�*n�>Mտ������o���%�y�׾C��>�@����H��PW�H,W�����r�������J5�uq����xR��e�ľ&Ҿ��־�Ѿ�ľ8�������n��2�V0���6�����(;�`巻�D����}�t�����8־%�G�n��a��?տ(w�^�!�D�>���Z�T?r��)���   �   \��wW���J���8��"�n�
���Ck�� ���qIK����峾@LW�qb��%k����8�����S�H�����;c��
��Ͷƾ=�V��Ll��#�� '�0�#������
�Uj�^�ľ(k��2@`�b��o���j�L�h�����e��,��U�� ��6"�6�J���L���>��Zu�DP#��k9�n�K� �W��   �   Z4���0��)'���lq� �h��������f��{%�q�ྫྷr��K�*�u0����]�^�6��x{�fҽP�*��Ȁ�Z���P�����4��O�h�c���p�Wu��Ep���b���M�l�3���uL�������~�;�(���ν
9v��2���Y������)������8�%�sf��Z��FX�����%���T�'��1��   �   B��@���������ڿ��^����q�b!5�I� �����r�Y�D��[H����c��˄�|4ѽxQ+�5���C¾'p�ڵ-��^W�}^��B���򞿽����g�� 9��JR���{�� �}�2�U�V|,�.}�����;7����)��1Ͻ�G��:&a��W���;���Y�^����5���r�Bf������ܿ�R��$;�BE��   �   #��޿؝ҿ����O_���Ð�H�k���7�i���T���z���%��tB�2��&����p�|�]8��Q����8�p[m����j������{ӿ��޿�&⿇޿[�ҿ���/b��Ɛ�y�k��7����X��W{�`���(��>D���������l�'|�!4��z��ڥ8��Vm�E����g������+xӿ�޿�   �   _d���5��5O���x���}���U��x,�Hz�K���4��F�)�],Ͻ�D���%a��Y��]>�~�Y�������5��r��h�����M ܿIV��&=�^G�b��R�������2�ڿ���������q�B$5�j� �����N�Y�t���I����c�QȄ�.ѽ�L+��1��?¾m���-�4ZW�/Y�@��_s����   �   �u�J@p�w�b��M�8~3�p���F�
�����~��(���νl0v���1���Y�� ����)��
��?��Ċ%�svf��\���Z���鿤'�����'��1��4��0��+'����s���ä�������f��}%�����t����*��2��@�]�"�6��n{�hҽ��*�ŀ��T��MJ�O��M�4�O�"�c��p��   �   <�&��#�����
��c���ľ�f���8`�Ԃ�f�����L��|�����e�0�R�U�h��$���J���b���Ǎ��v�R#��m9���K���W��\�<zW���J���8�Ρ"���
��m��w ���KK�����糾�NW��d�:&k�ܒ������NtS�i���	��lc����ƾC6񾁆�%h���#��   �   *z־��Ѿ�ľ���I���B�n�@�2��%��I.�����;�@·��B����}�:�����t:־�%���n�Sc��+տXx���!��>��Z��Ar�+�����M���q���Y�>1>�:�!�6o��Nտ𾣿��o��%�b�׾q�"@������C���)�hW�l���i��c���\C5�llq�����L��E�ľ�Ҿ�   �   �7����{��#i�LnL�BU(�� �� ��țB�<3��pv�;�!�<��)<Х����� �j��������<����Eط���~��E6�D�X���z��<��R���ә��"�������kz��X��[6������V���'ɇ��==�i����F���#�Rp��x��`�<P�o<��;�����J�JQ��TA��q*��HN���j��|��   �   ��R��n�ٽ�֦�@\��5Ѽ �9xp�<(y
=�/=�?�<țg�����3�γ���l��'N��b����ǿ����"�G��n��Q��i����i�������P��K����O��No���G�/#��/��ȿBR����O��������6��!�����̙<J�=ZX=��< ɷ����fc�C���ܽ��߰��   �   I����R���:��$c\����`Z��<$��<�5.=DK=�:=d��<��[�������>�`��a|�߶Y��1����ѿ~���*� VR��}����\����v��u��,s���ȧ�P��"P~�0S���+�>���Jӿ�Q���{[���+=���@B��d��D��L��<nR3=$D=PQ'=��<��;�Kt�l�Bxa����V���   �   �s��ҳs�$VO� (����� ꃹ��<�^=�J=&`=��H=<��<�{Y�鄩�4
C������D�T�]��ߝ��`տ�F
���-�RIV�+w��}�����k���h0����������Y��W���tFW��.�J,�.�ֿ>���_���[봾(}F���8t~����<�jA=�*Y=j�C=L�=Dِ< 3��嫼|���R�X�u��   �   [����R��;��8c\����`Z��<\��<�5.=�K=��:=��<��[�;�����>�f���{�ܵY�31����ѿ�
���*�"UR�ʤ}�A���b����u��`��r���ǧ�u���N~�/S���+�����Iӿ�P���z[�Q��/<��}?B�c��������<JS3=�D=�Q'=��<���;hKt�f�Rxa����.V���   �   *��b�����ٽ�֦�T\��5Ѽ '�9dq�<z
=1=�D�< �g����p3�����lk� &N�?a��D�ǿ�����"�BG���n�P�������g������N��y���+N���o�МG��-#�t.�a�ȿ�P����O����ޝ��p6���� ���љ<��=\Y=��< ����༶fc�"C����ܽ�����   �   �7����{��#i�anL�QU(�� �� ��x�B��1�����;&�<��)<蚄��썽�� �ݧ������<�����շ�'����B6�&�X���z�K:���O��+љ�; ��,����gz�ĉX�*Y6������󑸿PǇ��:=�����D����#��k���l��x�<8�o<���;�����J�%Q��PA��q*��HN���j���|��   �   ;z־ϜѾ�ľ���S���M�n�D�2�j%���-�������:������5��J�}�B������5־�%�P�n�`���տ"v��!���>��Z��<r�C(��4������q���Y��->�p�!��l�MKտ���6�o���%�ڡ׾`<�����86������V��~�Vi��#���PC5�ilq�����L��T�ľ�Ҿ�   �   F�&��#������
��c���ľ�f���8`��������ԪL��s꼼���e�'�ʐU������ ��J���w�������s��N#��i9��K�n�W�r\�uW��J�d�8�P�"���
�2
�-i��T����FK����⳾,HW�&\��k�@���`���XqS��������Lc�
���ƾG6񾅆�-h���#��   �   �u�X@p���b��M�@~3�u���F����p�~���(�>�ν,v���1�x�Y�)��L�)����I����%�pf��X���U���:$����2�'�4 1��4�f�0�T''����o����۟����2f�y%�����o��&�*��)����]���6�j{��ҽ)�*��Ā��T��FJ�N��P�4�O�+�c��p��   �   dd���5��;O���x����}���U��x,�Hz�:����3����)�I*Ͻ�A��4a��Q��&8�Y�Y�.ꬾQ	���5�E�r��c��	���ܿO��29�2C�$��*��ĩ�������ڿ0�����q�05�ڼ �����Y�6���A���c��Ą��+ѽ�K+�O1�� ?¾m���-�2ZW�2Y�@��dy����   �   
#��޿�ҿ����S_���Ð�N�k���7�d���T����z����!���8�:����eh�U |�,0��ד�v�8��Rm�ç���d��y����tӿ5�޿@�޿K�ҿ����Q\��������k��7�����P����z�"��a��(5�ȋ�p����k��|��3��n��ե8��Vm�E����g������1xӿ�޿�   �   F��D��«�����ڿ��c����q�`!5�=� �������Y����$D���c�)�Y&ѽmG+�.���:¾j�S�-��UW�T�-=��L잿8���a���2��L���u����}�B�U��t,�,w�m���M0����)��#Ͻ�=��"a�4S��H:�'�Y��n���5���r�Bf������ܿ�R��&;�FE��   �   \4���0��)'���nq��k��������f��{%�K��^r��;�*��,����]�.�6�|a{��ҽ�*�f���5P��LD����4�XO���c���p�Du��:p�A�b�7�M��y3����C@�������~��(�6�ν�!v�T�1���Y�-����)����g��-�%�sf��Z��EX�����%���V�'��1��   �   "\��wW���J���8��"�p�
���Ek�����mIK���n峾nKW��_�(k�4���ܩ���fS�y|��5����b�g��E�ƾ�/�Ƃ�d�o�#���&��|#�¾�*�
�]���ľ�a��1`��|�ϊ��p�L�Pd�L��e��)�=�U�� ��%"�/�J���M���>��Zu�DP#��k9�r�K��W��   �   ������z�q���Y��/>��!�,n�?Mտ������o���%�R�׾�����=�𝂽�4�������V��r�a��K���~<5�#dq���\G��M�ľLҾ�s־h�Ѿ�ľ-��W�����n�"�2����%��v����:� t���0�� �}�b������7־	%�C�n��a��?տ*w�`�!�D�>���Z�T?r��)���   �   ~ҙ��!��`����iz�r�X�|Z6�������I���[ȇ�o<=�¾��~E��N�#�sm���l����<�o< =�;􇒼��J��G���;��j*�gAN�z�j�Cy|��3���{��i��fL�vN(��	 �����~�B�������;(3�<��)<����1퍽�� �˨��g���><�����ַ�|��v���C6���X���z�l;���P���   �   �����O��m����N��.o�ܝG�n.#�/�d�ȿ�Q����O���������6� ������ԙ<.�=�^= �<����T�߼�Xc��:����ܽ����������n ��ٽDΦ��\��Ѽ :�9\��<�
=Z5=J�<��g�!��3������k��&N��a����ǿ��:�"�G���n��P��x����h���   �   ����r��ȧ�����O~��/S�t�+�
��hJӿvQ��l{[�����<��h@B�d��d�����<�T3=�D=�T'=��<��; 1t����oa����Q��3����M��(6��"Z\���8DZ�x<t��<�9.=�K=�:=��< �[�$�����>�����{�"�Y�g1��'�ѿ �4�*��UR�T�}�����ӻ��"v���   �   �)��D��_k���Z���m���F�hp"�Ң��
ȿ����`�N�r��<褾�1��ؓ��Eڻ�M=�IV=Ʀl=�X=�t'= ��<p��;��@��j�X�$�tE���N�@�A�(*���ӼX���p<x%�<f�2=�Sd=(�x=��b=�g=�KM������,�ʡ�f���!L����oƿ�u ��'!�&SE�~�l�����I��B���   �   =��6����Z����h���B���������Ŀ2���J��%�}v����-�4f���uݻ���<�I=^�X=ȳ==2�= �g<�TǻD�Լd�2��`k��t��<���څ�*`e�>�*�|-�� Ea����<��=�I=6�d=LU=�[=`oW�>B��P�(��r��	>�uoH�,�����¿���P����A���g�<!���ؗ�T;���   �   ����X��������}��S[��8�ܮ��x�lۺ������?�����1���Z3"�����@��Df�<�/ =��=G�<0�;4q����4��G���D��X��M��z� �!x����߽d����͉��(�P�q�@<���<��'=<L,=��<�d���D~�˹�Mє�
����=�AG��Q`�����`����7�|�Z���}�����x���   �   暋��V����~�d,e��yG�"�(�
q��߿�~���}{�{.���fA��0����q��m�  �<|��<(HH<`y����施#��S��8���R��wc��h��Ub���P�(�5�����ܽ���z�G����x<P2�<�Ț<PZŻF@d�5�����R���,���y�{����޿����(�b�G���e���;����   �   8q���k�\X]��yH�\�/���BB��]Qƿ2ᗿ�n]�F���žf�j�g����T�$W�@�: ��4�ռ�}y�l�ؽ�}!�2�Y��"�����6����ο���þ���$M��8������bU�7u��hѽZ�k� ټ���ͺ�hz;�+���H�}���g�cþe���Z\�/i���ƿ�_���\���0�gI��E^��Dl��   �   ��J�|F�fW;���*���J6���տ�:�����-i;�����������@���˽�~;��T������΋%�d7����'L�ǌ��t���ݾ)  ���L����J0�#�q����fھ�Բ��Z��2�G��1�;����M���Ø�fV2�8ǽfo>��o������]�:������x����ֿ<�������+�&U<�`G��   �   ��&�p�#���&�����[�׿Sӱ������TT���<X;̡���0�Q����.�l/
�ܲJ�5?��rZ�R�h��A��?8ܾ#�
�&�#4?�EnR��^��ub���]�+Q��=�;�$�'	��Hپ1΢�Ҍd��5�@2���UB����S(�N���������;�&�l�T��<���β��ٿ?���F����2A$��   �   �~����d����w=˿Hn���,���_�Ƅ&�ł�Ȳ����B��B��7���3�JzW��3��.��8�p��4��|���* ��G��rl�e���Tz��$���������f���ٙ��h2j�"�D�N�X(�"����m�L��_���ڧR��0�L�|����޲B����Bl�ca'�jn`�o<��.ۮ�P�̿R������k��   �   �Tҿ�cο��ÿ�����ҝ�ԅ�Y�Y���(�!���uꬾmYa�����8�L�qM�����'�	���b��?��Q���:*��[����TA���d����ĿPϿtXҿmgο	�ÿ����=՝�eօ�C�Y���(�����\^a�D���Ş���L��mM�Ĺ����	��b��;������6*��[�!��z>��{a��=�Ŀ�Ͽ�   �   ����������1����-j��D��J��"�n����m�(��1���̢R��0�֋|�����B�����p�Yd'�3r`��>���ݮ�k�̿�U翓����m�܀�����g��f��f@˿�p��/��,_�w�&���뾐���N�B��F὾:��3��sW��-�������p�`0�������
 �V�F��ml�����^w�����   �   �pb���]�@&Q���=�O�$��#	�GCپ�ɢ�$�d�1��+���MB�����T(��P��\��C��';2)���T��>��Ѳ��ٿ��������TC$�(�&���#�����������׿�ձ�V���rWT���1[;����43�S���.�z*
�@�J��7��U�yh�=��\2ܾ��
���&��/?�TiR��^��   �   Ӂ�G,�Y������`ھ�ϲ�^V��h�G��,��ꚽ���A������RX2�oǽbr>�>r�������;�(����z���ֿ���*����+�RW<��G� �J�\~F�|Y;���*�����7���տu<��x���=k;�O  ������@���˽;��M��(쥼8�%�/��f���L���o��@ݾ� �7��?���   �   ��þ�
���G��������	[U��n��^ѽ��k��¼���̺ �z;h+�H�H�ơ�g��þ���\\��j���ƿ�a��<^���0��hI�$H^�0Gl��q�R�k�~Z]�\{H���/���7D���Rƿo◿�p]����v
ž��j������T� W��Ǖ:Ў�@pռ�ly���ؽw!�&�Y�P���z�������ȿ��   �   ��h��Mb�
�P�(�5��
�H�ܽ^����l���8y<�<�<�͚<�YŻ�Bd���f����T�a�,�v�y�����9޿����(�ַG�t�e���^������X����~�.e�&{G�* )��q��߿���T{�|.�
�JB������q��g���<���<hkH<HJ�z���ܖ��㽖L��8���R��oc��   �   ]� �$n����߽�����ŉ���(���q�><��<t�'=\O,=���<Ph��@G~�
��SҔ�����&�=��G��@a���������7�� [�X�}�����y������Y������B�}��T[���8�n��oy�ܺ�����[�?�����ŉ���3"�ٿ�� ��Dk�<�3 =��=4V�<�\�;�Y���4��?���;�����C���   �   b����Յ�:We��*�����`�̊<¦=2�I=^�d=dMU=\= zW�*C��&�(��s���>�"pH�����g�¿�������
�A�Z�g��!��ٗ��;���=���6��s��sZ��r�h��B�X�������Ŀe��G�J��%��v����-�&f���nݻ���<I=P�X=��==�=@�g<�ǻȿԼʾ2��Wk�p���   �   ��N�B�A�L*���Ӽ8�� p<�$�<�2=@Sd=Ԕx=2�b=g=`WM������,�Fʡ�����!L����ƿv ��'!�BSE���l�����I��H���)��>��Uk��}Z��΍m���F�Rp"����p
ȿ����(�N�G���社��1�8ؓ�@?ڻHN=JV=,�l=<�X=Pu'=���<���;��@�Hj�4�$�VE��   �   t����Յ�TWe�2�*�0����`�̊<�=x�I=ҽd=$NU=R]=`[W��A����(��r���=�0oH�������¿������*�A�2�g�� ��.ؗ��:���<���5������Y��B�h�*�B��������
�Ŀ���P�J�2%��u��z�-��d���^ݻt��<�I=��X=�==8�=��g<PǻԿԼ־2��Wk�p���   �   n� �Dn����߽ٕ��
Ɖ���(���q� ?< ��<H�'=�P,=`��<�J��|A~�ɸ��Д����Z�=��F���_��������8�7���Z���}���x����X��	�����}��R[�0�8� ��aw�zں�]�����?���������1"�޼��0z�Lp�<P5 =��=tW�<�_�;@Y����4��?���;�����C���   �   ��h��Mb�"�P�<�5��
�R�ܽS����l�켻�y<�@�<0Ԛ<�0Ż�:d������tQ���,��y�����v޿����(��G�
�e��� ��������U����~��*e�VxG���(�p�%߿u}���{{��y.�z��?�����@�q�hR���<8��<�pH<�F�����ܖ���㽘L��8���R��oc��   �   ��þ�
���G��+������[U��n�~^ѽB�k� �����̺��z;��*���H�]���f�xþ���X\��g��+ƿ�]���[���0�@eI��C^�fBl���p���k�$V]��wH���/�.�
@���Oƿ�ߗ��l]����8žހj�����T�hW��K�: ���mռ�ky�\�ؽ�v!��Y�R���z�������ȿ��   �   ہ�P,�b������`ھ�ϲ�`V��X�G��,� ꚽ���8��L����M2�fǽJl>��m������P�:�@���1w����ֿ�������+�S<�G�B�J��yF�BU;���*�j���4�_�տ�8�������f;����������@���˽Ft;��?��㥼d}%�3.��"���L���o��Bݾ� �=��F���   �   �pb���]�K&Q���=�V�$��#	�LCپ�ɢ���d��0�]*���IB����8J(��H��=������;�$���T�';���̲�<ٿ.��������?$���&�R�#���T�[�����׿�б�����|QT�m	��T;0���-��J��>�.�x#
���J�Q6���T��xh��<��P2ܾ��
���&��/?�[iR���^��   �   ����������7����-j��D��J��"�]��M�m����7���h�R�x0�h||�"{གྷ�B����0h쾮^'��j`�K:���خ�^�̿�N�;���j��|����Z`�����g:˿�k���*����^�ˁ&�;~�j�����B�B;� +���3��lW��+�����3�p�@0�������
 �T�F��ml�����aw�����   �   �Tҿ�cοǝÿ�����ҝ�ԅ�^�Y���(����Vꬾ�Xa�>�������L��bM�r���t�	���b��7������3*��[�����;��r^����ĿXϿdQҿ~`οl�ÿ�����ϝ��х�0�Y�?�(�̜��j款bSa����`�����L�ldM�������	�p�b��;������6*���[���}>��a��C�Ŀ�Ͽ�   �   �~����d��#��|=˿Ln���,���_�Ą&���뾗�����B�j@��/�`�3�hW��&�����5�p�$,��0���" �:�F�il�����zt��|������ ������z����(j���D�G�)������m���򯽐�R�v 0�|��	�B�L��l�Xa'�dn`�m<��.ۮ�Q�̿R������k��   �    �&�t�#���(�����a�׿Vӱ������TT���X;�����/��M��b�.�  
�ʜJ��/���O�#rh��8���,ܾ5�
���&�+?��dR��^��kb���]�b!Q�&�=�E�$�B 	�v=پŢ��~d�n+��"��@B����vI(��J��t������;�&�c�T��<���β��ٿ@���H����4A$��   �   ��J�|F�jW;���*���N6���տ�:�����+i;�����Y�����@��˽dv;�(<��tץ�>s%��&������L�5����i���ܾ �o��A���}�G(����y���ZZھ!ʲ��Q���G��&��ᚽ`��*��D���N2��ǽ�n>��o��g���U�:������x����ֿ<�������+�(U<�bG��   �   :q���k�^X]��yH�`�/���EB��aQƿ4ᗿ�n]�?���žփj�j����T�X�V��˖:����Vռh\y�<�ؽ�p!�f�Y�����u��񟳾�¿���þ����A��󦞾���SU�Ah��Sѽ��k�H��� �˺ ?{;X�*�l�H�r��!g�5þY���Z\�.i���ƿ�_���\���0�gI��E^��Dl��   �   蚋��V����~�f,e��yG�$�(�q��߿�~���}{� {.���5A��~���q��R���<T��< �H<�����Ӗ�T��`F��8�N�R��gc���h��Eb�]�P��5�f�V�ܽ!����]�P����+y<�L�<�ۚ<�$Ż�;d��������R���,���y�{����޿����(�b�G���e���;����   �   ����X��������}��S[� �8�ޮ��x�oۺ������?���������2"�$��� ~��r�<\8 =��=�d�<`��;LC����4��7��E3��Q��9��X� �8d���߽������6�(�(�q� e<��<��'=�T,=x��<@B���A~�Y��,є�����	�=�AG��Q`�����b����7�~�Z���}�����x���   �   =��6����Z����h���B���������Ŀ2���J��%�pv��Z�-�~e��0dݻ���<,I=��X=�==R�=(h<��ƻ\�Լ��2��Nk�]k������-х�8Ne��}*����@v`�|׊<��=>�I=��d=NPU=�^=`MW��A���(��r��>�soH�,�����¿���P����A���g�<!���ؗ�U;���   �   *�����������q���Q�j1����E鿱���X�4|7���s	�����2�]�`}�;�(=N�q=)�=rt=z(G=^
=0:�< M:�X`�pf̼����������Ȼ���1�0��;���<0�=��Y=�y�=�ʌ=�Ă=�><=8z,<��F�}��1��]`�!�4�$*���s�����V��h�/�.�P�*@q��Ɔ�X~���   �   櫐�R��=�����l�L�M�^�-�Nh��^忁��������4�*A꾝싾ze�Z;W�`�;��!=�e=�1t=v[=�'=$��<�~�;(�F��0漆	&�v�E��O��)A�R{�XUμx]���"<,|�<RC:=�in=Q��=�Ly=x�5=P�)<ָ@����5�����VD1�&��M���[ �?�n�,���L���l�����W���   �   r��3[���w�T_�B�B��%��T��ڿ/����pu��)��Zܾ	������E��K�;b =��@=>�<=�8=��<�8����T��۔�3�[�ʽ��н�ȽeA��T`��PE�H�Ǽ �e��^�<�C#=.�O=��S=�V!=��<��0�M;��3�Wbؾ՚'��r������\ؿ���t$�H9B��_���w��y���   �   (�s��|n���_��J���1����!����dȿ���	�_�/Q�r�ƾQj����`O,� �U;�&�<�X�<���<@![;�<���c��鶽O}��l>�&�2��}A��F�	@�.0�������R���JO��ә���<<2�<��=�3�<��;�r�%���d�W�þ�}���]��}��(kǿ���Lq��2�(;K��`���n��   �   �T�|P�*%D�2����$���,߿�䱿����c�D����/��� H���Ƚ�� �ɹ��M<P��;H H��3�B3������9�7j�����?%��G���0_�����t��0�����d���3�F��������И��X/@<���<`�f;������ğC�-e���J�jyC�)������N߿�$��9���3��E�T�P��   �   �4���0��_'������E�h�DK��r�f���%����X���X"�����x��� '� �߻��ͼ>Au�7�޽0�,���r�Ꝿ�����#�$���X��.G�74�6����C޾IG��:���8jl��B'���Խ�kc��1��@�X��,��x�ۼ����P�d+���V߾�d%���f����������j��N/�^(�r�1��   �   ���Z���@��I���6�7t��4%���z�:D<�������3�]��K��4�u��Nݼ�0���;�:����P���ZF�8P������Ty��kI��w)�X�:�e�E�e*I�1�D�%\9��'�D@��}�-���6���.A�t�񽹃���������'˼�n������\�"���5�8�<�h|�{9��pÿK5俦� �
/��p��   �   N��rW��#ο�9�� ��h}���E������;���]�#�^_����6�%�V4�v_�������wM����+�־�^�I�0�SrR�GGp����x ���M��sx���ǂ��m���O��%.�dL�ԚӾPc��k�I���/݅�U���ڼ 3�ၲ���#�蜇�@
ϾH���uG����ì�����пb��M>��   �   ׼��3���Y��[)��猿W3n���@�,��T�پ�����>��޽$�m�hJ��4	�йp��:ὴA�5���ܾ_��+C�	q��}��1�������빿Vڼ��6���\��,���錿�7n�$�@�����پ6����>�ʒ޽L�m��K��1	�:�p�.4ύ�@��1���ܾL}�]C��q� {��R��������繿�   �   �J���u���Ă�H�m�P�O�J".�WI���Ӿ�_�� �I����|؅�bP���ڼ>3�g���Y�#�����;Ͼ����xG� ��;���S���	п����A�����Z���&ο1<��o�� l}���E�:��'�;E����#�c��f�6��!�X.�Z������rM������־�[�a�0��mR�DBp�b��������   �   �%I���D��W9��'��<��w�(���2���(A����}��@p�� {��,)˼�n�����4�\�0���V��<� |��;��
ÿ;8�L� ��0��r����2���B��L���9⿛v��6'��X�z��F<����������]��O���v��Mݼ (���2�{���G��*TF��K�������r���E�cs)���:���E��   �   }C��0�c����=޾�A�������bl��<'�3yԽP^c� ���jX�����ۼ��S��-���Y߾�f%�|�f�e���0���v�����0��_(�l�1���4���0�da'�R�D��?H�\����L���f�i�%�������Z"�����0���0�0x߻t�ͼ@2u��޽��,�f�r�$坾�{��3�(�������   �   �Y������o��������d�}3�����������F���J@<���<`�f;�����`�C�4g��XL�m{C�]*�������P߿&��:�Z�3�zE�V�P��T�tP��&D�L�2� ��8��a.߿h汿�����D�҄�˼��
H���Ƚ�� �ȹ��M<���;��G�3��)���{�|�8��.j���� �����   �   h
F��@�H�/�D}�g�� I���:O�X��� �<p@�<��=�8�<� �;*u�ڢ�:�d��þ�~�@�]��~���lǿ���Rr� 2��<K���`���n��s��~n���_���J� �1�t������fȿ����i�_�)R���ƾ�Rj����8P,���U;�-�<�c�<�и<��[;0!�� c��߶��q���7��2��vA��   �   ��н{Ƚ�8��X��HBE���Ǽ �[��n�<�I#=��O=��S=�W!=p�<�0�h<��5��cؾϛ'�:�r������]ؿ���ju$�<:B��_�R�w��z���r���[��0�w�`_��B��%�U��ڿ͐���qu���)��[ܾ�������E�`S�;�"=>�@=x�<=|?=D��< ������J�T��Ӕ�z鵽>�ʽ�   �   ��N�2!A�Hs��FμPC�x�"<���<G:=�ln=I��=�My=ҽ5=��)<z�@���N6��w���D1����υ��� �n?���,�4�L�2�l���hX��O���eR��������l���M���-��h�'_�����ҕ��;4�yA��싾�e�2;W���;��!=�e=j4t=�y[=:�'=���<@��;ȍF�!�"&���E��   �   ������ɻ��1��;��<�=<�Y=�y�=hʌ=�Ă=D><=�w,<��F�i}�$2���`�S�4�B*���s��
��j��~�/�H�P�@@q��Ɔ�\~��*�����������q�p�Q�T1�����D鿍���9�|7�s�:	�����F�]� ��;(=��q=M)�=�t=�(G=�
=�:�< M: X`�Hf̼����   �   ��N�F!A�bs��Fμ�C�`�"<���<G:=�ln=���=~Ny=�5=��)<��@���5��E��D1������� ��>�&�,�@�L��l�Y���W��|����Q������L�l���M���-��g�-^�����:���Z4�=@��닾�d�H8W����;>�!=��e=�4t=�y[=t�'=���<��;��F�0!�.&�ФE��   �   ��н�Ƚ�8���X��\BE���Ǽ �[�$o�<DJ#=j�O=�S=�Y!=��<�~0�^:��2�raؾ0�'��r�X���\ؿ���t$�|8B��_���w�9y��Zq��uZ����w�$_�B�B�%��S��ڿS����ou��)�jYܾ��� �E�@p�;%=ȫ@=v�<="@=��< ������:�T��Ӕ��鵽O�ʽ�   �   y
F��@�\�/�U}�|��'I���:O�й����<�B�<P�=|>�<PF�;�m�6����d���þ�|�0�]��|��jǿ���lp��2��9K�f�`��n�B�s�{n�4�_���J���1����g���pcȿ튙�C�_��O���ƾ<Nj���H,��V;(4�<,h�<�Ӹ<`�[; ����b��߶��q���7�$�2��vA��   �   �Y������o��������d� }3�������4���<��hS@<�<`g;`��}��I�C�qc���I��wC��'������"M߿�#�P8�0�3��E�`�P��T�zP�N#D��2�H������*߿O㱿E���T�D���󸫾��G���Ƚ�� �Ź��M< ��;h�G���3�0)��n{�h�8��.j�
���& �����   �   �C��0�s����=޾�A�������bl��<'��xԽ�\c�P��@-X��솻�}ۼ����N�r)���S߾�b%�6�f������������-�T\(���1��}4���0��]'��l��aC�B�{I����f�[�%���������T"�{���H������0V߻��ͼj0u���޽r�,�D�r�坾�{��6�1�������   �   �%I���D��W9�
�'��<��w�(���2���(A���|���h���n���˼��m�����
�\�Z���L���<�*	|�}7��ÿ�2�� �R-��n�ؽ�~��?�?F��4⿩q��#��|�z�^A<������s�]��D����u��9ݼ����.����/F���SF��K�������r���E�es)���:���E��   �   �J���u���Ă�S�m�W�O�O".�ZI���Ӿ�_����I�����օ�vJ���ڼ3��{����#�6����Ͼ���grG�
��o������}п���:�����S�T� ο�6������c}�7�E���z�;����~#�dX����6����'��W��.����qM�������־�[�\�0��mR�GBp�e��������   �   $׼��3���Y��a)��!猿^3n���@�.��J�پ凕�.�>�u�޽��m��A��'	���p��,���@�7.����۾mz��C�;q��x�����������乿�Ӽ�a0���V���&���䌿�.n���@�����پ[���&�>�Ƅ޽��m��>��(	�r�p�O2�"�@�`1���ܾD}�VC�q� {��V��������繿�   �   S��yW��#ο�9��#��#h}���E����~�;�����#�]��Z�6�h弎#�bS������:lM�A�����־�X���0�|iR�j=p���������H���r��R�]�m���O�p.�F�Ӿ�[���{I����х�2D���ڼt	3�^��Ǫ#�����
Ͼ;���uG������������пe��Q>��   �   ���^���@��I���6�;t��8%���z�:D<�����󲾨�]��I���u��;ݼ���l'�&���o=���MF��G�������l��&B�_o)���:�"�E�!I���D�aS9��'�9��q�b#���.��J"A�e��u���V��he��X˼,�m�����q�\�򩲾&�1�<�b|�z9��oÿJ5俨� �/��p��   �   �4���0��_'������E�m�FK��u�f���%�ޟ�$���GW"�����<���p��+߻��ͼ�"u�&�޽L�,���r�`���Yv����S������?� -�����;7޾%<������jZl�@6'��nԽ�Mc�,�� �W��҆�$~ۼ}��� P�$+��~V߾�d%���f�����
�����j��N/�^(�t�1��   �   �T�~P�,%D�Ĕ2����&���,߿�䱿����b�D����
�����G���Ƚ� NŹP�M<`�;��G��s3� ���u�w�8�l&j�l����릾^T�����j������Q�d��u3��� �צ��.�������r@<�̇<�'g;�����*�C��d���J�cyC�)������N߿�$��9���3��E�V�P��   �   *�s��|n���_��J� �1����%����dȿ����_�+Q�^�ƾ�Pj����(K,� V;�8�<<q�<��<�w\;�����b��ն�of���1�>�2�WoA�F���?�^�/��v����9?���)O������&<�R�<��=�E�<�Q�;�n�Ǟ佀�d�8�þ�}���]��}��(kǿ���Lq��2�(;K��`���n��   �   r��4[���w�T_�B�B��%��T��ڿ1����pu��)��Zܾ��,�t�E��l�;@&=��@=ڸ<=JF=0��<�G���k�T�T��˔��ൽR�ʽ��н�ȽO0���P��4E���Ǽ <Q�x��<Q#=��O=��S=B\!=�<�~0��:��3�EbؾК'��r������\ؿ���t$�H9B��_���w��y���   �   櫐�R��=�����l�L�M�^�-�Nh��^忂��������4�%A꾐싾Le�:W�0�;r�!= �e=�6t=�|[=0�'=<��<���;�sF�H��%�R�E��N��A�k�P7μ�'���"<��<vK:=Ppn=ִ�=xPy=F�5= �)<~�@����5�����SD1�$��M���[ �?�n�,���L���l�����W���   �   ��v���q�l�b��;M���3��:�'~��ďʿ�>��4�b�����Ⱦd�j��[�,��\͛<n}N=	Ň=M��=D��=$�i=b4=���<�z<@-2;��XTS�`Gl���:��A�����;���<T�=r2P=�ۃ="4�=v��=���=�n=`��< zϼZ�ֽ��a���þ��_�2:��=Xȿk<��R5�3���L�T�b�Цq��   �   ��q�$�l�Nf^��cI�@�0�(���A���!ǿn����^^�U���ľoe����\�@v�<�I=�x�=3È=j�{=�)N=�O=T�<��;��"�Di��\߼\�ĩҼH]�������<�8�<�!.=��k=�F�=�q�=�*�=9h=�f�<�ż��н��\�����5�[�Ĥ���ſ�<��^���0�nI��Y^�.�l��   �   l�c���^�b�Q�r�>���'�&&�9�쿒+��0���KR��G�M�����U���ν0b伸��<� 8=�]d=��`=4l9=�g�<��&<�l/��t����H�8��.���b����]��(su�P7�H;Ҽ���L�<:�=��W=�/=cM�=��U=�Q�<p����Ͽ�F�M������O�[�����5��Р��Z'��>�`
R��)_��   �   �N�&�J�@)?��4.������f�ٿ����>���n?����6�����=�s(��H���T��<�"=�r+=�=�Z�< 9һ���ɂ�5�������:��Pv�����	�M��߱�4)k� h� #>:�9�<�.)=��G=Χ4=��<HƂ�u��h�6��$��5� �j=�t<��O����Lٿ��&���.���?���J��   �   R$6���2�f�(�w�r��2N����������h��~'�6�⾦������������H2k<�F�<�M�< ^s;�|ż��t�~ν ���=�2�c�����<鉾����݈��L}��,^��A7�����|����W�t���0�)<�5�<��=� �<@t3����V��|���
�}J&�)�g��s���������^[	��A�v�)��3��   �   ��`�<�@��Ũ�A�ɿ���B���<E�#��p黾��g��?����\���9�0�<(�<j�T���^��t��+E��[���;��B���l"Ҿġ߾��#\޾D�Ͼzr��������|�n=��!�����bd� g�`�c<`�U<�^�phL�6���/id�����O+E�M]��q̦�`�ʿ+V���
�����   �   �Q��U�8�ݿ$RĿ�h������V�) �cCᾌ���2�0�����(c� }ֺ�pj��\8��&��Fu��Hk�/���M�;G�����)���m(�cg+�V�'�v�[��3���ɾ�s����c����Ʊ��$��R&��'�:����9�����0��֓���ᾅ� �XX��&��}㨿�&ƿ��߿"��" ��   �   9/ҿ>(ο�Nÿ����uz������~Y�?N(�l���1_��D�[�=&����z�Z¼�����5��7���i$��}�0ҳ�����ݭ3���M�(b�F�n���r�X�m�D`��_K�H1�3���D����sqw�lu��T��П(���e� ���43���y�����]��������1�)�ld[�Z���:��`��+�Ŀ��ο�   �   �g���+���p�� ��C�q�ҟK���#�����@T��Ǉt�B��aw����8^�0yc��3�w��2F���x��������=&�d}N�u�������� נ��j��a.��[s��{���r���K���#�����X��X�t�&��j|�� �  ^�Xoc�<-�����A��x���������:&�lyN�vu��}��ޠ��MԠ��   �   ��r�w�m�k?`��[K��1����b?꾝 ���jw��p�cN��p�(���e�����@:���y�q���~]��������. *�h[����A=���b��"�Ŀ�οS2ҿF+ο�QÿS����|��ɇ���Y� Q(�����Nb����[��+��� {��^¼���X���5�p0��cd$��}��ͳ����3���M�W#b�U�n��   �   Cc+�M�'�0r��������ɾ�o����c�l��f���B�$��8&�@��:����r=�]�J�0�Eٓ�7���� �~X�o(���娿)ƿ��߿;��R$ ���3T��S���ݿ�TĿ�j�������V�d ��F�� ��� 2����Ԭ��a��ֺ@Rj��P8�5���o�zAk�����;���%��@��ti(��   �   ����U޾V�Ͼm��������|�^g=�{�����VX� ]� �c<P�U<�j�jmL������ld�̍�����-E��^��UΦ���ʿ�X���������,��������+��P�ɿ�������>E�ƈ��뻾Ʒg�OC��X�\��9��<p�<p �4��V���y��$E�7W���6������ZҾg�߾�   �   P���Xو��C}��$^��:7�����r����W�Ȉ���*<�A�<f�=0"�<�{3��8Y��~��t�@L&�v�g�pu��v�����꿎\	��B���)�\3��%6�H�2���(�Rx����P꿁���ѵ����h�b�'�P����W��M�����h9k<HO�<T[�< �s;@bż��t��ν���S�=���c�����䉾�   �   �o������	�M��"ֱ�lk�@Lༀ�@:K�<�4)=0�G=
�4= �<hʂ����k�6�n&��Q� ��k=�o=������,Nٿ��.�ȭ.�V�?���J�~�N���J��*?��5.����l����ٿ�����>�� p?�Ι�Z����=��)���������<�%=~w+=�=Xm�<p�ѻ�r�=�����������δ��   �   R����U��6du��7��"ҼPǒ��]�<H�=�W=�3=�N�=��U=0Q�<(����ѿ���M�M �����F�O���	���M��x��r['�Ԏ>�lR��*_���c���^�Z�Q�F�>�B�'��&� �E,�������KR�~H������U���ν$c�X��<�8=4ad=��`=Fr9=Tw�<�'<0@/�[����H�����9����   �   �L��ҼO���x�� �<�B�<&.=2�k=�G�=�r�=0+�=d9h=�e�< �ż��нȦ\�Ӯ��6��[�5���ſI=�����j0��I��Z^���l�n�q���l��f^�`dI���0�h��`B��3"ǿ�����^^���D�ľ\oe����@��w�<�I=�y�=^Ĉ=j�{=�-N=lT=H�<p=�; �"��Z��߼�   �   HGl���:�pB�����;L��<&�=<2P=�ۃ= 4�=T��=]��=tn=(��<�{ϼ�ֽ�a��þ�I_�P:��_Xȿ�<��b5� 3���L�`�b�Ԧq���v���q�^�b��;M���3��:�~����ʿ�>����b�~���Ⱦ��j�,[�V���Λ<�}N=5Ň=y��=i��=n�i=Lb4=L��< �z<@/2;���SS��   �   �L�ؚҼ@O���x���<�B�<&.=R�k=�G�=�r�=~+�=r:h=�h�<�ż��н_�\�ɭ��O5��[�����BſF<�� ���0�I�pY^���l�,�q���l��e^�hcI�ȯ0� �OA��V!ǿ�����]^���0�ľ�me��ས� {�<I=z�=�Ĉ=ֲ{=�-N=�T=��< >�;�"��Z��8߼�   �   `����U��bdu��7�#Ҽ`ǒ��]�<x�=��W=r4=BO�=��U=4W�<�*ο�+�M�O��y��W�O����u���_��L��Z'��>�n	R��(_�F�c���^�P�Q��>�Ɨ'�v%��쿠*��k����IR�G�������U��ν8Y��<�8=�bd=��`=s9=Px�<h'< ?/��Z����H�����A����   �   �o������	�h��2ֱ�xk�LༀA:(L�<�5)=��G=��4=�
�<t��������6��#��[� ��h=��;��U���|KٿH��>���.���?��J���N���J��'?��3.���������ٿV���=��;m?�ɗ�����6�=��$����̶�<�(=�y+=` =Lo�<��ѻ\r�������������ִ��   �   Z���dو��C}��$^��:7�����r��p�W�����*<�E�<��=X,�<�\3�%�T�s{����I&�9�g��r��4�����HZ	�L@��)�.
3��"6��2���(��u�@��L�-��������h�}'���⾴�����'��������Ok<�V�<``�<`t;�_ż��t��ν���H�=���c�!����䉾�   �   ����U޾c�Ͼm������|�[g=�h�.���W����c<��U<@&�v`L�-����ed�����v�&)E��[���ʦ�W�ʿ�S�H�����l�����������9���ɿ�����:E�:���滾��g�i9���z\���9�(�<��<�
�P��rU���y��$E�(W��}6������^Ҿo�߾�   �   Kc+�T�'�8r��������ɾ�o����c�F��˽���$�0*&�  ;`c��T0��趽(�0�0ԓ�*��L� �}X��$��bᨿ$ƿ;�߿$��! �~��M��C�_�ݿ�OĿ�f������V�� ��?ᾶ��d2����F��=��<պ�Aj�@N8�J��Lo�BAk�������;���$��C��zi(��   �   �r���m�t?`��[K��1����f?꾘 ���jw�hp�iM���(�p�e�@���� ���y�����]�f�������o�)��`[�L	��e8��_]��K�Ŀ��ο$,ҿ3%ο Lÿ�����w�������Y�AK(������[����[�=����z��D¼`��x	���5�/���c$���}��ͳ�����3���M�[#b�Z�n��   �   �g���+���p�� ��L�q�ڟK���#�����4T����t�Ԁ��u������]��Jc��"�/���=��yx��������a7&��uN�u�{��8����Ѡ�e���(��n��������q��K�O�#�����P��b�t�o|�p����P�]��Nc��'����KA�vx�l��~���{:&�hyN�uu��}��᠘�PԠ��   �   =/ҿD(ο�Nÿ����yz�����Y�AN(�c���_����[��$����z��L¼p������ 5��(��J_$�=�}�Sɳ����U	��3�B�M��b�x�n��r���m��:`�?WK��1����9�����cw�8k� F��R�(�Pre�`}��%��
y�]���]�s�������'�)�dd[�W���:��`��-�Ŀ��ο�   �    �Q��[�=�ݿ(RĿ�h������V�) �VC�j��2�w����A���Ժ�(j��C8����j�b:k�)���k~;������o��oe(�*_+�D�'�Xn�R������\ɾ�j��W�c����d���*�$��
&� ^ ;�]�� 3�춽�0�o֓�c��z� �QX��&��{㨿�&ƿ��߿&��" ��   �   ��b�@�D��˨�D�ɿ��C���<E� ��Y黾R�g�?>��N�\� �9���<�<���xt�FM��.t��E�S���1��3���fҾ"�߾?�㾏O޾X�Ͼ�g���|��b�|�O`=���X����I������c<8�U<@&绶cL������hd�����
�H+E�J]��n̦�^�ʿ+V���
��
���   �   T$6���2�j�(�
w�t��6N�����������h��~'�(�⾆����ޥ������Qk<�\�<l�<��t;�Gż�t��ν���0�=��c������߉������Ԉ�;}��^�j37�T��zh��|�W�m���A*<�S�<�=L0�<�^3��dV��|���
�vJ&�$�g��s���������^[	��A�v�)��3��   �   �N�&�J�@)?��4.������i�ٿ����>���n?���!���N�=�E'���������<�*=�}+=�&=x��<pzѻ~d�����.��������~��fi�a����	�&��"̱�k��.� �C:_�<=)=��G=֯4=@�<����.���6��$��,� �j=�r<��P����Lٿ��&���.���?���J��   �   l�c���^�b�Q�r�>���'�&&�9�쿓+��1���KR��G�A�����U��νX]����<�8= ed=z�`=fx9=D��<@;'<x/�xB����H� ���c���`����M��@Uu���6��	Ҽ@o��Hp�<(�=��W=9=�P�=��U=Y�<p塚Ͽ��M������O�Z�����5��Р��Z'��>�b
R��)_��   �   ��q�&�l�Nf^��cI�@�0�(���A���!ǿo����^^�U���ľ�ne�b��6��y�<RI=�z�=|ň=R�{=81N=�X=X%�<Pl�;�"�XL��H ߼t=��Ҽ�@�� C��X�<PM�<�*.= �k=zI�=t�=\,�=�;h=0j�<��ż�н��\�����5�[�¤���ſ�<��^���0�nI��Y^�.�l��   �   ��I�Z�E�<�:��6*��S�ʦ �K�Կ�h��'耿@W:������O��5�J�� B�6!=�	q=�	�=m��=fȔ=N=�=\�[=��*=hV�</�<@[B<���;�#�;`%<�p�<��<v =�R=Lʄ=Z.�=X�=i�=v��=�^�=v�5= #˹���0�)����������7��K~�n���aӿ���������)� �:�$�E��   �   ��E�
B��K7�|@'�������FHѿ�y��t*}�Y�6������ǜ��g0�B����-��C=h�l=ӡ�=���=k��=��p=��>=�E=p �<8�< 2\9@7���2û��3�0ȓ; �x<���<�(0=�4l=�#�=��=O�=֩=j��=R�4=��:�����%��Q�����3���y�fˤ���Ͽm���xV�^'�G7��B��   �   P;�L�7�~�-����v����ƿ��2�o�>�,��������#�[͌��i���=.�^=%�=
R�=r _=��(=@�<�r�;����'Ǽ$R�dv.�>$5��{%�0� �Ե��@2����<jF=ڪX=4��=)��=�=˃�=n�1=��[;�	q��K����h��)�)�� m�������ſ����K����d�-���7��   �   �w+�.<(�nO�(��K+��7ݿꗶ������Z����o�ҾC�����J�i��x��� =��E=�T=�a9=d*�<��/<x�Q�z��<�{��+����ʽ�$߽l��$�ڽͦ��6��
[���������<�$-=,�h=W�=�q=�#*=0x�;rTF��7��a}���ξ%����X��ڏ����_ݿ�X�"1�8��2�(��   �   �-�ZW����H��6���Ŀ6ա��-��?�fW�J�����]����(�/��TX;�a�<zI=��=}�<@O������Ҍ�I}ֽ���l.�m�F��AV�g�Z���S�rGB�t�'�b���tý~_p���ü���;���< �6=��D=XP=��7<ڥ���ܽg�W�x鲾�.�d�>���~���o.ſ���@[��&�����   �   R�S� �8���߿m�ſk����3��ލX�qf!��(㾛���� 1�Z���Ȧ伈V<��<Ĵ�<�6.<`�}�0,T�'�Ľ\t�O�J�h;~������᧾0���w��<���VJ���b����u�jA��k��ϰ�t�,� �λ@~�<�+=�e=hhh<����in��rX-�����I�aZ!��Y��Ί�շ��C/ǿ��%D��~��   �   )�ڿ��ֿ�S˿e	��5#��<R����b��30�����$��#�f�Q���r�h�_��/< f�<`�;�B���z��B齥B5��X}��F����Ⱦ��9��)	�����_��w���tľ�O���xs��+��׽��Z��qc�ع=<��<@$w<�'�p�g���&\f�R���؎��f1��d�����ϫ��ӝ���̿�Q׿�   �   }��3����G���4ς�ԡ\�2����8�ƾC����U&�l����8���ʺ��,<`ԋ;x����hx�^W�LD�e���v��*������(�:���D��3H�i�C��E8��}&�)�j�-8���E��^�<��R���b��y� d�;�pU< x9�R�쭱���'�R@��Bɾ�
��I4��b_�qW��>r���|���B���   �   �쇿�%�� R{�%Nd�FG���&�V���Iɾ玾Ƨ:�0׽�D��r/����;@��;h�G��N��޽��?�����D;g�Re)��&J���f��l}�����(���V{�KRd��IG�̪&����MɾIꎾ|�:��6׽��D���/����;��;X�G���N�Hx޽g�?�-��@@;?d��a)��"J�;�f��g}������   �   s/H�F�C��A8�Iz&��%��d3��CB���<��J彦vb��y� ��;�rU< E���d����(�4C��% ɾx�
��L4�af_��Y���t��'��rE��$
��̘��/J��`���8т�Q�\�2�����ƾ����jY&�O���@>� '˺ �,<���;�����\x��N�FD��������r��6��G�(�:���D��   �   +��R\�fq��#�Dľ`K��yqs�C�+��׽�zZ�HMc���=<4��<�"w<h '�εg�� ��`f�l�����/i1�T�d��������F�����̿�T׿�ڿn�ֿ.V˿���L%��T����b�(60����['���f����r���_��/<|l�< ��;0/���xz�69�~<5��P}�6B��K�Ⱦ���5�y&	��   �   ,r������WE��^����u��A� f��ư�l�,�p�λ���<�/=xg=�ch<���Dr���[-�G���M�x\!��Y�PЊ�����o1ǿ/��F�������� ����P�߿x�ſ.���/5��A�X�Mh!��+㾌���<#1����� ���T<X��<X��<�U.<(�}�\T���Ľfn�$�J�3~������ܧ�����   �   w�Z��S�@B���'�n��Sjý�Np��mü�;�;P��<p�6=��D=Q=��7<����ܽP�W��벾,0�Y�>��~�b���/0ſ���`\��'�γ�/��X�ғ�X���忪�Ŀ�֡�(0�ϸ?��X�����]�y�4�/��HX;�d�<M=D�=̍�< ���T��ʌ��rֽ����e.���F��9V��   �   z��j�ڽ�����,���	[����`��<J,-=��h=�X�=ڼq=$*=�j�;bXF��9�Od}�u�ξk��^�X��ۏ����� ݿ�Y�2�F��R�(��x+�F=(�rP���,�59ݿ ���o���O�Z����߼Ҿ9���%����i������ =*�E=6�T=�g9=H:�<H�/<pPQ�����{�"��J�ʽ�߽�   �   �5��n%��� �\����涺��<�M=�X=���=⤙=3	�=P��=0�1=��[;q�BM�������%�)��m�a�����ſ��ￒL����2�-���7��P;��7�>�-���� w�����ƿ���o��,�������#�1Ό��m黊�=��^=�=�S�=�%_=��(=H"�<P��;X���Ǽ4E��h.��   �    �»�(3����;`y<p��<-0=f8l=%�=4��=�O�=�֩=���=�4=�g:Ԟ��ǩ%�AR����򾣹3���y��ˤ�7�Ͽ����V��'��G7�pB�l�E�r
B�BL7��@'���%���Hѿ�y���*}���6�ޢ��Ȝ�h0�y�����-�D=l�l=���=��=���=��p=��>=jJ=�*�<��< xb9 ���   �   0$�;X%<�p�<���<T =��R=8ʄ=H.�=:�=�h�=R��=_^�=�5= �˹������)�.�������*7�L~������ӿ���������)�*�:�(�E���I�R�E�2�:��6*�|S��� �-�Կbh��耿W:�=���[O���5����HB��!=*
q=
�=���=�Ȕ=p=�=��[=��*=�V�<\/�<�[B<���;�   �   @�»�)3�p��;Py<p��<-0=~8l=%�=S��=P�=�֩=��=L�4=��:9�����%�`Q�����ȸ3�|�y�)ˤ�[�Ͽ���8V�'��F7��B�|�E��	B�jK7�@'�b�����Gѿy���)}���6�����*ǜ��f0�Ċ����-��E=��l=���=��=�=$�p=
�>=�J=D+�<��< �b9����   �   �5��n%��� ����� 綺��<N=$�X=ɐ�=:��=�	�=-��=֑1=��[;�q��J�Y���u�侁�)���l����9�ſ���hK�@����-���7�,O;�p�7���-�R���u���	�ƿ ��o�;�,������%#��ʌ��I黔�=��^=E�=�T�=p&_=��(=H#�<���;0��|Ǽ&E��h.��   �   ���w�ڽ�����,���	[�d�漠���<�,-=��h=�Y�=4�q=�'*=���;�OF�r6��_}�$�ξ%��`�X��ُ�{��ݿ0X�B0�:���(�fv+�;(�^N�.��m*�a6ݿ����z���7�Z�T��t�Ҿӱ��֎���i�`"��� =,�E=Z�T=6i9=�<�<Ь/<�MQ�����{��!��>�ʽ�߽�   �   ~�Z� �S�)@B�ɱ'�x��YjýrNp�mü�@�;���<2�6=|�D=�U=��7<ޟ���ܽ̏W��精s-���>���~����,ſ��4Z�~%�D���,�V�l��&��/��J�Ŀ�ӡ�y+��?��U����Y�]����n�/�@�X;�n�<�P=о=|��<�ꆻD���Ɍ�Wrֽ����e.���F��9V��   �   1r������aE��^����u��A��e��ư���,��}λl��<�2=Tl=��h<����j���U-����+G⾋X!��
Y�<͊����>-ǿ}ΰA��(����� ���󿙊߿?�ſ����2��*�X�Od!��%�0���1��������@u<���<,��<�`.<0y}��T��Ľ*n���J��2~������ܧ�����   �   /��W\�rq��.�LľcK��wqs�2�+�̵׽fyZ��Ec�`�=<�<�@w<��&��g����Wf�|�����d1��d�㗌�����{�����̿O׿j�ڿ�ֿQ˿���!��MP����b�10����Y!��R�f�����r���_��#/<�w�<�Ѱ;�)���vz�x8�6<5��P}� B��>�Ⱦ���5�{&	��   �   y/H�J�C��A8�Pz&��%��d3��=B��ȩ<�TJ��tb�xy� ��;��U< @���ݧ����'��=���ɾ�~
��F4�*__�jU���o��(z��7@���������8E����͂�"�\�
2�8��A�ƾ;���+Q&������-�@�ɺ�-<�"�;𦠼�Yx��M�TFD�v������\��/��E�(�:���D��   �   �쇿�%��
R{�.Nd�"FG���&�X���Iɾ	玾��:�I/׽d�D�Xa/��;���;��G��N��p޽h�?��
��<;�a��^)��J��f�hc}�K���ꇿF#��jM{��Id�HBG�L�&����Eɾ�㎾\�:��'׽N�D�8I/��"�;p��;H�G��N�w޽��?���#@;4d��a)��"J�:�f��g}������   �   ��7����G�� �7ς�ڡ\�#2����1�ƾ,���bU&�C����4�@'ʺh-<�;�;����(Ox��E��@D�𞎾%���������(�$ :�_�D�<+H��C��=8��v&��"��^��.��m>���<��A�6hb�`Vy���; �U< ����m���V�'�$@�� ɾ�
��I4��b_�pW��=r���|���B���   �   ,�ڿ��ֿ�S˿j	��9#��?R����b��30�����$����f�ٷ��
r���_��/<|�<p��;@��8jz��/�w65�gI}��=��	�Ⱦ�龖2�#	�����X��j��(
��ľ�F���is��+�/�׽�jZ�@c�x�=<t�<�Cw<0�&�ƪg�%��[f�.���ʎ�yf1��d�����ϫ��ӝ���̿�Q׿�   �   T�U� �?���߿p�ſm����3��ߍX�qf!��(㾅���H 1�#����估n<���<���<�{.<XQ}�(T��Ľ�h��J��*~�L����ק�����l������N@��nY��f{u�h�@�`�������,�@#λ���<:8=�n=؁h<����l���W-�ߊ���I�XZ!��Y��Ί�ӷ��C/ǿ��'D�����   �   �-�\W����J��8���Ŀ:ա�.� �?�eW�<���n�]����*�/���X;do�<*S=��=h��<����ؤ�3���2hֽ���_.���F�	2V���Z�P�S��8B��'�T���_ý�<p�PüP��;��<V�6=f�D=VW=��7<|����ܽ�W�Y鲾�.�^�>���~���m.ſ���@[��&�����   �   �w+�0<(�pO�(��L+��7ݿ뗶������Z����g�Ҿ/������2�i� D��� =��E=��T=nn9=K�<x�/<�Q���8�{�����ʽ߽��併vڽm���@#��x�Z��t� H�'�<�4-=��h=�[�=��q=�(*=`��;RF��7�za}���ξ����X��ڏ����]ݿ�X�"1�8��4�(��   �   
P;�N�7���-����v����ƿ��4�o�?�,��������#��̌��X�&�=��^=B�=$V�=�*_=��(=�1�<0�;��8�Ƽx8��[.�
	5�"a%��� �����@���ೋ<V=·X=i��=8��=1�=��=��1=��[;Rq��K�𮍾Z��&�)�� m�������ſ����K����f�-���7��   �   ��E�
B��K7�|@'�������FHѿ�y��u*}�X�6�~����ǜ��g0�򋜽�-�$E=��l=Y��=��=���=��p=v�>=�N=�4�<�< �h9`Р�P�»��2�*�;X'y<���<�10=d<l=�&�=���=Q�=�ש=���=�4=��:c���Ψ%��Q��
���3���y�fˤ���Ͽm���xV�^'�G7��B��   �   ��!����N��D�	��7��c�п?!��������L��m��Tľd�q�o���B�04�;�d.=k%�=Y7�=z5�=Sϙ=��=,ew=R=r.=nM=���<X^�<4��<��<�=J&9=��d=�c�=��=Q,�=d��=���=�Q�= N�=־~=��<���E�"_d�����Y]�b�I������Ӫ�(�ϿC|�β	���l���   �   ��&�z�r���#��dͿ�(��j����'I�܉��(���l�m.��8c9�p}<$/=o��=m֕=��=�p�=�S�=^�_=��5=��=���<��<�χ<���<�ˣ<���<�W=��C=�w=zÕ=���=A}�=��=R'�=���=6�}=���<�X�gj޽�
_����Р�pXF��<�������x̿��$t���"/��   �   f��Z�<��.� �JQ�!*ÿ������|��>�+(����bZ[����\M��u8<�`0=�oy=gb�=���=��w=@-L=:K=p��<8�&<�Җ� ���yl�Pyu� !6��cG��< A�<��=Z`=��=�=<U�=�g�=Hä=V�z=�R�<�[ż��ʽ��O�5���Ҭ�߼;���z�������¿���� �����u��   �   |�
�va��Y����ѿ�(��� ����f���,��3���<��OA��½�V� w�<�S0=�)g=��q=@�Z=f�)=���< �;('\�j�t�G� T{�>ی��ꏽR��8_a�ډ!�� ���Z�:��<1=�_w=���=�]�=���=p2s=+�<�l��� ��Ty7�����/z�+�a�e�����t���(ҿ$��6��*���   �   �I������8�v�ҿ�n��O���������J�J��*ӾFu��)� ��ꗽ���̬<$�+=.�I=e:=��=�Z<�:��_ ��F���Ľ	��JH���������Ů�.���f�^�\ü���;�k�<pL="�}=Ov�=:6e=B�= ���υ����w��%�о����pJ��ہ��(��9&����ӿ�	�CC��   �   AտMѿ�ƿ�-��0����|��FP\���*�������֜]����H;Q�@�X�\��<�*=У=��<0��;Hwͼ�z���Ͻ���^<���`��
}�S��Չ������v��W�V�0�^������*?�0n(����<d�%=��Q=��M="'=r�;7��/�ybZ�a4�������m+��V]�,K���ˠ�L���
ǿe�ѿ�   �   ���k���#Y���𕿩����)^��U3�.�	��YȾ����t�&�k���\=� P<d��<~F=P�<@߼:��u����k��;�NHx�9}�������Ǿb�ԾOaؾ|�Ҿ{�ľ��� ��k+l�}�.���<4��s���SL<b�=�)=�=Fk<(oƼ���tD&��L��G�ɾs�� 5�O`��섿g*���Y���@���   �   ����[�������&n�<P� >.�O� `Ӿ����_E��S㽼�H�@⾻�7�<`��<�G�<@6s;����N�����bU�'����*��^��d$�!����������x����/߾tw�� Ό��J�ޕ�Ir������R-<���<B�=�{�<@�����L��2�GGI��J����־`v�l�0���R��p�F􃿲B���   �   ĘX��S�G���4�l��`����̾�c��	R�F��J��������[<T�<���<0�4<�G����P4���Y������Ҿw���Z�>�6��gI���T�̜X��T�}�G��4�s�������̾�f��TR�!��O�����`�[<�Q�<���<��4<�8��S ��40��Y�+�Ҿ���rW���6��cI���T��   �   ,����ou�.���*߾s��{ʌ�J�d���k������j-<��<Ė=tw�<0骻��L��9��KI� N����־�x�x�0��R��p�a����D��ݖ����������)n��P��@.�bQ��cӾ���(dE��Y���H�����3�<���<�N�<`�s;�����G����IU�S���@&���~�^!���g���   �   �[ؾ��ҾA�ľ������5$l���.�����,��]��@rL<@�=X�)=v=x:k< {Ƽգ�� H&�PO����ɾ��m5�FR`�Vp,���[��(C���������B[����h����,^�X3�,�	��\Ⱦ������&������G�F<\��<�H=Z�< ۽:�t�ض���f�ԩ;��@x��x���{��S�ǾʆԾ�   �   �Љ�z�����v���W���0�����x���?��?(�࡞<|�%=<�Q=�M=T&=�W�; �7��4�fZ��6�����p+�5Y]��L��t͠�N��ǿ��ѿ�տ	ѿ�ƿ�/����,~���R\���*�����L��	�]�<����@Q�@�X�L��<,=��=H��< ˝;P_ͼ��z�Q�Ͻ����<� �`�x}��N���   �   +��E�� �ʣ�o�����^��?üpܦ;\}�<�vL=��}=�w�=�6e=�=�ҽ�҅��Xy����оu��sJ��܁�**���'��|�ӿ��UE�K�����:�4�ҿ@p����������m�J����",Ӿ�v��"� �C헽�
��Lˬ< �+=ުI=�i:=F�=�=Z< �9�jQ ��=���Ľ����5B�����   �   �ᏽVI���Na��z!�d���֞: ��<4$1=*fw=	��=E_�=���=�2s=t(�<,s�����e{7����D|��+��e��������)ҿ�����
��^�
�Rb�PZ����ѿ�)��m��n�f�Ԯ,�-5���=���PA�"�½[꼠u�<rT0=�+g=�q=�Z=Դ)=4��<�_�;��[� \���G�C{�cҌ��   �   PLu���5��F��<XR�<:�=�`=m��=��=�V�=�h�=�ä=B�z=|P�<�`ż՜ʽP�O�^�������;���z�t�����¿��r� �T���v��n[�Ы��� �1R��*ÿ����� }��	>��(����t[[�P���N��s8<,a0=qy={c�=B��=�w=�2L=�Q=Ǿ<��&<�������pMl��   �   �<p֣<���<l\=�C=|�w=�ĕ=���=5~�=���=�'�=���=��}=���<,\��k޽�_�9��M��YF�=��U���y̿���vt���~/��j&������-$�EeͿ )�������'I��� )��Al��.���c9�p}<�/=՝�=�֕=|�=�q�=U�=��_=��5=
�=|��<��<�ڇ<�   �   `��< ��<�=4&9=��d=�c�=��=@,�=M��=���=�Q�=�M�=f�~=��<��F彁_d�����~]���I������Ӫ�A�Ͽ\|�ز	���p����!����F��8�	��7��H�п#!��������L��m��Tľ�q��n�&�B��8�;Le.=�%�=|7�=�5�=nϙ=��=rew=PR=�.=�M=���<�^�<�   �   �<p֣<���<n\=�C=��w=ŕ=��=M~�=���=�'�=F��=�}=\��<�V��i޽8
_�4�����$XF��<������5x̿����s�8��.�P��%�"���%#�bdͿ?(������&I�Z���'���l��,���`9���<�/=c��=nו=��=r�=SU�=
�_=��5=D�=���<4�<�ڇ<�   �   �Ku���5���F�Ъ<dR�<H�=�`=���=4�=W�=�h�=~Ĥ=��z=TW�<�Vż�ʽ��O�k���F��"�;���z������¿��^� �$��Hu���&Z������ �;P�0)ÿ/���h�|��>�V'�����X[�M��8I���8<d0=0sy=Hd�=ꝉ=�w=l3L=�R=0Ⱦ<h�&<��������Ll��   �   �ᏽTI���Na��z!�T���ڞ:P��<|$1=�fw=u��=�_�=���=�5s=2�<�d��F����w7�T󜾉x�g+���e����e��G'ҿ���l��P����
��`��X�
��ѿY'��q���0�f�G�,�U1���:���LA���½�K�Ā�<pX0=�.g=\�q=ښZ=F�)=���<@h�;X�[�x[�f�G��B{�PҌ��   �   (��H��
 �ң�p�����^��?ü�ަ;�~�<�wL=@�}=�x�=�:e=��=`����˅�z�v���о���8oJ�~ځ�f'���$����ӿ�>A�oG������6濛�ҿm��Ӻ��h�����J�����'Ӿds��f~ ��旽�����ج<��+=j�I=Xl:=^�=�DZ< �9�0P �o=���Ľ����!B�����   �   �Љ�|�����v���W���0�����x��Z?�=(���<>�%=��Q=&�M=�,=��;D{7��*� _Z�2�������k+�T]��I���ɠ�3J���ǿ3�ѿ տѿ�ƿ�+��]���{���M\�p�*�#���c��ޘ]�����42Q��SX���<V1=��=L��<�ݝ;�[ͼ�z���Ͻ���l<�ݕ`�d}��N���   �   �[ؾ��ҾG�ľ������7$l���.�r�轐,���Z��XyL<�=��)=�=�`k< _Ƽԙ���@&�xJ��,�ɾs�?�4�L`��ꄿu(��W���>��g��&����V���ӯ��S&^��R3���	�NVȾ���z�&�h����*��o<8��<JN=b�<�=�:Dr�絙�,f���;��@x��x���{��J�ǾȆԾ�   �   .����su�2���*߾
s��xʌ��J�@��%k��h���u-<D��<�=��<P}����L�.,��BI��G���־�s���0�)�R�=�p�:򃿉@��s���-�������5"n��P�;.�sL��[Ӿܐ���ZE�3L��H�𗾻$H�< ��<�X�<��s;ؔ���F������U�,���!&���~�V!���h���   �   ȘX��S�ȘG���4�o��c����̾�c���R���II��������[<�_�<���<��4<�$������,���Y���Ҿ��dT�D�6��_I���T���X��S���G�&�4�F������̾�_��JR�Ȁ�C���w��P\< d�<���<��4<�1��	����/���Y���Ҿ���iW���6��cI���T��   �   ����^�������&n�BP�">.�O�`Ӿ����_E�%S㽨�H�Ⱦ��A�<���<�]�<�,t;�����@��_��>U������!���y�h���������-r�.��O%߾en���ƌ�� J�j���c��hﵼ�-<���<��=���<����ЍL��1��FI��J����־Rv�a�0�~�R���p�G􃿴B���   �   ���n���&Y���𕿬����)^��U3�-�	��YȾ����6�&������7� a<,��<�O=$j�<��:h�㮙��a���;�n9x��t���v���Ǿ?�Ծ Vؾb�Ҿ��ľ���o���l�@�.�S�轥$��C���L<̝=��)=�	= Zk<hƼĝ���C&��L��$�ɾe�� 5�
O`�}섿f*���Y���@���   �   FտOѿ�ƿ�-��2����|��HP\���*���������]�J���&9Q� �X�ȳ�<2=l�=ܯ�<��;�Eͼ��z���Ͻ���<�z�`�H�|�mJ��N̉�+�����v���W��0�����n��n?��
(���<�%=r�Q=v�M=�,=���;�7��.�bZ�?4�������m+��V]�(K���ˠ�L���
ǿg�ѿ�   �   �I������8�y�ҿ�n��R���������J�H��*Ӿ6u��� ��闽�����Ԭ< �+=Z�I=$p:=R�=�eZ<��9��B �:5���Ľ����)<�H��������������dy���^�H"ü?�;���<�~L=~�}=�z�=n<e=��= ����ͅ�F�|w��
�о����pJ��ہ��(��9&����ӿ�	�GC��   �   |�
�xa��Y����ѿ�(��� ����f���,��3��}<���NA���½�R��|�< X0=�/g=��q=�Z=�)=���<p��;`�[�N�>�G�<2{��Ɍ��؏��@���=a��j!�0餼�b�:,ջ<-1=�mw=��=�a�=���=�6s=�1�<Xh�� ��y7�n���z�z+�^�e�󢒿t���(ҿ%��6��*���   �   f��Z�>��/� �LQ�#*ÿ������|��>�+(����NZ[����,L��|8<�c0=�sy=e�=3��=��w=:8L=|X=�־<0!'<�[���� !l�Xu�`�5�@F�h�<Xd�< �=~`=T��=i�=�X�=>j�=GŤ=B�z= W�<�Xż(�ʽ��O�$���̬�ڼ;���z�������¿���� �����u��   �   ��&�|�r���#��dͿ�(��i����'I�݉��(���l�H.���b9���<r/=_��=�ו=b�=�r�=mV�=��_=R�5=B�=��<�<�<|͇<�< ��<:a=t�C=d�w=�ƕ=x �=r�=���=�(�=���=��}=���<<W�'j޽�
_�x��͠�nXF��<�������x̿��&t���$/��   �   �����h��Ӓ쿒�ؿ ���U��F`��:�P����۾���i+�;��HY����<N�@=�\�=���=��=��=�;�=��{=*d=nwN====�2=�R0=�B7=�G=da=xi�=w��=�ة=I�=�;�=�F�=���=�&�=r0�=�m�=�9G= #G;B�{��=��h���Ծ���4hN�k���Y������tؿ����m���   �   d���>��!��Lտ�B���>������0�L�Zy�+�־@�����&��ߢ�`Ȣ��O�<�FB=/��=i�=�!�==`��=B�i=�/N=��4=� =�e=e=�="y&=�mA=�
e=<y�=]��=#�=��=J��=l��=���=)%�=@�=8yI=�C�;�Hq�p"�}_���bоg��l�J���������ỿn�Կ����K���   �   ud�+�sݿ�pʿ�ǲ�� ���x�ُA�M���Cɾ"���C��x����f�t��<�1F=�k|=���=���=��w=ڛW=F�1=��
=���<��<ضM<�)<H�9<t��<|�<�	=��<=��s=�:�=�<�=%&�=��=.��=���=��=�O=��<��R�X3	�y���þB��O�?��v�S�������@�ʿ�Mݿ�O��   �   �Nڿ�[ֿ2˿�㹿F����^b���/���������Kh��=���g������,�<�J=�er=p*x=�/d=��==v�
= ��<P��;���x����������x	㼤����k����7<�t�<fF@=�j�=�?�=��=h%�=���=�W�=ptW=`�s<P�#�H5��]�2����b ���.�)�a�W���%���@����˿'�ֿ�   �   �¿Is���b��ʤ����Eu�(�F�b����ྨ����tB��Uӽ�I ��·;��=v`L=��`=�Q=|�&=��<��;��z�T�� �l�i��{���ޥƽ>ɽy<�����Ԍ~�*J$�������<�b=ZDY=<�=:֠=�Ť=Y��=p�^=��<��Ҽ�O���:�\ꗾr߾sI��F���u�����i���󴿄ʾ��   �   �v��G���q���ǌ���v���O��m'��W ��ӹ��cz������������<�t!= wH=�C=d�=��<�i���-� ꁽn�ý�1�����1�H�>�~�A��X:�d)��8�1⽹�����,�`��4�<�2=v�w=)�=���=�ab=���<��%�������Նx�繾*� ��\(�^:Q�ԋx�♍��!�������   �   �t������\^~�y$g���I���(����[̾fK����=�0�׽�t4� ��7�3�<�1= �;=�0=�)�<����,,�v��l��HG0��_]�&����������$A�������7����y��"O�ϒ���ݽ�C��d\����;<�=z�[=��t=��_=&=p��;��)�IE׽{�?����V�ξ���`�*���K�_i����"���   �   k�Y�V U��H�͟5�������jξs����S����E]����v��&�<��=�9=��#=l�< ���7.�}��}��j�R�^����G�ľ�Eھ*����뾹��}�־����F��������xC����蘽��开�<�c=~�H=��S=0M,=t��<\z���Y�����~W[��ߝ�K!ӾI?�!	 ���7�HNJ�}�U��   �   �$��� �$��)��`��]����X���V�\��g�����μ �;<[=��==P=8= ��<@Ǥ;�	�"s��d&�T2b�������ž}M�,'
������!�J�$��� ������*��t���>\��+%V���������μ�q;<�W=��==(>8=8��<���;�	��l�� "��,b�����ž�H�b$
������!��   �   Q��b��p�־���4���e����rC��������$��`�<�h=N�H=��S=�K,=���<�����^��7��R\[�"㝾?%Ӿ�A�� �	�7��QJ�  V���Y��#U�*�H�Ϣ5����
���nξq�����S�P��7b����v���<�=(�9=H�#=��< ����,.�F	��ˊ���R�ƪ��Y꨾��ľ�@ھ����   �   �<��.���f3��h�y��O� ����ݽ^<���D����;<x�=��[=��t=��_==�d�;
�)��J׽V�?������ξ�����*���K��i����a$���v��S����a~��'g���I���(����^̾�M��\�=�`�׽|4� ��7�.�<��1=��;=�4=�5�<����,��n���{�|A0�Y]�T������!����   �   ��A��Q:��])� 3������,��s�8��<D�2=��w=�*�=I��=~ab=���<��%�������x��鹾�� �_(��<Q���x�����#��h����x���H��qs��Ɍ���v���O��o'�pY �_ֹ�\gz�R��x�������X��<&t!=�wH=��C=�=4�<� ���!��⁽t�ýR,�&��P�1���>��   �   �Ƚ�2����P{~��:$��ۀ���<l=�KY=��=&ؠ=�Ƥ=���=��^=\�<H�Ҽ�S����:�8엾�t߾K��F�,�u�k���k��1���,̾�w¿�t��"d��kˤ�K���Gu��F�ϓ����E����vB��Xӽ�M �ஷ;��=�`L=`�`=*�Q=v�&=0�<`F�;(�z����\�l��������כƽ�   �   z�������0	���8<���<�N@=Bn�=�B�=���=�&�=H��=�W�=�sW=��s<~�#��8��]�·��d �0�.���a�V���&��?B���˿��ֿ4Pڿ7]ֿH3˿�乿N򣿵���_b���/�p������Mh�?�B�g� ����*�<�J=�fr=�,x=<3d=d�==
=ȯ�<P��;���~��l�����   �   X�9<8��<h��<��	=��<=ΐs===�=�>�=�'�=�=��=2��=��=�O= <��R��4	�My��þ��Z�?�X�v��������+�ʿ�Nݿ�P�xe�,�[ݿ�qʿ�Ȳ�����x���A����Dɾ���~D�z��P�f�0��<�1F=�l|=x��=���=��w=�W=\�1=��
=��<���<��M<>)<�   �   p�=r}&=�qA=He=�z�=���=Q$�=���=��=���=��=J%�=!�=txI=�8�;Kq�;#�`��Ecо����J� ������b⻿��Կ��YL������>����迳տ)C��?��������L��y���־~���,�&��ߢ�8ɢ��O�<�FB=f��=mi�=7"�=���=k��=֛i=�2N=.�4=� = j=di=�   �   �B7=�G= da=vi�=o��=�ة=�H�=u;�=�F�=v��=�&�=R0�=�m�=j9G=�G;�{� >��h��)�Ծ��[hN�$k��Z������tؿ����m�������h��ƒ쿀�ؿ�B��2`���P�e���۾����i+��:��X����<��@=�\�=̛�=��=��=<�=��{=J*d=�wN=6===��2=�R0=�   �   ��=�}&=
rA=^e=�z�=���=\$�=���=4��=$��= ��=�%�=��=�yI=`J�;�Gq�"�>_��)bо)���J�l��G����ỿ�Կ!��OK��ۣ��y=������տVB��N>��^�����L��x�^�־������&�,ޢ�Ģ�hS�<hHB=��=�i�=�"�=��=���=n�i=T3N=��4=L� =Fj=�i=�   �   P�9<���<���<�	=�<=��s=V=�=�>�=(�=W�=o��=���=��=ԂO=��<��R�g2	�7y���þ�����?��v��������s�ʿ�Lݿ�N�sc�*�uݿ�oʿ ǲ�0 ���x�ŎA�p��XBɾ$��)B��v����f�x��<�4F= o|=f��=���=\�w=,�W=l�1=��
=L	�<쳐<p�M<h?)<�   �    � �⼸��� ��`8<\��<�N@=nn�=�B�=X��=X'�=*��=Y�=|wW=8�s<�#�l2��]�߄��b ���.���a�|���$���?��~�˿ֿ̚jMڿxZֿ�0˿I⹿ ����S\b�0�/�j�����fIh��;���g�`���(5�<�J=�ir=V/x=�5d=T�==��
=ಡ<��;���0}��$�缂��   �   ��Ƚg2����>{~�x:$�pۀ��<ll=<LY=q�=�ؠ=Ȥ=[��=t�^=���<��Ҽ?L����:��藾�o߾
H�Q�F���u�ׇ��0h����Ⱦ�"
¿�q��a���Ȥ�� ��OCu�!�F�����ྨ����qB�;Qӽ�B ���;��=�eL=4�`=T�Q=*�&=��<�V�;�z�T���l�&��������ƽ�   �   ��A��Q:��])�3��⽵j�,�@r����<J�2=$�w=�+�=��=�fb=,��<�%������,�x��乾�� ��Z(�8Q��x�X���# ��Ԫ��u��EE��p���Ō��v��O��k'�V �1ѹ��_z�������0y��\��<�z!=}H=��C=\= ��<��|��ၽ�ý�+���"�1�e�>��   �   �<��,���f3��g�y��O���b�ݽ+<��`C����;<�=�[=D�t=*�_==�;�)��?׽�~?�q��&�ξ�����*���K�;i����� ���r�������Z~�2!g���I��(����-X̾�H����=���׽�j4� �
8XA�<��1=��;=�8=�<�<P����,�em��({�A0��X]�5���z������   �   N��_��p�־���3���a����rC��������8��x�< k=��H=��S=jS,=д�<�h���S�����R[��ܝ�zӾ�<�q ��7��JJ��U��Y��U���H���5�7��X���fξ+�����S�߿�W���v��6�<�=��9=v�#=�< i���).�	��B���R�����4꨾q�ľ�@ھ����   �   �$��� �&��,��c��]����X���V�<������ ~μ��;<N^=��==vD8=T��<@9�;\�	��e����''b��{����ž�Cﾧ!
����]�!��$��� ���_��b�����AU���V����'����iμ��;<�b=��==pD8=ؽ�<p�;�	��k���!�H,b��~����žkH�Y$
����~�!��   �   n�Y�Z U��H�џ5�������jξm�����S�����\��`�v��,�<@�=P�9=��#=��<�5��$ .�|������R�0���.樾ܖľ�;ھb��������H�־U������������lC�����ؘ�̙���<�p=p�H=d�S=�R,=讟<�s��EX����W[��ߝ� !Ӿ8?�	 ���7�ENJ�~�U��   �   �t������_^~�|$g���I���(����[̾\K����=���׽ds4� `�7�:�<h�1=��;=�;=�F�<�Q��6�+�Hf���v��;0�6R]�����e������A8��ˠ��8/����y�O�)��t�ݽ4���)���<<8�=��[=�t=�_=�
=��;�)�/D׽�?����/�ξz��T�*���K�\i����"���   �   �v��G���q���ǌ��v���O��m'��W ��ӹ��cz����[���Є��<��<Ny!=>}H=��C="=� �< ��v��ځ�wý�&�&����1���>���A�K:�(W)�!-��l圽Ж,� ?���<�2=Իw=�-�=��=*gb=D��<��%����d��|�x��湾� ��\(�V:Q�ϋx�ᙍ��!�������   �   �¿Ms���b��ʤ����Eu�'�F�b����ྞ���xtB�PUӽ.H � Է;ғ=LeL=T�`=�Q=|�&=L*�< ��;�z����"�l�����B�����ƽ��Ƚ^(���製di~�v*$�p���`<4v= TY=n�=
۠=�ɤ=��=��^=��<`�Ҽ O����:�:ꗾ�q߾hI��F���u�����i���󴿈ʾ��   �   �Nڿ�[ֿ2˿�㹿H����^b���/���������Kh��=���g� ����1�<t�J=vjr=1x=v8d=��==B�
=h��<�H�;�e�le���缶��
q�,��̄��𣡻�38< ��<6W@=�q�=�E�=���=�(�=5��=�Y�=nwW=�s<��#��4�`�]�����b ���.�&�a�V���%���@����˿'�ֿ�   �   yd�+�tݿ�pʿ�ǲ�� ���x�؏A�K���Cɾ���C��x�� �f�x��<�3F=o|=冈=e��=�w=��W=�1=��
=x�<�<P�M<(b)<��9<4΀<��<��	=X�<=V�s=@�=A�=�)�=��=|��=���=��=΂O=��<��R�"3	�Vy���þ>��K�?��v�R�������A�ʿ�Mݿ�O��   �   f���>��!��Lտ�B���>������0�L�[y�+�־=�����&�hߢ�hǢ�DQ�<�GB=�=j�=#�=���=� �=��i=�5N=��4=҉ =$n=�m=ԫ=́&=$vA=8e=�|�=w��=�%�=���=��=܋�=���=
&�=��="zI=0I�;ZHq�T"�r_��zbоe��j�J���������ỿo�Կ����K���   �   ~���������^���؏�?1s�}E�Ȃ�QZྑ�����G���xSJ��ɹ����<.*-=�+X=�l=��p=��l=��d=>�[=BT=J�O=VaO=��S=$:^=��n=�v�=o��=�&�=L�=���=��=J��=V��=hP�=T��=P��=��=��=�'=�E����+�2������WھqK�RwC�Qr�h���ei��K��#���   �   �<��DԹ�� ������K����n��ZA�����۾H���/�B�<Sܽܒ?� �y����<T0=��X=jzj=l�l=�f=Z�Z=��N=hhD=V�<=�9=HE<=�E=(�T=�k=��=�r�=R��=u�=�|�=��=8]�=��=���=X��=||�=�Y�=F=�=r������7.�=L��j�վ�q���?�k�m�	��~������O޹��   �   �����r�����(l��3ᅿ��a�j�6�����+ξ�ˍ��3���ƽx[ ���:���<��7=�'Z=Ze=��_=TQ=�== �'=@�=N=p��<�<�r�<�=��=��;=T`c=k�=��=���=$r�=��=�O�=��=��=�k�=?�=��=��v���!!�p���9Mɾ�+��5��[a�0̅� }��;-�������   �   �פ�ġ�����v��Ȑt�h�M��%�R���N��:�{�G�*���hl߼xd <j}
=x�B=KZ=�Y=�jH=@�+=t�=,[�<�z< ��;@��: E/���j��ߝ����;��^<(��<�* =R�\=!r�=~=�=pg�=��=��=c<�=�M�=2�=ZN,=�����v�����
q�莵�:����W%�@�M�P�t�����vM����   �   �ؑ��
��5)��Z�u��W�OT4�o��U[ܾ�q���S�ƭ��H�r��.I���<�$=hhM=�`V=�4F=�&#=�K�<��f< Q��z�t���F&��G��CV��Q�a8�Jd��r�� �x�(]�<�=�j=ʉ�=���=��=�g�=�N�=��=
l@=��<�i2�Zo�Z�L�Ξ���۾�����4���W���v�����yH���   �   z�x�؊s�o�e��tP�ߗ5�e|�&�lƵ��q���$&� ����L��9�;<"�<$�==@�T=`?K=�&=��<X_<��Q�+�`�n�*l���4ɽbM����������a˽�ʢ��b�xE�@�ֺ�^�<�@=��=2?�=�ڬ=∩=t�=^�S=���<H�μ�|����#�������?-�x��67���Q�)�f��#t��   �   �QK�-G��Y;��^)�����D���͍���B����6g��t0�ȭ�<"�,=|�T=�8V=>�5= ��<�%<�R���F�XC��������^2�!H��U���W�p|O��=�j "��� �]���Y�4#��БW<\!=��q=���=J1�=� �=��c=p9�<py߻X�f��A���/H�S\���Kþ+:����9!+���<���G��   �   �%������WE����XӸ����M�2�Jڑ��߼�0cY<B=TeU=�@e=��N=tU=X�c<pԁ��U�|��,}�4H>��Dl�nh���#��ʣ��W��`u������̬���[��)��X�r����=� *�;�=*�`=ƅ=x�=��l=�� =00'<��ᵤ�_�4Z�i+��@̾�2'羸}����za��   �   5�7�8�׾����垣��v���?E�����L���P���<�)=�qX=v�v=��m=��<=T��<������:�Ľ��Ќ���V�)t��Ǌ���ƾG�۾����羽�׾Ɨ�������y���DE����nS��@d���<x$=�nX=��v=ȅm=j�<=���<�r���}:����������V� q������ƾ��۾���   �   |S��Tq������H���l�Z���)��O�I~��L'� o�;t�=��`=]ǅ=��=�l=� =�'<X������b��8Z�Z.���Ͼ�a+���8��,d�L(��������G�����ָ�����N��"��ߑ��＼hLY<~=DcU=j@e=�N=VX=8�c<�Ł���U�����x��B>��>l��d������ţ��   �   ڝW��uO�n=��"�t� ��
��x�Y�d����W<�!=��q=���=L2�=/�=j�c=d3�<�߻@g�sG���3H��^���Nþ>��Y���#+���<�k�G��TK��G��\;�a)�6��6�G��Ѝ�{�B�% �^>g�`�0����<��,=|�T=9V=B�5=���<�<<pB���F�[<��������"Y2��H�Z U��   �   �������;X˽������b��)뼀Iպr�<8$@=��=VA�=Yܬ=���=r�=��S=<��<,�μ �����#����n"��r0�h��t7��Q���f��&t�T�x���s��e��vP���5�5~�%��ȵ��s���'&�0����R�@�;�<��==4�T=�@K=ή&=P%�<px<ȵQ�< �.�n�ed���+ɽ�C������   �   ��Q��Q8��U��W����u�@r�<�&=~�j=���=���=1�=�h�=O�=���=Xj@=H�<(o2�Js��L������۾f����4���W�*�v�Ǔ���I��ڑ����i*����u��
W��U4�ϊ��]ܾ�s��j�S�w�����r��=I� ޣ<�
$=
hM=xaV=�6F=�)#=�T�<�f< O�xS�Hl��9&���F�x4V��   �   ����0L�;(_<\��<Z3 =�\=[u�=$@�=�i�=l��=  �==�=!N�=��=�L,=@m��T�v�N���q�����P����X%���M��t�󻋿�N��'��ؤ�š�����w��d�t���M�:�%�������E�{���R���xr߼0\ <.|
=��B=\KZ=2�Y=�lH=f�+=ԝ=pf�<��z<`:�;���:��.���i��   �   �=��=R�;=xfc=7�=m��=�¶=�s�=D��=�P�=���=�=�k�=� �=:�=����w��$#!�_���vNɾ�,�܋5��\a��̅��}���-��i��������s������l���ᅿ��a�/�6�G���,ξb̍��3� �ƽx] ����:���<��7=�'Z=
e=B�_=XQ=�==��'=��=�=<��<�*�<|��<�   �   ��T=@k=B�=t�=���=7v�=�}�=��=�]�=4�=��=|��=l|�=�Y�=
E=8Dr�����n8.��L��,�վxr�}�?��m�o	��䞠�^���޹�X=���Թ�#��L���GK����n�3[A�`��_�۾������B��Sܽ��?���y����<20=��X=�zj=�l=�f=��Z=��N=�jD=��<=��9=tH<=�E=�   �   ��n=�v�=s��=�&�=L�=���=��=<��=H��=\P�=@��=8��=��=鳏=('=LG�����r�2�道��Wھ�K�swC�qr�w���oi��T��'��}���������R���؏�1s�_E���� Z�e���>�G�����RJ�ƹ����<l*-=�+X=�l=��p=��l=��d=f�[=NBT=t�O=�aO=��S=B:^=�   �   ޖT=lk=S�=t�=���=Dv�=~�=��=�]�=Z�=D��=ȱ�=�|�="Z�=�F=0:r�'���07.��K��	�վ�q���?���m����/�������ݹ��<���ӹ�] �������J����n�DZA����0�۾����@�B��Qܽ��?���y����<�0=
�X=|j=>�l=�f=��Z=��N=|kD=��<=��9=�H<=H	E=�   �   n=�=��;=�fc=O�=���=�¶=�s�=t��=Q�=���=��=]l�=�=��=p���t��� !�����LLɾf+��5��Za��˅�~|���,��ߊ��ﹳ��q��&��nk��������a�f�6����R*ξ�ʍ���3�8�ƽ�W � }�:��<��7=t*Z=te=v�_=bQ=�==B�'=(�=�=X��<�,�<ȁ�<�   �   �l��0P�;�_<���<�3 =4�\=�u�=Z@�=�i�=΁�=� �=�=�=9O�=��=fQ,=������v���xq�����t���zV%���M���t����yL���֤��¡�~���u����t���M���%�!��������{�<����|b߼Hu <<�
=:�B=OZ=��Y=�oH=:�+=`�= k�<�{<H�;�ۙ:��.���i��   �   ؛Q�0Q8�VU��V����u��r�<�&=�j=��=W��=��=�i�=wP�=���=p@=��<�c2�ek潾�L������۾����4���W���v�U���4G��jב�^	���'���u��W�uR4�އ��Xܾ�o��ˁS�����r� I���<�$=,mM=�eV=�:F=z-#=h[�<`�f< ^N��I�@h�"8&�L�F��3V��   �   J������X˽������b�)� =պs�<�$@=X�=B�=\ݬ=	��=��=�S=�ˡ<L�μjx����#�%���s��8*��� 7�5�Q���f�!t��x��s���e�rP���5�jz���õ��o���!&�����D��m�;�-�<��==� U=�EK=8�&=`-�<8�<��Q�B���n�Oc���*ɽC�h����   �   ��W��uO�V=��"�d� �z
���Y�`
��0�W<�!=J�q=���=�3�=n�=ܢc=�E�<@=߻��f��;���+H��Y��{Hþt6������+�N�<���G�OK�RG�&W;�$\)������PA���ʍ�{�B����+g��S0����<6�,=`�T=�>V=L�5=���<@M< ;��ĂF��:��C��>���X2��H� U��   �   jS��Fq������B���_�Z���)��O�~��&�v�;ʓ=��`=�ȅ=)��=.�l=� =�N'<�t�ԯ��?[�2/Z�p(���Ⱦ�#�c{����^��"�I��u���B���ᾤϸ���n�M�,��ӑ��˼���Y<=�kU=,Ge=��N=:]=��c<Ľ���U���!x�LB>�*>l��d������ţ��   �   *�0�5�׾����➣��v���?E�t���L���N��<x+=�tX=x�v=��m=��<=���<�(��r:�n���I��$�V��m��S����ƾ�۾	�I�]羖�׾^������qs��:E� ���E��X9�8�<J1=�xX=� w=�m=��<=���<�R�� z:��������V��p��݆���ƾ��۾���   �   �%����
��VE����VӸ���m�M���ّ��ݼ��iY<�=�hU=Fe=8�N=t_=P�c<������U����t�L=>�28l�Ha���������JO��1m������������Z��)�fF�mv����`��;Ԛ=�a=yʅ=���=*�l=8� = @'<��V���b^�j3Z�%+��̾�'羨}����ua��   �   �QK�,G��Y;��^)�����D���͍���B�7��,5g�0o0�ȱ�<�,=ҹT=�>V=��5=���<�a<,���xF�V4��3��l��.S2�nH���T��W� oO� =��"�$� �X����Y�񔼰�W<b!=$�q=���=5�=��=b�c=PA�<�^߻p�f��@��>/H�\��^Kþ:����/!+���<���G��   �   �x�ڊs�s�e��tP���5�e|�$�fƵ��q���$&�̄���K� F�;'�<��==B U=PFK=h�&=5�<��<H�Q�,��n��[��G"ɽ�9�]�������E��/N˽����*b�T뼀�Ӻ$��<-@=��=bD�=�ެ=��=��=P�S=Lǡ<̗μ�{��j�#�Է�����-�j��,7���Q�%�f��#t��   �   �ؑ��
��7)��]�u��W�PT4�o��S[ܾ�q��ЄS�������r��)I���<�$=JlM=*fV=$<F= 0#=�c�<8�f<��L��$�R�r+&�L�F��$V�~�Q��A8��F�l;����r����<J0=��j=.��=���=��=�j�='Q�=���=&o@=��<�g2�sn���L�������۾�����4���W���v�����zH���   �   �פ�ġ�����v��ʐt�h�M��%�P���J��*�{�.�䍤��j߼�i <\
=D�B=�NZ=L�Y=�qH=��+=P�=du�<�{<���; ��: �-��$i� �� ��;H1_<x��<z< =�\=�x�='C�=l�=���=��=�>�=�O�=��=�P,=�џ��v�@��L
q�ˎ��#����W%�;�M�M�t�����uM����   �   �����r�����)l��3ᅿ��a�h�6�����+ξ�ˍ��3�d�ƽ�Z � 6�:��<��7=(*Z=�e=p `=Q=�==v�'=&�=�=d��<�8�<���<4%=�=0�;=�lc=%�=��=Ŷ=�u�=���=:R�=د�=(�=�l�=(�="�=8���u���!!�Z���(Mɾ�+�݊5��[a�0̅�}��<-�������   �   �<��EԹ�� ������K����n��ZA�����۾G���(�B�"Sܽ��?��y����<40=��X=|j=��l=Vf=��Z="�N=HmD=��<=�9=�K<=bE=�T=�k=� �=�u�=��=�w�=�=��=�^�=��=���=��=}�==Z�=�F=P;r�~���z7.�4L��c�վ�q���?�j�m�	��������P޹��   �   �q���Ԉ��G��Vk�tcM�M(,�[
�)LӾm_�� JQ�����������@C-�Pn<�A�<<��<TZ�<�A�<Ty�<��<�(=>�=�%$=�]9=B�Q=>�m=�΅=��=<T�=�U�=�t�=$��=��=���=��>n>O�>��=���=1�=d�v=�t�<в���Ƚ$.:��E����;^\� +���L�\�j��C���׈��   �   q����b��g�}���f���I�H�(��V���ξ�╾��K�g2���ǋ�`�� <H�hj�<p��<do�<(��<�7�<�;�<̴�<,-�< '	=�=��*=�EA=�\[=<�x=p�=��=<p�="C�=���=�[�=6��=���=��>�N >RW�=+�=jT�=�'y=�H�<�,꼍���ġ5�@#���ɾ�����'��I�ڢf���}� j���   �   dā�4�~�FYp��DZ�Ch>�<?����U���[Ƌ�Sd<�̀�lIs�'��@��;(�<C�<ȥ=j(=t��<���<��<��<$��< L�<���<��=h�#=�b>=.+^=L�=PQ�=iU�=�M�=:�=4-�=�\�=���=H��=0/�=��=��=��=�E�<�ƺ�����n�(�$������E�����B>��^Z�g�p��~��   �   Lm��]h�-[���F��-��E����<ݭ�Bx��$�o½Vt:�`�'��eW<���<�M	=j�=@o=p��<�r�<Q�<Ļ�<�wT<��9<P`7<H<Q<�O�<D��<D�<��=vLM=�+==>�=��=�l�=��=��=�~�=f�=��=��=�N�=�*�<He�����b@�; n��'��
���@�(R-�3G���[�ԟh��   �   �\P�x L�E@�Z�-�N��o����2ƾ�k���P�AH��3��X��@�b;ܪ�<��=� =Db=��=�e�<dĒ<�<�F/:�3��F[�P���a��������p������d;8r�<Ħ=<&D=a�=H��=��= C�=��=���=���=a�=��=��= 5P�~b�����^K��ѓ���ƾ�������.���@�X�L��   �   ��/�9,���!����0����ϾB���9�o�N�"�>�Ľ@*;��l����<.�=��2="�7=L�&=X�=H��<�p�; [ֻ4a���{��^D��*n��܄��ĉ����&Rj���7����x����@<n=�V=I܎=T�=��=���=�J�=���=6�=��0=		<��TO���+$��s�����p<Ӿ�}��Cr���"���,��   �   �e�&��^��꾭�Ⱦ������{�$4����X�w��p��h�Z<� =�'B=��T=�*K=�7*=T��< �H<0��$��R�P�����z���q�̖����������zwܽ�㱽R(}�,����ػ`��<��0=
�=�؜=���=;j�=�Ԧ=!�=�F=�ܞ<����o��մ����>������Y��A�;C�,������   �   ��۾�־o�Ǿ�ݱ�����`q�6)4���:ዽ��ϼP�<bG=$VN=ʉo=8�q=��W=�!$=|��< �Q����zLl��������4}���7�:}L��uX��LZ�*�Q�}�>��#��.��麽LS`�,����4<v�=,yi=q�=���=u+�=�g�=��T=d	�<��f%�ǯ�V�P�F�tM��f*��ռ���˾d(ؾ�   �   2q�������Տ���|��R�V�"�^i佊j��L3ؼ ��;H7=�Z=��=Gg�=ư�=V�Z=��=�i@<<˖�Q]�q	�����~�:��=f��W��5���=���t��z����؏���|�L
R��"�q��p��`Gؼp��;<1=&Z='�==f�=P��=��Z=@�=�w@<���I]����-���:�I8f��T���1��`:���   �   �FZ�D�Q�߻>�À#�	*��ẽ�E`�H��Ƚ4<d�=~~i=h�=���=:,�=�g�=��T=`�<�]�%��˯���j�F��O��c-��=���׻˾S,ؾ��۾�־#�Ǿ�౾��eq�z-4���拽��ϼ�<hB=xRN=N�o=q=��W=�"$=p��< �P����zCl���������x���7��wL��oX��   �   >������Mnܽ7۱�}����ػ�͡<4�0=��=ۜ=Z­=Jk�=>զ=�=F=�֞<����r�����\ ?�ٿ���\��{�;�F�,������g�;��`���گȾd����{��4����,�w��~����Z<��=�$B=֣T=�)K=>8*=\��<��H< \�(����P������s���i�������   �   ����"Cj�@�7����X���
A<j'=��V=Lߎ=��=P��=*��=�K�=ܘ�=�5�=�0=H�<P��GS��j.$���s�ׯ��<?Ӿ���t���"���,��/�/;,���!����3����Ͼz���Êo��"���Ľ�0;����4�<<}=��2=��7=��&=�=@��<���;�1ֻHS���r��SD�n��Մ������   �   h^p��y���e;���< �=X.D=ׂ�=*��=��=�D�=:�=��=��=t�=M�=��=�lP��!b������K��ӓ���ƾ�������.���@�L�L��^P�e"L��F@��-��������4ƾom��XP�4J��6��x���wb;P��<��=�� =�a=��=0h�<�Ȓ<`< �0:���'[��	��HM���}���   �   Pǲ<@&�<|�=�SM=`2="A�=f�=�n�=���=�=��= �=R��=��='N�='�<�e����B��"n�")����B�yS-��4G��[�w�h��m�=_h��.[��F�-��F�n�徑ޭ�Yx�J $�vq½x:���'�p\W<��<^L	=��=o=���<�u�<�U�<�<��T<��9<z7<�XQ<L_�<�   �   �g>=T0^=�N�=�S�=�W�=�O�=��=�.�=�]�=���=���=�/�=$��=��=ҟ=�B�<�˺�������(�	��F����F��ǭ��C>��_Z���p�K�~��ā�Z�~�XZp��EZ�i>��?�A���?���ǋ�de<�k���Ks��*��p~�;��< A�<4�=,(=��<0��<���<T��<���< S�<Ȝ�<�=^�#=�   �   ҝx=Hq�=��=dq�=&D�=l��=b\�=܁�=���=ѱ>O >pW�=
+�=<T�=�&y=|F�<X0�ÿ����5��#��иɾ���q�'�^I�r�f���}�qj������8c����}�V�f�V�I���(��V��ξH㕾��K�3��`ȋ���� hH�0i�<h��<�n�<���<8�<P<�<H��<h/�<z(	=��=��*=�GA=B_[=�   �   �΅=��=DT�=�U�=�t�= ��=��=���=��>�m>J�>��=���=�0�=�v=�s�<(���OȽf.:��E����;v\�& +���L�n�j��C���׈��q���Ԉ��G��Ck�^cM�5(,�D
� LӾJ_���IQ�̬�F������ ?-�n<�A�<x��<�Z�< B�<�y�<T��<$)=p�= &$=�]9=h�Q=h�m=�   �   J�x=wq�=��=�q�=>D�=|��=x\�=���=���=�> O >�W�=^+�=�T�=\(y=pJ�<�*����T�5��"����ɾM����'�kI�b�f�b�}��i�� ����b����}�@�f�^�I���(�.V���ξb╾��K��0���Ƌ���伀�G�@m�<4��<\r�<P��<\;�<�?�<@��<2�<�)	=��=r�*=�HA=�_[=�   �   �h>=�0^=�N�=�S�=�W�=�O�=�=�.�=^�=���=8��=0�=ʞ�=���=v�=J�<P������X�(�p��4���bD��8���A>��]Z�U�p���~��Á��~�Xp��CZ�Ag>�[>��������_ŋ��b<�c~罒Es�� �����;\�<XH�<��=~+=P��<0��<���<���<p��< W�<��<p�=n�#=�   �   �ɲ<(�<&�=>TM=�2=bA�=��=�n�=ܯ�=r�=p��=� �=@��=
�=�O�=d1�<�d�!����>�n�F&��Y���?��P-��1G��[�9�h��m��[h��+[�7�F�z-��D���徙ۭ��x��$��k½2o:��'��tW< �<bQ	=j�=�s=`��<�}�<�]�<�Ɂ<��T<��9<0�7<X`Q<8b�<�   �   Yp��q껀�e;ć�<x�=�.D=��=l��=J�=fE�=��=���=4��=�=��=�=`�O��b������K�Г���ƾ�����U�.���@�k�L��ZP��L�#C@���-��������H0ƾ�i���P��E�50���㼀c;@��<�=�� =hg=N�=�r�<�Ғ<(<��1:���@[�x�� I��Pz���   �   ٠��Bj�x�7����0���A<�'=�V=�ߎ=&�=���=��=�L�=���=L8�=
�0=�!	<R���J���($�N�s�>����9Ӿ�z��up���"�k�,���/��6,���!�� �O-���Ͼȩ��)�o��"��Ľ";��6��|��<j�=�2=��7=J�&="�=̛�<p��;�	ֻJ���n�HPD�8n��Ԅ������   �   ��x����mܽ�ڱ��}������ػϡ<��0=��=�ۜ=Bí=�l�=צ=��=*F=,�<�����i��������>�=���W����;e?�,������c���\�4�N�Ⱦ������{�4�c���}w� `��h�Z<�=Z-B=X�T=�0K=�>*=���<�I<�/����Z�P������q��Hh�Ō��x��   �   �FZ��Q���>���#��)�`ẽxE`�,��p�4<B�=�i=G�=3��=�-�=Nj�=��T=`�<�� � 	%����������F��J��D'��T���N�˾c$ؾ��۾�־��Ǿڱ�񻖾C[q��$4�r��ۋ�d�ϼ0�<RN=>\N=��o=�q=b�W=�($=X��<�{O��⼐>l��������x���7�0wL��oX��   �   q��傛��Տ���|��R�<�"�+i�Ij��2ؼ���;h8=LZ=��=�h�=��=��Z=N�=Ș@<0���
=]��������:��2f��Q��c.���6���m��a��5ҏ�B�|�:�Q�b�"��`低c���ؼ�$�;
?=LZ=�	�=&j�=���=��Z=�=��@<ĵ��4D]����0��9�:��7f��T���1��6:���   �   ��۾�־b�Ǿ�ݱ�����`q� )4���������ϼ@�<�H="XN=��o=P�q=��W=Z)$=0��< �N����h6l���������s�!�7��qL��iX��@Z�~Q���>�R{#�(%�ٺ�`7`��룼 �4<��=��i=v
�=���=�.�=�j�=@�T=��<�� ��%��į�c �v�F�M��*�������˾C(ؾ�   �   �e�!��^��꾨�Ⱦ������{�4���罼�w�Xo��8�Z<$=*B=�T=R/K=�>*=���<pI<p�D��ХP�(���Kk���`�������������dܽDұ��}�����Bػt�<��0=�=ޜ=ŭ=�m�=�צ=��=VF=��<ܖ��,m������>�D����Y��	�;�B�������   �   ��/�9,���!����0����Ͼ<���$�o�8�"���Ľ�);�e����<�=��2=�7=��&=��=재<���;`�ջD=��^f�"FD�Ln��̈́�����]���3j���7�@���v�@8A<J1=��V=��=�
�=���={��=�M�=��=I8�=غ0=x	<����M��+$�y�s�L���:<Ӿ�}��5r���"�|�,��   �   �\P�y L�	E@�\�-�N��l����2ƾ�k���P�'H��3�����@�b;ȭ�<��=� =df=(�=Pt�<�֒<�4< �2:��x�Z���,5���d��x,p���`Gf;L��<ع=(7D=���=s��=��=ZG�=N�=ʐ�=���=[�=v�=��= P��b������K��ѓ���ƾ���t����.���@�V�L��   �   Lm��]h�-[���F��-��E����6ݭ�5x��$��n½�s:�p�'��iW<��<�O	=b�=:s=���<��<�a�<�ρ<��T< �9<��7<|Q<4q�<8ٲ<�7�<ڼ=�[M=�9=\D�=5�=q�=���=��=���=z!�=���=@
�=�O�=X/�<(�d�ɩ���?��n�{'�����@� R-�3G���[�ҟh��   �   dā�6�~�HYp��DZ�Ch>�<?����R���XƋ�Jd<����Is�&�����;�<�E�<��=
+=D��<,��<���<���<<��<D]�<���<��=�#=�m>=�5^=NQ�=0V�=�Y�=�Q�=��=(0�=,_�=���=���=�0�="��=π�=N�=�H�<ĺ�!���/�(�
�����xE�����B>��^Z�g�p��~��   �   q����b��i�}���f���I�H�(��V���ξ�╾��K�[2���ǋ���� &H�Xk�<���<8q�<���<;�<�?�<��<�3�<�*	=F�=,�*=�JA=b[=��x=�r�=D��=�r�=OE�=t��=J]�=���=>��=!�>OO >�W�=�+�=�T�=l(y=0J�<�+�D�����5�3#���ɾ�����'��I�٢f���}�!j���   �   S?�NW;��n0���Dc
�3��Q���/����F���A�����N����A���qM�@lQ�p0z�贒��n������ha]���л �M;�-k<���<f� =�]T=�C�=%V�=�?�=���=���=�]�=�v�=�+>�(>Z�	>a3>W�>��=���=�s�=��S=h�T<���ǽ!9.�F4��n����6㾯�	�nN��c0��Z;��   �   ֈ;�C�7��-�Gq�i���+�����򆾆�A�t���ϥ��cC�Sؼ�Rs�P|,��A2�pt]�L1��@}��l�� X��Kػ X;�S<ps�<��=�H=J�y=���=���=xT�=���=���=4��=x>4d>CF>z>>���=hr�==�0V=`�g<���P6���*���~����9�޾��TH��-�T�7��   �   1�ʇ-��F#��o�<��TbӾ���� {� u2����E����"�ܵ��H�� @��Pᱻ`��h�E��|m��tr��uL�@�� i﹨�<tA�<���<Zi$=*mR=E�=�.�=2��=�.�=,(�=J��=�j�=|>��>ޥ>`	�=�x�=T��=9$�=�U\=$ō<4�����3-���n�������Ѿ�������r#�M�-��   �   W� ���=�h�	H澼轾#����]�>��V�ǽj7g�d!߼���@٘:@�;��<;�S�� w�����8�D�X�F�Xi$� ��� p͸[�;�4|<8��<��=��9=��g=�ҋ=���=6��=���=0��=H�=��=�~�=
�=�7�=x�=A�=h�d=<��<����"�����X�U����/㽾����z����   �   �Z�6?	��� �UM�o�ƾ8���Q�|�Լ8�Z���ԗ�\��8�7����;��]<X�~<�%V<P< s�:������ �(�Z��Ax�P?y���^���(��ڮ� ��:� <��<t� =��4=��k=�}�=��=r��=&�=У�=�F�=t��=���=��=���=�Ml=�p�<P�;���p���f07�G��褾[8ɾ���/���	��   �   ȥ꾹��I־\i��b=��;,��L�I���^-���B���|�0��;T��<D��<��<���<��<�< �*�h��Y���gǼ<��W	�tZ��t�d��� �ɼ�y�`dB��i=<��<�5=�Mw=n��=ַ�=�D�=�<�=|l�=x��=��=}��=�p=�-=@��$B/�r�������S�tF�����jlþ��ؾ�z��   �   �?������W���8��*}�2I��g�F�Ž
	^��N��P4�;���<&O=(+=~�%=ح=��<@2d<�P�:(�J�T-Լ����Q�b~{� ͍��ر�����hay��B�?���0�%<�D�<LM=歈=���=@2�=R�=j��=���=�G�=�o=L�=�?�;�6�]���b��-�&���Z��S��-m��X���%P���   �   d��������l|�O�\��6��j�"���
�_��袼X�<T��<4:=�I[=�9c=��T=��3=��=XJ�< 3�w���"�rv������\ɽ�Z轾��������(�]ӽ�ۨ�@�m�c�Ы��D�<�*=�-r=�H�= ��=�=PX�=���=v�d=t�=�	Z<x�v�{C����8����>&���L���n�/T��Z���   �   I���?���-�����h齏��ڋ@�T|��DK<�)=*$V=Á=E.�=���= `}=PQ=@�=d�< [��� �ֺq����-G�8�"\,��]>�YH� I���?���-�+ ��p�E"��<�@��y|��%K<(#=�V=���=�,�=�ߊ=�]}=�Q=��=��<�I���	 ���q������A�5�X,�Y>�QTH��   �   Z��9 �mӽ\Ԩ���m�pW�@\����<�*=j3r=,K�=��=��=|Y�=ε�=>�d=,�=@Z<X�v�T�C��"��_���:B&���L�(�n��V����/�������8r|�$�\�6�tn�`���`�_������j<�u�<t	:= F[=66c=��T=��3=F�=�I�< �빰q�� "��v�X�DWɽ�S�Q�������   �   ���Sy��B��&��Џ0��D%<�U�<^M=۰�=��=>4�=��=���=~��=H�=o=X�=P-�;�>�y�������&�<�Z��U���o�����S���B������Z��;���"}�I�k���Ž�^�]����;��<�J=�+=f�%=P�=��<h.d<@U�:0�J�'Լ���Q��u{��Ǎ�0얽g����   �    �ɼP�x� �A��=<X �<l5=RTw=M��=D��=�F�=V>�=�m�=j��=���=���=��p=@,=@�ẾF/�շ�����S�UH�����nþ|�ؾ�}�̨꾭��־�k���?��&.����I�����1���B�(}�0_�;$��<���<h�<ܰ�<X�<P< �*����pU��<aǼ���>Q	��R��k�t����   �    @<��<@� =4�4=��k=���=���=���=�=Z��=�G�=h��=F��=~��=���=�Ll=@m�<��;�F�p�0뽬27�8�hꤾ}:ɾ�龂����	�\��@	�D� ��O羆�ƾ����F�|�:�8�2���ח�t��x�7����;(�]<��~<�V<� <�6�:Љ��x� ���Z��9x�2y�h|^���(�������:�   �   l�=2�9=,�g=3Ջ=h��=f��=���=���=��=�=^�=�
�=8�=Dx�=+�=��d=ě�<�#���$��w��^�U�^����佾����8{�/���� �>��T�	i��I�2꽾E$����]������ǽ�;g��(߼0�� ~�:0͌; �<;����0��������D���F��d$�0��� dǸ0z�; G|<���<�   �   �pR=�F�=�0�=짭=_0�=�)�=���=�k�=�>S�>&�>�	�=y�=b��=$�=U\=<���v���`.�8�n�����%�Ѿ���އ�rs#�)�-��1���-�mG#��p�Q=��]cӾy��?"{�v2�C���F����"�8���h��O���ﱻ�����E�؀m��vr��uL�@�� ��0�<hF�<t�<�l$=�   �    �y=���=���=VU�=f��=x��=Ԙ�=�>ld>pF>�>>
��=Vr�=���=>0V=�g<`��e7��B*���~�+���޾b��H�U-���7�J�;���7��-��q����,�t�����A�����Х��dC�Uؼ�Vs� �,��E2��w]��2��H~������X� Iػ c;�S<�u�<H�=��H=�   �   �C�=1V�=�?�=���=���=�]�=�v�=�+>�(>S�	>X3>Q�>���=���=�s�=b�S=��T<����ǽV9.�f4�������6���	�zN��c0��Z;�T?�GW;��n0����4c
���1����.��дF������T�N�H���@��xqM�@lQ�00z�д���n��X����`]� �л��M;�.k<h��<�� =�]T=�   �   ־y=ڭ�=ē�=~U�=���=���=��=�>zd>F>�>0>R��=�r�=J��=�1V=H�g<����5��*��~�4����޾���G�}-���7�a�;���7�-��p����*�s���,򆾮�A�����Υ��aC��Oؼ�Ls�hv,��;2��m]��-��Xy��<�� X��8ػ��;H�S<�x�<Z�=��H=�   �   rR=rG�=1�=:��=�0�=�)�=���=�k�=>o�>K�>,
�=�y�=��=%�=�W\=�ɍ<P��񁰽,�A�n�������Ѿh���c���q#�w�-�+1��-��E#�/o��:��aӾ���{��s2�,��C��>�"�����(���)��pʱ�ػ��E�8nm��dr��dL����� �P�<�K�<�	�<Zn$=�   �   D�=��9=D�g=�Ջ=���=���=ʻ�=��=��=V�=��=4�=�8�=Ny�=��=��d=���<��� ��G��H�U�є���὾Q�����x����"� �����f�F�罾�!��^�]�L��*�ǽ,2g�p߼`��@U�:��;�=;�ĉ�PP�����h�D���F��N$�P���  �����;�R|<X��<�   �   �H<�<�� =2�4=��k=U��=
��=��=b�=���=dH�=��=0��=���=m��=�Ql=dz�<8�;���p����-7�"��椾26ɾ��ݔ���	�;Y��=	��� ��J�)�ƾ8�����|�
�8����ї���p�7�@�;�^<��~<P:V<�<@4�:pK��hn �X�Z��x��y�ph^�؋(����@=�:�   �   |�ɼ �x� �A�H�=<"�<05=Uw=���=���=G�=�>�=�n�=k��=��=���=��p=z3= ���9/��������S�`D��y
���iþ��ؾ�w澬�꾥��[־�f���:��*����I���q(���B� �|���;\ȫ<���<��<D��<���<<<��(�Ȃ�F��SǼ����K	�N�"h�d}���   �   � �� Ry��B��$��x�0��G%<�V�<M=9��=���=�4�=��=���=�=J�=|o=��=p|�;�$������|�&�O�Z�NQ��vj��k���M���<������T���5��H}���H�.d�;�Ž�]�4>��m�;\��<�T=�+=n�%=>�=�(�<�Qd<�i�:��J�hԼ��^�P�4p{��ō�Qꖽ���   �   ���d��ӽ�Ө�*�m��V�W��D�<T*=F4r=�K�=���=��=�Z�=���=��d=`�=p)Z<H�v�<pC�u��ޔ���:&���L�R�n�bQ��n��l�������hg|�*�\�+�5��f�<���r�_�<բ� �<T��<n:=�O[=T?c=��T=R�3=�=�Z�< x繠a���	"��v�R𣽭Tɽ�Q轗������   �   � I�b�?���-�����h�D��H�@��Q|��GK<\*=.%V=�Á=2/�=@�=�c}=@Q=��=&�<@���$���X�q��}���9�0�TS,��S>� OH���H�v�?���-�8���`�?��B@�H)|��hK<41=�*V=Ɓ=1�=��=,f}=�Q=��=x%�<p��x �Эq������>��3�*W,�NX>��SH��   �   4��������l|�)�\��6��j�������_�h碼`�<8��<n:=�K[=�;c=��T=�3=f�=�Y�< �L]���"��v�0죽hOɽzK�]���&�������ҽQ̨�x~m��J������<�*=H:r=2N�=�¢=A�=,\�=���=��d=��=p%Z<`�v��tC���������=&���L���n��S�����   �   �?������W��r8��}�I��g��Ž�^��M���:�;���<~P=
+=(�%=��=�$�<�Ld<@b�:��J�<Լ���$�P�h{������䖽����;����Dy��rB����8_0�p%<dh�<|M=V��=��=�6�=` �=��=���=�J�=o=^�=0o�;H+㼴�������&���Z�\S���l������O���   �   ��꾩��?־Si��X=��0,��7�I����$-��2B��|����;|��<@��< �<`��<��<�4<�)�P��DC���MǼ0���E	��F�l_�8j���ɼH�x� A�x�=<4�<:5=\w=��=$��="I�=�@�=�o�=~��=ތ�=��=��p=�2=� ẜ=/�S�������
S�F�����1lþ��ؾ�z��   �   �Z�2?	��� �SM�l�ƾ1���F�|�ü8�+���ԗ������7�pȪ;h�]<��~</V<�<@��:�V���p ���Z�Px��y�0X^�w(��W��@�:�f<�.�<B� =��4=f�k=m��=���=T��=T�=^��=�I�=$��=��=L��=���=�Ql=|x�<��;��p�A뽯/7���V褾%8ɾZ��!���	��   �   U� ���<�
h�H澸轾	#����]�+��-�ǽ7g�� ߼�� ��:��;��<;@���_��h����D�@�F�(L$�p��� Թ� ��;�c|<���<��=�9=��g=>؋=2��=쭺=ý�=���=^�=��=���= �=p9�=�y�=��=X�d=ؤ�<����!��i����U�ߕ��㽾�����z�����   �   1�ˇ-��F#��o�<��RbӾ���� {��t2�u��qE��6�"���� ���9���ر����ТE��rm�Hhr�@fL�p��� ����<�O�<��<Pq$=RuR="I�=�2�=橭=22�=B+�=��=
m�=~>��>��>�
�=z�=`��=6%�=�W\=�ȍ<��������,�^�n�p�����Ѿ�������r#�J�-��   �   ֈ;�E�7��-�Gq�h���+�����򆾀�A�n���ϥ�ncC��Rؼ�Qs��z,��?2��q]��/���z��8��@X��9ػ �;p�S<Pz�<z�=ҢH=N�y=���=���=JV�=J��=L��=���=>�d>�F>�>V>���=�r�=a��=�1V=؉g<���5��^*���~����.�޾��PH��-�R�7��   �   vJ��w�/@��nʾ3,���]��$�a�)C*�H������!󁽚�R��9H��>\���/	��큰�����lƽ�E���ܭ�3����V�
0�����I<�=��V=q-�=��=��=�a�=4(�=U�>D�>pe>^�>�t><>>/ >��=B�=G��=>B<=p<)<R��o��� ����R�2���(��֨ɾ����   �   ^��?�4�ܾ�'ƾqZ������\�F�%����cA��,�w�AG��#=�B�P�(Ox�F퓽�B��*Y�������'������ �����R��= �@�"�P�:<�==r�O=��=���=�D�=�'�=(0�=u">q >�
>��>�f>w4>���=���=�6�=�Q�=rG==�5<~!��_��l:�V6N��U��m�����ž��ܾ�P��   �   ��d&ݾ,(ϾR����G���q��`�K������ؽrr��"�T��P&�v��L#0�AV��D��XM��1������k���9՝��+���I� L����:��A<�E�<8�9=X-}=�W�=k�=LF�=� �=�E�=�8>5�>W�>�'>Le>P�=t��=���=�A�=�?=��W<@u�06�����QA����*�������ŘϾrݾ�   �   ̾`=Ǿ;���r���	����f��Q2��j�����2�n���P��kԼ�|��4.!���M�ʂy��ݍ��(���Ж�o����r�:>�����0'p��j;���<��=*Q=�R�=���=�0�=v��=З�=���=@��=�X>�>���=���=p��=�[�=饔=<�A=�u�<p��Ş��̍�L�-�I�f��=�����������Ǿ�   �   +5������ԟ����_sp��@�J���Dνwd��@"�����ȇ@� �%��*m��A��t�	�LJ5��Z�`>r�~�z��2r���Z�ؾ6��w	��ƫ� ��`W�;`��<0�=�kH=�C�=j	�=�ȳ=���=���=���=l!�=���=�o�=���=�/�=��=`h�=��?=�8�<��{�*�_� ʽ����G��?x�E����u������   �   �B��،�L���oe��i?��.�G�ڽ�I��$~#�l����� ��;x2<��l;`N����w���ռ�� �3�G�f�N��I�^+:��!�PF�� ���F� �ʹ��J<4a�<*�$=~_=��==�=�4�=\��=���=���=V��=8d�=���='S�=YX�=f�7=8I�<�J!���2�dF������A&���N�U�q����� ���   �   �Sc��Z���G��-���ycӽD��l^��QQ����;\��<ؐ�<���<���<xgh<�i;P�����H$�����5�^�F�;O��|O�R2G�v�5����@0����� �|��0:<��<X3=��q=F�=�=ɺ=�e�=�0�=��= ��= Ȗ=��p=�c%=�J�<�uԻ��}˅��Ƚbp�7%���@��^U�sa��   �    "'�8*�.��	'�󰶽(�x�v�`�뻸9i<`��<�7(=^<=�:=X�&=>=�<��	<��<����@����,�,5W� :{�f��������^���������| b�h1)��4ȼ`��Ȅa<��=��I=&E�=�'�=���=\g�= ~�=�`�=��=h I=x�=� k<�4ѻ���X�U����Fн�C�����P� �X�'��   �   U(⽑Ͻ�ʰ��Y��D~7��z���e�:�<�9#=h�X=�fz=��=�f�=fl=��F=2p=�a�<0B�;��'�tiἴH8�p�~����D����cս�z��3��.�Ͻ%Ѱ�u_���7�썮��W�:���<�3#=�X=�az=Y�=�d�=Hl=��F=�l=�[�<�.�;�'�xi�G8�Ԣ~�@���o���4_ս_u��-��   �   ����|b��&)�L ȼ�Ҹ�H�a<= �I=�G�=**�=8��=gi�=��=�b�=��=8#I=� =&k<�2ѻ��X�फ़�UJнjH��n���� ���'��%'��-�����-����x����/컠i<t��<H2(=Y<=L�:=��&=��=l٬<�	<������ C��|�,�3W�46{�����ơ��cZ�������   �   ������A|�hR:<D��<b#3=��q=��=n�=.˺=og�=�2�=V��=���==ɖ=��p=�d%=�K�<�{Ի\���ͅ��Ƚr��%�щ@�dbU��va��Wc��Z���G�$-�8���hӽ�H��|f��mQ���;P��<���<��<���<�Sh< oi;`*������*������5���F��8O��xO��,G���5�����   �    �ǹ�K<o�<��$=��_=e�=��=&7�=Z��=^��=n��=���=pe�=���=T�=�X�= �7=�H�<8Q!���2��H��m���*D&�r�N���q�����"���D��ڌ��M��0se�m?�L1���ڽ�M����#�4"��@���0��;�<@>l;v��X�w�H�ռl����3���G�4�N�b�I�d*:���!�~B�����E��   �    ��<^�=2qH=�F�=��=˳=���=V��= ��=�"�=���=�p�=���=�0�=^�=�h�=��?=<7�<��{���_��ʽW��V�G��Bx�ٜ���w��t	��7��즫��֟����=vp���@�f��PHν�g���'�\��0�@���%��<m�K��,�	��N5�0Z�JBr���z��4r���Z���6�Fv	�����0���y�;�   �   �=�Q=�T�=���=P2�=��=J��=���=j��=KY>��>���=>��=���=\�=	��=�A=`s�<���j���-���-�G�f��>��������{�Ǿ�̾�>Ǿ�<��?t���
����f��S2�l������n�����`sԼ����22!��M�Ԇy��ߍ�P*��Җ�����D�r�d:>�����P!p���;��<�   �   f�9=�/}=�X�=���=rG�=�!�=�F�=V9>��>��>(>�e>��=���=��=�A�=l�?=0�W<�xἌ7����,SA�`����������Ͼ7sݾ�⾆'ݾ=)ϾH����H��Fr����K� ��S�ؽ�s����T��S&�,��&0�
DV�NF���N������$������֝�A,��\�I��K��0�:�PG<tI�<�   �   ��O=��=`��=LE�=>(�=�0�=�">� >5�
>�>�f>�4>��=���=�6�=�Q�=�F==��5<�"��`��;�7N�V��󮨾E�ž6�ܾBQ뾤^�h@뾼�ܾ(ƾ�Z����j\���%�r��B����w�nBG�%=���P��Px��C���Y��;���?(�����<�����R��= �(�"�X�:<�>=�   �   ��V=�-�=��=���=�a�=<(�=V�>H�>qe>]�>�t>6>;/ >t�=(�=$��=�A<=�:)<�������-���R�2���(���ɾ���vJ��o� @��nʾ ,���]����a�C*�������󁽌�R�:H��>\� ��<	����������lƽ�E���ܭ������V��/������I<P�=�   �   ��O=��=���=�E�=p(�=�0�=�">� >H�
>�>g>�4>J��=(��=:7�=\R�=|H==��5< �_���9��5N�FU�� ���3�ž
�ܾP�_]�*?뾌�ܾ�&ƾ�Y��>���\���%�d��W@��h�w�h?G�"=���P�vMx�^쓽�A��X��b���l&��P���������R�T; ���"� �:<H@=�   �   j�9=R1}=�Y�=��=�G�=�!�=(G�=t9>��>��>$(>�e> 	�=N �=��=�B�=T�?=��W<�n�L4�����PA����B���������Ͼ�pݾd�)%ݾ�&Ͼ5����F���p����K����h�ؽ�p��ڃT��M&�r��2 0��=V�C��gK������������ҝ�>)����I�lB���u:�T<�N�<�   �   ��="Q=~U�=l��=�2�=���=���=,��=���=vY>��>4��=܋�=���=*]�=���=�A=~�<����囆�q��T�-��f�`<��:���t���;�ǾP�˾�;Ǿ}9��bq��^��A�f��O2��h������n�\��
�\cԼ�s��~)!���M�@}y��ڍ�b%��Q͖�����r��2>������p� �;�
�<�   �   �ũ<��="sH=HG�=i�={˳=���=���=���=0#�=,��=Dq�=d��=�1�=��=�j�=��?=,D�<��{���_���ɽ��>�G��<x������s�����!3������ҟ�0��(pp�<�@�����@ν�`����쫼�r@�8o%��m� 6��0�	�lC5�pZ��6r�@z� *r���Z�ܵ6��n	�̴���󻀛�;�   �    �Ź�&K<hs�<~�$=�_=��=B�=�7�=ļ�=̈�=���=`��=Cf�=��=�U�=�Z�=`�7=�V�<H,!���2�hA��B����>&�~N�l�q��������\@���Ռ��I���ke��f?��+���ڽ.E��fv#����@J�� �;�I<��l;���@�w�X�ռ���$�3��uG�z�N���I�� :�P�!�x;�(����E��   �   ��<����|� Y:<̑�<b$3=��q=s��=��=�˺=�g�=J3�=.��=���=�ʖ=µp=�j%=TZ�<0ԻT��ƅ��Ƚ�l�|%���@��ZU��na��Oc���Z���G��	-����R]ӽ�>��>U� 2Q����;$ţ< ��<D��<LǷ<Ђh< 4j;x���t����H����5�̘F�/O�JpO��%G���5�����   �   �����b��$)�0ȼ�ȸ�h�a<�=��I=aH�=�*�=���=j�=ـ�=�c�==:'I==Bk<��л��LvX�����?нK<�����"� ��'��'�&�0����I���L�x�2�����Xi<,��<�=(=4d<=0;=��&=0=4�< �	<����,����*���,��(W��,{�����k����W��T����   �   �&�^Ͻ�ɰ��X��2}7��x���|�:��<�:#=@�X=�gz=?�=�g�=vl=X�F=�s=�k�<�u�;(c'�`TἎ;8�p�~�����Lｽ�Wս�m��%�h ��	Ͻ{ð��R��r7��d�����:��<4A#=��X=�lz=��=�i�=�!l=R�F=�w=hr�<��;`\'�pSἬ<8�b�~�
�����1\ս�r��+��   �   z!'��)�̅�u&�}���`�x�����뻀<i<���<�8(=0_<=j�:="�&=�=��<ذ	<�š�����.��R�,�0'W��){�Ɤ�隔�_S��p��������b��)�|ȼ0|����a<�=|�I=FK�= -�=��=l�=ł�=�e�=�=8*I=�= Ik<��л\�켦xX�7���Cн�@��N��B� ���'��   �   |Sc���Z���G�l-���&cӽ�C���]��OQ����;ع�<���<D��<���<�oh< �i;�	�P}��������5���F�L-O��lO�� G�\�5�`���̇��@�{��z:<���<�+3=8�q=D��=L�=�ͺ=�i�=5�=���=.­=̖=
�p=,l%= \�<�1Ի����ǅ�UȽ�n��%���@��]U�lra��   �   bB���׌��K���oe��i?�v.�
�ڽqI���}#�P��@���@��; 6< �l;`A��؟w�زռ&��2�3��xG���N���I�N :�f�!�.8����`�E� �¹�AK< ��<*�$=P�_=��=��=�9�=ɾ�=���=���=���=�g�=@��=�V�=�[�=h�7=,W�<�/!�@�2�cC��:����@&���N���q�h�������   �   
5�������ԟ����Esp���@�2���DνDd���!�������@��%��&m�0?��Ɗ	�H5��
Z��:r���z��,r�L�Z�\�6��m	����0��@��;�Ω<��=,xH=�I�=��=�ͳ=��=z��=��=�$�=h��=hr�=h��=p2�=w�=k�=`�?=�C�<��{�>�_���ɽ���1�G�8?x������u��j���   �   � ̾Q=Ǿ;���r���	����f��Q2��j�v����n���x��jԼ`{��X-!���M�8�y��܍�6'���Ζ�O�����r��3>�����p� �;��<��=R%Q=:W�=0��=�4�=��=��=n��=ص�=�Y>,�>���=���=f��=�]�=䧔=6�A=T}�<�������4�콘�-���f�l=��z���������Ǿ�   �   ��]&ݾ&(ϾM����G���q��T�K������ؽVr���T��P&����"0��@V�kD���L���������T����ӝ�*���I�C��xt:��W<PQ�<"�9=J3}=�Z�=2��=�H�=�"�=H�=�9>�>�>o(>�e>�	�=� �=>��=3C�=n�?=`�W<xp�5�����~QA�j�����~�����Ͼ�qݾ�   �   ^��?�1�ܾ�'ƾoZ������\�@�%����WA���w��@G�j#=��P��Nx�퓽�B���X��#���!'��쪩�)�����R��; �`�"���:<�@=`�O=s �=*��=F�=�(�=T1�=�">� >q�
>�>$g>�4>���=`��=n7�=�R�=�H==Х5<N �b_��0:� 6N��U��[�����ž��ܾ�P��   �   �l�����@���2�j�H���#���w�Ƚ䠟�m����{��ud���Oý�i����ˊ0��G�2V���[��V��*F�|Y-�����Fսv��x	� lp��/�<�\=��=�B�=��=Rs�=+4>mq
>�>�\>w3>�v
>d�>_�=.��=]��=fی=fl1=p+V<(i���Iz���ӽ�����A��"h��J��{���   �   |>��?퉾���Ne���B��������h����E]���I���䗽�<�����0]���+�\B���P�KcV�5Q�y�A��)�X�
���н�C���b���e�Pz�<�fY=Θ= ��=<��=���=\�>R1	>u�>�;>�>�X	>��>�)�=���=@�=s��=V0= #X<Ա����t��TϽpa��=�l@c��~��g���   �   ��������o�2�T���3�B����⽣�����(�d�"}d�����Щ����ս������|3��B���G��5C��25��������Ľੁ�G��@q��L��<��N=�ڑ=��=���=ք�=t��=�e>�S	>�
>�	>��>µ�=Xn�=�}�= H�=�0�=tN+=0�Z<X���h�d���½$l
��	2��5U���p�:���   �   ��k��e�<T�|�:�9��!����载�ዽ�P�b�+�Z�+�j�N�n��4C���W⽎��5����*�_�0�h�-�f"����������x}n��r�Y�p�<�C:=Ne�=0�=Re�=�c�=�.�=8��=@>"�>8�>� >t��=T��=�Q�=�7�=.~=2!=@S<�ь���N�����H��r{ ���?�;X��qg��   �   �H�"�A���1�\���K����Ľ����-D�z ��OƼ,&Ƽ�j���<����������۽�� ��!�`��N~���
�����^ν�L���CZ�H�����Hǌ<�=D_d=#h�=�Q�=4��=f`�=&��=�F�=�"�=jo�=`�=���=5��=��=)��=��c=�;=��1<<����48�� ���qڽ~V�
�%���9���E��   �   �!�����x콟ɻ�C8����3��ɼ�>2� �z� d{���-�ȷ��L�#�tq��̟��~½��ܽ��� ,��Ͻ�p���荽�N�t��H;8����;���<Nq-=Em=���=�߬=���=���=�u�= �=���=*�=F��=J'�=Z�=���=�b<=��<��;����`t(��ȇ��溽n�꽜�	����&C!��   �    .���!��rǽxȡ���m�V������ @�6�RA<�$�<���<`'B< &k:�Xb�Xd���WD�&���T㜽l���Ʃ�����Ԫ��~���ς�R�P�(��ȴ�І޻P�<�{�<p�!=��\=�X�=wl�=���=�=k�=nQ�= u�=3-�=8�=�=��E=�=�	}<��(�<Ԯ�l&��t�����½�ݽ8�q���   �   }۫��>��Zix�~�3� eϼЪۻ�+*<���<�<=j�!=�^!=�5=�P�<X�@<��V� ��(���B���l�����ތ�\X��N7��HD���=h��cF�L_�<�ڼ�$]� :<��<�� =��;=Lp=y�=qJ�=I�=�|�=)�=آ�=�nh=vE4=`��<�Co<��E�i��h����z6���k����K��ƪ�����D���   �   �2W�<)��@5@�p��;��<�=�{C=D�e=
�v=.�u=-c=��@=��=���<0;�;p1���~�������8�<�\�z�x����� I���؋����n�x��:W�"D)�h"��T@��u�;��<��=�uC=̽e=��v=��u=�'c=,�@=��=$��<��;pd����������8�.�\���x������G��֋� ����x��   �   ��ڼ�	]� `�:ȹ�<2� =�<=�p=�=�L�=hK�=�=��=S��=�sh=�J4=$��<hXo< �D�a�������y6��k�����L������A��` ���߫�0C���rx�D�3��uϼ��ۻ *<(��<�6=��!=�X!=0=8D�<��@<@W�� ����� B�R�l�^	�������Y���7���C��;h��_F�Z��   �   �a޻h�<���<��!=
�\=4[�=�n�=ք�=��=m�=rS�= w�=G/�=]�=3�=غE=�=p}<�{(�,Ѯ�X&�n�t�����½� ޽2<�>v���2���&��wǽ͡�*�m� ����� ���:A<$�<舑<PB< �i:�tb�Ds���_D�,���N眽-����������֪����=Ђ�<�P���\����   �   p��;��<�u-=jIm=��=��=���=���=�w�=�!�=H��=�+�=��=�(�=�[�=��=�e<=���<���;����bu(�	ʇ��躽X��v�	�����E!�n�!�v!���0}��ͻ�<����3���ɼ�U2� �z���{��-��Ľ�8�#��{q��П���½��ܽ��뽰/��� ϽFr��Z鍽�N��q��`18��   �   �ˌ<��=jbd=�i�=�S�=Ȼ�=�a�=���=�G�=�#�=�p�=��=��={��=Y��=K��=��c=�<=8�1<ၼ@68�m���sڽ�W��%���9���E�V�H���A��1�����O���Ľ���63D��%�ZƼx0Ƽ�o�z�<����*�����۽� ��#�E����n�
�m���{`ν�M���DZ�h��0���   �   T�<�E:=hf�=\�=|f�=�d�=�/�=@��=�>��>��>= >f��=0��=|R�=�8�=4/~=�!=@S<4ӌ���N�o���o���| ���?��<X��sg���k��e�6T�N�:�ڰ����5뽽K䋽D�P���+���+��N��p���E���Z�.�����d�*��0���-��"����������v~n��r��L��   �   $��<�N=�ۑ=N�=���=���=.��=�e>�S	>Q�
>>�	>�>T��=�n�=~�=�H�=>1�=�N+=�Z<L���"�d�˞½�l
�2�	7U��p��:�����Կ��a�o�}�T���3�F��z��D������0�d�D�d�:���������ս����}3��B�3�G�7C��35����.��y�ĽH���TG���b���   �   �{�<\gY=wΘ=l��=���=��=��>~1	>��>�;>">Y	>��>*�=��=_�=��=60=�!X<l�����t��UϽ�a���=�"Ac�2������>���퉾y����e�&�B�z�����Pi�����^��{J���嗽�=��ݔ��]���+�B�T Q��cV��5Q���A�p�)���
���н	D���b���e��   �   `0�<R�\=��=�B�=.��=\s�=14>rq
>�>�\>x3>�v
>a�> _�=$��=C��=Eی=l1=�)V<j��:Jz���ӽ���ǫA��"h��J��}���l�����;����j�H���#���X�Ƚࠟ�o����{���d�� Pý�i����ފ0��G� 2V���[��V��*F�fY-����xFս9��	��Tp��   �   �~�<�hY=�Θ=¸�=���=D��=��>�1	>��>�;>6>Y	>�>H*�=Z��=��=��=�0=�(X<����t��SϽ�`�r�=��?c�j~�����>���쉾����{e���B�J�����ug��-��o\���H��䗽�;��ʒ콨\�d�+��B���P��bV�14Q���A�:�)���
��н|B��f`� e��   �   ��<4�N=oܑ=��= ��=���=x��=f>
T	>m�
>]�	>D�>���=Xo�=�~�=TI�=O2�=bQ+= �Z<@���n�d�H�½�j
��2�N4U��p�G9��"��=���Y�o���T�c�3���y�⽱���[����d�zd����������ս�����/{3�B�|�G�\4C�015����%���ĽY����=���為�   �   ���<�H:=�g�=J�=2g�=de�="0�=���=�>��>��>p >���=���=RS�=�9�=$2~=�!=8/S<�ƌ���N������ ��py ���?��8X�Hog�q�k��e�
T�f�:�R�������彽Pߋ� �P���+���+��{N��k��q@���T����T����*�F�0�D�-�@"�������:�Vvn�te�`���   �   �Ռ<��=Ped=�j�=VT�=f��=db�=���=JH�=L$�=q�= �=���=B��=`��=���=l�c=�A= �1<�с��,8�����mڽ�S�^�%���9���E��H�T�A���1���G����Ľ��2'D����DƼXƼ�d�|�<�V ��ߡ����۽�� �n�Ь��{�N�
������Yν�G���:Z����Pܢ��   �    ��;(�<�x-=�Km=���=��=<��=��=�w�=$"�=¹�=D,�=���=�)�=�\�=���=�i<=��<@�;,p��k(��Ç�{ẽ��꽚�	�����?!���!���%�s콳Ļ��3��ҿ3� |ɼ%2� ?z�`{�0�-� ���#��kq�ȟ�zy½L�ܽ$��E&����Ͻ�j��㍽
�M�H`���8��   �   �5޻�<x��<j�!=��\=�[�=jo�=Z��=z��=�m�=�S�=�w�=�/�=A�=_�=�E=�
=`,}< (�D����&���t�2���_½�ݽ�1�k��{'��G��lǽ�¡���m�L��T �77�mA<l1�<<��< BB<��l:h9b��R��ND�ݕ���ݜ�v�����������Ϊ�ix���ɂ���P���L����   �   d�ڼh�\��:h��<� =X<=�p=��=UM�=�K�=��=�=���=�uh=M4=��<�go< DC�(T��\���xo6���k��~���D��C���#�����ի�_8���]x���3��Qϼ dۻ K*<���<:C=�"=�d!=x<=�^�<�A<�V���������B�̴l�V ��W،��Q���0���=���0h�DWF�PS��   �   .W�R8)����,@�`��;\�<��=�|C=�e=��v=�u=.c=�@=d�=쪳< Q�;���8u�����T�8��\�V�x�b�vA��Ћ�����x��&W�l0)�@��@�P��;P�<`�=��C=��e=�v=@�u=^3c=��@=.�=8��<��;p����h������8���\���x�S�YB���ы�7��x�x��   �   j٫��<���fx���3�`bϼ��ۻ /*<@��<l==8�!=n_!=�6=�R�<�@<@zV�H�����B���l�T���ڌ��S���1���=���.h��SF�zN���ڼ��\� ��:�˄<t� =l<=�p=�=�O�=0N�=܁�=v�=p��=�zh=RR4=̟�<8}o< B��K��Č��vm6�D�k�{��?F��̦��s������   �   P,��O ��qǽ�ǡ�n�m�h������  �6�UA<&�<앑<�*B<�bk:Tb�4a���UD�י���᜽E����������Ъ��y��sʂ��P���ج��p޻0<��<̐!=$�\=s^�=�q�=���=���=�o�=�U�=�y�=	2�=Z�=��=@�E=�=P;}<��'�H���&&���t������½+�ݽj5�zo���   �   <�!�h����w�0ɻ��7���3��ɼp<2���z��Z{���-�@���V�#��rq��˟��}½e�ܽ!���)�佊Ͻ�l��-䍽��M��^��8����;<�<�|-=�Om=��=��="��=���=�y�=�#�=`��=�-�=H��=�+�=�^�=H��=�l<=8��<��;Dn��Tk(��ć�3㺽G��K�	����LB!��   �   p�H�ĉA�[�1�*��BK��O�Ľt�� -D� �OƼ8%Ƽ�i��<�X��+���E�۽�� �d!�����}���
������[νDI��F<Z���꼐բ�0ٌ<��=hd=fl�=�U�=���=�c�=d��=�I�=�%�=`r�=f�=ֺ�=���=���=洖=��c=fC=��1<tс��-8������nڽKU��%���9���E��   �   }�k��e�T�W�:�������v载�ዽ��P��+���+�
�N��m���B��hW�Z�����X�*���0���-��"�����뽪���xn��f� ��T��<DJ:=�h�=L�=>h�=xf�=(1�=���=c >:�>P�>� >���=���=@T�=�:�=�3~=� !=�1S<�ƌ�N�����R���z �J�?��:X�5qg��   �   ������ށo� �T���3�2����⽂�������d��|d�i���������ս�����Z|3�WB���G��5C�I25������'�Ľ*���|?�� ������<�N=�ܑ=��=���=���=��=ff>XT	>��
>��	>��>J��=�o�=T�=�I�=�2�=R+=��Z<����B�d��½�k
�n	2�Z5U�V�p��9���   �   r>��6퉾���Ee���B�������vh����9]���I���䗽�<����� ]���+�JB���P�*cV��4Q�B�A�ɝ)��
���нC�� a��$e�h~�<�hY=Ϙ= ��=.��=���=��>�1	>��><>X>@Y	>0�>�*�=���="�=\��=&0=(*X<�����t��SϽ!a�ڠ=�7@c��~��V���   �   1Q�,o�������;�Ž]���u��(�v��2��� ����ɽ�M��Z2�o�b��{��H�������\���.0ž�����4�������釾d�X����G�ҽ�\��5.��W�<&?i=m�=�f�=��=�>�%	>�@>U�>�]>��	>��>>��=A�=���=kP�=�C�=NT1=��<���@"��x��챽2{�)f�F��   �   n��x��l� ��A⽄���|����[����j�^]t����m�½�&�4�-�W]��@�����R����ϼ�"���ռ�I~��?L������$T����.�ͽ�PV�P� ����<>�h=�{�=��=�=�� >Z)>50>�b>�>�d>�h>�+�=H��=�g�=���=L�=��,=���<�dŻ���j�s�fg����ܽLa �#���   �    ���E ��'뽊�̽;r��;ǉ�3a��RH�MQ��Ҁ�����k)�k���L�g�{����0W��D����+��;P��T˥�rɓ�z�V%G�Ǫ�mο�:�D� d��`��<�f=rn�=f��=��= 8�=0>x�>]�	>�>>�B�=f��= �=:��=��=\n=��=�[�<���]��uh�B�����νʃ�U���   �   �6轿޽�Ƚہ�� �����X�Hx)�4��-�j�F��ٌ�P`ȽHh	�rj3��^�T^���Ǔ�����¢�7���#R��\/��;ha�a3����#��B/+�`蕻t�<z�_=���=e��=�=�`�=���=�8>I�>�[> 1�=���=�f�=��=?��=ԍ�=�M=��= �@<�P�2� ���Y�{���b����սSe��   �   �����]���������PF�����Vļ�
���榼t����E��-��|�ڽ���9�p�]�V{����㲋��S��2Հ��>f�BC��a�J��I������d���<p�S=�ܓ=��=��=P��=J(�=.��=2l�=^9�=���=�~�=���=��=d�=T�Z=R`=L�<`uc;8-o�?��?N�����d��D�������   �   ��Nф���\�2&�$�ټ��a� 膻 @E: -�X���D˼�B�{e����ܽ�*���/���I��\��Bd���a�"�T�4�>�"���;̿�Ґx� ��I�����<N�==�(�=Iޤ=Pܽ=T�=Rb�=Z��=l��=�l�=�W�=�3�=eܜ=#R�=�8K=�N=���<Pʪ;�b���¼^R�j�L��x�┍�����y���   �   r�S�DO-�����`���0!�� :<xs�< ��<z�<P[< �6�)����1������^ʽ�[ ��S���'�T0�p00��'������XVԽ�[����S���ټ@"F�T��<�L=X�`=��=Џ�=�ж=�/�=v[�=H�=y5�=ʸ�=I��=�c=�,'=���<�".<��l������$�J��_@�T\�f�o��Lz��y�?m��   �   ~	�$߱�������;�$�<DS�<.e=�l+=��)=��=���<`U<��;�vo���m��M����ͽ� �_��B�� #���s�u�ͽ�'��%����2?�����N���<87�<��)=�ia=w�=\#�=*��=Z��=�+�=�͎=br=<P:=�G�<x�P<`m���⤼z���O:��O]��pt��3��P����z���j��qR��1��   �   N��P��� �*<�c�<X�=b�G=Z�h=d!{=�|=DPj=�E=\�=��< }߹H0���W#�^�j�D]��ަ�n���/������������޻p��I>����T���ߍ�0�*<(Z�<b�=|�G=p�h=t{=�|=�Jj=��E=��=Dڗ< ��(C���a#���j��b���㦽%���3��+����������p��H>�����   �   hE�x�<�>�<��)=�ma=8y�=�%�=^��=���=5.�=KЎ=\!r=�V:=�V�<�Q<@(��(Ѥ�����G:� H]��jt�N1�������z�F�j��sR���1� 	�h鱼�� q�;��<�H�<�_=�g+=�)=�=���<�7<p�;��x��m�@S����ͽ��e�����'���w齂�ͽ�)��<����2?�t���   �   �F�� �<�O=��`=;�=���=�Ҷ=�1�=r]�=:J�=�7�=X��=Č=�c=�3'=��<`?.< !l� �������2\@��\���o�pNz�d�y�hCm���S��T-�����X��� P���#<lh�<��<�n�<�f[< ���9����1��Ɛ��dʽ�^ �W��'�ZW0��30�ֽ'������XԽA]��2�S���ټ�   �   �;��\��<R�==�)�=�ߤ=�ݽ=��=�c�=���=(��=�n�=�Y�=6�=�ޜ=�T�=`>K=T=���< �;HS�L�¼�P�d�L���x�I������-|�����NԄ���\�@
&�ؐټ0 b�`�� �C:���8��(R˼��B��i����ܽ�-���/���I�J!\�Fd���a���T���>���"�W�Bο��x�����   �    g�t��<҃S={ݓ=��=��=t��=|)�=r��=�m�=�:�=j��=���=���=��=,f�=R�Z=
d=��<��c;8'o��>��@N����Kf��`��%���u���}`��㷝�֦���UF����l`ļh����h���:�E�1����ڽ�İ9�Z�]�7Y{�����w���bU���ր�OAf�0C�Nc�^�K������   �   �땻�<R�_=#��= �=��=�a�=j��=89>ȣ>\>J2�= �=<h�=T��=���=4��=LM=��=з@<XN�x� ��Y���������Ԧս�g�9�<޽l�Ƚ>���] ���X�`|)�:��1���F�;܌�McȽj	�rl3�&�^��_��Lɓ�{���FĢ�~���NS��_0���ia�Pb3����$���0+��   �   0f��ܖ�<f=�n�=��= �=�8�=|>��>��	>�>>`C�=H��=�=��=꧚=�n=�=�\�<0�廲]� wh�0�����νP��0��	���F ��)�H�̽�s���ȉ��5a��UH�$PQ�VԀ������+�Nl�C�L��{����+X��D ���,��)Q��-̥�-ʓ�Dz�D&G�r��MϿ�(�D��   �   � �(��<��h=!|�=��=P�=�� >~)>]0>�b>+>�d>�h>T,�=���=h�=���=`L�=^�,=̼�<�fŻ���P�s��g��D�ܽ�a ���������� ��B�O���>���C\��4�j�_t������½.'��-��W]�>A��(��ܤ��&м����ּ��~���L����*%T�Ί���ͽ�PV��   �   �3.��X�<|?i=0m�=�f�=*��=�>�%	>�@>W�>�]>��	>��>4��=A�=���=UP�=vC�=T1=0�<�����"�Hx��P{�4f�F�4Q�,o�������2�ŽW���u��@�v��2��� ��&�ɽ�M�
[2���b��{��W�������d���/0ž�����4�������釾:�X�x���ҽT�\��   �   0� ����<�h=�|�=R�=��=�� >�)>o0>�b>=>�d>�h>�,�=���=hh�=j��=�L�=��,=��< VŻ��f�s�Jf��[�ܽ�` ����͇�؄�Ҿ ��@�x��������Z���j��[t�R�����½&���-�jV]�f@��8��أ��ϼ�����Լ��}���K��6���#T������ͽNV��   �   �C��t��<�f=�o�=���=��=9�=�>��>��	>>�>�C�=���=x�=���=���=�n=��=8c�<�u��X�fqh�����,�ν\�������D ��%�n�̽Lp��rŉ��/a��OH�JQ�р����'��i�z�L���{�9���>V��@����*��&O��Eʥ�nȓ�0z��#G�@���˿���D��   �   0���\�<�`=q��=�=�	�=:b�=ܪ�=f9>�>?\>�2�=� �=�h�=���=���=F��=
M=8�=x�@<�8��� �N�Y�����_�ս�a�D3�g
޽ïȽ�~��h�����X��s)���L)���F�7׌��]Ƚ�f	��h3���^�]���Ɠ�����t��������P���-���ea��^3��� ���(+��   �   ���|��<�S=ߓ=+��=��=��=*�=���=�m�=>;�=���=>��=T��=Ҿ�=*g�=��Z=\g=0��<��c;o��6�07N���G`�����F���q����Y��"���u����IF����pKļ ��ܦ������E�.*����ڽh���9���]��R{�c������R��rӀ��;f�&C��^�%�FE������   �   @@�����<ܖ==�+�=��=�޽=��=vd�=���=���=Fo�=&Z�=�6�=�ߜ=�U�=�@K=�V=̽�< �;8<���¼FH�>�L���x�ŏ������t��P ���̄��\�J�%��vټX�a����� �F:������l7˼��B�$a����ܽ�'�T�/��I�)\��>d���a�H�T���>�L�"���vƿ�j�x�����   �   ��E� �<nT=�`=��=���=RӶ=|2�=�]�=�J�=D8�=޻�=�Č=R c=v5'=��<K.<��k�����輨x�vS@��\���o�NAz��y�^4m�L�S��E-������o���䁻�U<p��<ḫ<h��<��[< �7�����1�o���Yʽ`X �HP���'�"P0�n,0�$�'���T���OԽaU��b�S��ټ�   �   �&�`�<�G�<�)=tpa=0z�=E&�=�='��=�.�=�Ў=d"r=X:=|Y�<�Q<����ˤ���C:�fB]��ct�-�����~�z���j�fR� �1�.���˱�(���ߟ;�3�< a�<�k=s+=��)=f�=���<�t<p�;�\e��m�)G���~ͽ>��PW��R��1��l�'�ͽ� �������&?��l��   �   �?��������*<,j�<��=$�G=��h=�"{=�	|=Qj=��E=Z�=��< �޹-���U#���j��[��uܦ�����,��+��B	��|���l�p�@=>����9��`s��`�*<�s�<z�=��G=|�h=P'{=�|=dVj=��E=�=P��< �ڹ����K#�\�j�WV��Cצ����(��������ګ���p��=>�����   �   V	��ձ����0��;�(�<\V�<Zf=�m+=|�)=ֻ=T��<Y<��;�Vn�&�m��L����ͽJ��I]��(��I ��fp齓�ͽ(#��'����'?��k�h�x�<�N�<��)=xta=F|�=](�=��=Z��=1�=Tӎ=$(r=�^:=�g�<h-Q< Ӊ�ع��6���::��:]�(]t�*��/��ķz�Ĺj��gR�8�1��   �   R�S�JK-������{�����?<�u�<���<�{�< �[<  16((���1����e^ʽN[ �jS�<�'�dS0��/0���'�r�Z���RԽnW����S�\�ټ��E���<�V=��`=$�=B��=ն=H4�=�_�=�L�=v:�=M��=kǌ=\&c=<'=��<�g.<�sk�,�����s��O@��\���o��Bz���y�p8m��   �   ���τ�4�\�v&���ټ��a��ᆻ mE: �����C˼r�B�*e��E�ܽ�*�C�/�F�I�v\�2Bd�ʣa�<�T� �>�{�"�`
��ȿ���x����@G����<j�==�,�=�=�=��=�e�=��=H��=q�=&\�=�8�=�=LX�=FK=�\=�Ȥ<P=�;+�`�¼8F���L���x�됍��	��w���   �   ���e\�����^���OF�ҏ�\Uļ�	���妼������E�Q-��;�ڽ����9�<�]��U{�𩇾�����S���Ԁ�&>f�LC��`���G����������<��S=�ߓ=���=��=&��="+�=��=Do�=�<�=p��=���=8��=���=Di�=,�Z=hk=`�< !d;�o��5�Z7N�u����a����������   �   �5��޽O�Ƚa��������X��w)���.-��F�sٌ�!`Ƚ*h	�Tj3�^�C^���Ǔ�����¢�	����Q��/���ga�9`3�9���!���*+��ĕ���<`=Δ�=��=,
�=�b�=���=�9>j�>�\>�3�=��=j�=m��=��=đ�=�M=��=�@<�3�~� ���Y�꥖�;��� �ս�c��   �   ʫ��E �~'�I�̽r��ǉ��2a��RH��LQ��Ҁ�v���H)��j���L�V�{����"W��3����+��P��2˥�Eɓ��z��$G�5��+Ϳ�~�D�@M��`��<�f=�o�=ؿ�=�=�9�=�>*�>�	>g> >�D�=���=l�=���=���=�n= �=�e�< p��X��qh�����-�ν�������   �   H��Z��V� ��A�d���h���n[����j�<]t����_�½�&�,�-��V]��@�����L����ϼ���{ռ�:~��*L�����~$T�>����ͽZOV��� ����<��h=�|�=c�=��=�� >�)>�0>�b>d> e>i>�,�=f��=�h�=���=]M�=��,=|��<PRŻ����s��f��ڝܽa �����   �   �yO���G�,�4�@!��V�z� �V����H��R���߽�o"���a������2��\��[�E��L��P�G�|��6���⾋ǹ����� N�ɉ������l���<2g~=�{�=T��=N��=��>��	>�P>��	>�>>s� >j��=Κ�=pU�=�[�=�ۗ=��u=��7=��<�I<�I��t
���B�2�-��G��   �   ��G��L?�N[+�p������D�������=�.���Y2ؽ����\�v!��D����>��a����d<��
�s��d�/�޾�
������@�I�p;�G����1V����<�s=�B�=�0�= ��=�>\�>��	>�Y>�]>غ�=N&�=pg�=��=�Ƭ=�f�=d�k=b�.=<_�< �4<�R���֝��8��A)���@��   �   |&2�h�&�
��LF���ü�T���yּ�K��y��H½F��L�K��3���G���HҾ[���z��>��N�
R�������Ѿ"C����fq<�t��2eo�����H�<���=bX�=���=��=�m>�l>��>;�>~`�=и�=F��=8��= �=���=Q��=�FL=��=�g�<`��;�����������Ԫ��/��   �   ���I���мdי��[��9�P(s��"ռ�+?���T��32��qq��ך�9漾��۾����҆�Lk����2�����ܾw���ϧ�� zm�sg(���ҽ�H��Cg�w
=<$�=^�=��=Dj�=D��=�d�=J�=P��=($�=���=��=�t�=|W�=�K|=��H="�=�T�<��8< �D�HDC�D뱼|���I�����   �   L9ڼ������[��,Ļ hθ`�; ���&����*h��5½N���3J�����zۡ������Ӿ�h�(�羽g�S�վ���^���������L������8Y�`<;H�=��=W��=X��=|}�=��=>��=��=���=���=Jչ=���=��= Z=�7%=���<�˃<0�;���� <W��\���ּ����v� �Hi���   �   ����`� _	�H<�Rp<���<ܿ�<�~<@^ ����Fͅ�:ڽ����~R�{���i��CǮ�u������T�����.���*��x�^�SK)����;i����ڼ�+<�=֗~=��=P�=�M�=23�=�a�=ԕ�=5��=M��=ћ�=N/d=p)&=��<@�9<�ܲ�8�F� 0���S߼���b������.�������˼�   �   ��2� �:��A<g�<�J�<r>=�g	=���<X�f<�Lѻ���r���߽�� $H��|p�@����ȓ��~���e��j͍��W���Z�:p1��D����(�R�i��@�V<�?=�vq=�/�=��=�~�=��=�U�=�v�=���=:Hx=ָ4=�T�<@P�;8�)�=ؼFv"�*�J���d�^To���l��^�d.G�R>(��b�p����   �   0�޻�
<hR�<��=��3=��J=
<O=܎==M=�Q�<�i����P����ͽJ9� �,�� H��[��.d�ҕb�*�V��1B�� '�R��wͽ�U�����!�h�r<�X=$�Z= ǈ=u��=%��=�Ϥ=R��=i�=N�S=8�	=�WO<�%�l���`�b�����]�ƽ�yν%˽AԽ��Ψ� ��@j_�������   �   @�л�Z<4_�<lI9=Zg=�n�=b!�=e��=VGh=3=Ĝ�<`&&;h�ļ�`W�g����ܽ:����������<\�p�GJ�|ǽ,����O�@m伀�лxZ<8[�<�F9=.g=�l�=X�=��=�Ah=�3=���<`�%;X�ļ�lW��m��f�ܽ>����������_���ZO󽝀ǽ���R�O��p��   �   (!�X�r<�Y=�Z=eȈ=���=� �=�Ѥ=���=>�=��S=
=�|O<�%����*�`�������}�ƽsνN�ʽEϽ��ʨ����Df_���� �P�޻p�
<M�<R�=��3=��J=�7O=̉==*G=D�<�?j����hV����ͽ$=�b�,��H��[��3d�K�b�I�V��5B��'�����ͽ3X��f��   �   �l��P�V<z@= xq=�0�=��=`��=ʂ�=�W�=iy�=ҳ�=�Nx=��4=Df�<0��;�)��&ؼ�j"�,�J��vd�FKo�&�l��^�4*G��;(��a������2� O:ȯA<�_�<�B�<*:=c	=h��< �f< �ѻv���w��8�߽�	�(H�"�p�����~˓�,���2h���ύ��[�2�Z��r1��F������R��   �   ��ڼ�'<�=��~=��=D�=�N�=�4�=jc�=җ�=�¿=� �=힏=Z6d=21&=@�<�9<@Ʊ���F�� ��`F߼v��X��`��x-����X�˼@���X(��<
�<�Bp<Dؒ<���<�i<8v �����х�,?ڽ�����R�}��l���ɮ���������V�����4���,��A�^�tM)���Ak���   �   �[���;;�=��=؜�=
��=d~�=��=���=��=���=���=�׹=���=��=t�Z=:>%=��<؃<��;�x��P-W��W���ּ<���T� ��l��X>ڼ����(�[��IĻ ָ�G; 7���(&���鼨$h��9½���l6J�C���jݡ�,����Ӿ�j⾐��j�v�վs������+����L��������   �   H�H��Ug��v
=X$�=��=h��=�j�=��=�e�=j�=���=�%�=h��=���=�v�=�Y�=|P|=.�H=\�=P\�<ؘ8<�D��>C�0걼4��K���� ��L� �м�ݙ��[���9��6s��*ռ�0?����� X��52�Dtq��ؚ��缾��۾����؇�Rl��������r�ܾԣ�����{m��h(���ҽ�   �   �fo����lH�<���=�X�=���=���=�m>$m>��>��>xa�=���=���=���=�!�=h��=���=�IL=�=0k�<`��; �绬���ȟ����j�/�^(2�v�&�F���J�ü�Y���~ּ�N�.y�K½���سK�t4��I��
JҾ���{��?��O��R�4��,��ܙѾ�C��U�Hr<�����   �   ����@2V����<8t=�B�=�0�=`��=�>��>��	>�Y>^>j��=�&�=h�=���=�Ǭ=}g�=��k=T�.=�`�<��4<�Q��`ם�49��B)���@���G�N?�x\+����������P��<�=�4����3ؽ����	\�"������ྠ��������<��
����Zd���޾��������I��;��   �   \��Ⱥl���<�g~=�{�=r��=^��=��>��	>�P>��	>�>>t� >l��=̚�=fU�=o[�=�ۗ=\�u=��7=��<�I<�K���
��&C�`�-��G��yO���G�(�4�B!��V��� �|���H��R��8�߽�o"��a�ڍ��3��x��[�O��R��P�B�w��,�����pǹ�댏�y N�����   �   쉄��(V�<��<�u=>C�=P1�=���=�>��>��	>�Y>^>���='�=Fh�=���=�Ǭ=�g�=|�k=��.=dc�<P�4<@B���ҝ��6��?)���@���G�K?��Y+�ږ���������B�=������1ؽe��p\�!�����V���	��8��;�5
����c�t�޾	
�����H�I��:��   �   �`o� ��HO�<$��=�Y�=���=��=�m>Jm>�>ˀ>�a�=>��=Ԝ�=��=�!�=���=l��=PKL=D�=�p�<��;�a� ���(���¦���/��"2�؀&����(@��üxO��tּ(I��y�KG½H���K��2��G���GҾ!��&z�>�0N�FQ�Β���󾘗Ѿ�A���򃾺o<��}��   �   ��H�@�f�|{
=&�=��=b��=�k�=���=*f�=��=���=&�=ʡ�=^��=Rw�=XZ�=R|=&�H=��=`b�<��8<��B��)C�Pޱ�����C���4��D���м�Ι�@�Z�`�9��s��ռ�'?���Q��H12��oq�4֚��伾C�۾����΅�?j����%�����ܾ����B���rwm�0e(�+�ҽ�   �   xQ�@k<;��=��=f��=.��=>�=���=��=��=���="��="ع=��=��=�Z=@%=T�<�݃< 1�; U���W�K��|�ռ@����� ��Z���+ڼМ��x[�pĻ Pĸ �; ���(&�,��h��1½���0J�����١�퀽�r�Ӿf⾣��;e��վE��H��� �����L����ﯽ�   �   \�ڼ�I<T=T�~=@�=��=�O�=X5�=d�=H��= ÿ=t�=g��=z7d=�2&=|�<�9<�r����F�����<߼���t������$�H���l�˼ؙ���� ���-<�ip<��<�ʄ<��<XF ����;Ʌ�/5ڽ���x{R�
y��g���Į�Ν��H���VQ��������(��n�^��G)����d���   �   V�� �V<�F=�|q=F2�=�=T��=���=NX�=�y�=M��=�Ox=��4=�h�<`��;H�)��"ؼbh"���J��rd�RFo�0�l��^�J"G�3(�bX�h���@g2� �:h�A<Ht�<�V�<2D=jm	=���<�g<0ѻ���m���߽h��H��wp�����HƓ��{��c���ʍ��R�5�Z�l1�A�P�� �R��   �   �� ���r<<`=ȲZ= ʈ=B��=��=tҤ=O��=��=��S=
=��O<��%�B����`����������ƽ2qν��ʽo̽�3Ǩ�6���]_�����ٹ���޻�
<Da�<J�=��3=��J=�AO=��==TS=$`�<�6i����J���ͽ`5���,�(�G��[��)d���b��V�-B�F�&�:��-
ͽhO��h��   �   `5л�=Z<�j�<�M9=~g=�o�=?"�=��=nHh=�3=���<�4&;p�ļ�_W�xf���ܽ�9�d��"�����,[�,�DG�9yǽS����O�|[��:л�?Z<�m�<P9=V!g=�q�='$�=8��=bMh=�3=���< �&;��ļ�SW��_����ܽ�5�F�� �����}W����A��tǽ(��V�O��V��   �   0�޻ �
<�\�<F�=n�3=��J=�=O=�==�M=�S�<�i���-P��h�ͽ9�Ќ,�� H�j[�J.d��b�D�V��0B���&�֤�ͽ5R����x� �h�r<a=\�Z=9ˈ=���=��=_Ԥ=���=[�=�S=b
=(�O<��%�޼��s`����������ƽ�jν��ʽ"ǽ��¨��	��<Y_�����׹��   �   pl2��`:��A<lm�<(O�<(@=i	=���<��f<�Fѻ.��%r����߽���#H�S|p�����ȓ�j~��ze��͍��V���Z��n1�JC��
����R�X[��P�V<�F=�}q=3�="�=���=%��=1Z�=(|�=�=Vx=��4=ty�<��;��)��ؼ]"���J�hd��<o��l���^��G�0(�W������   �   ȝ��
����X<@Zp<��<���<��<x[ �0���̅��9ڽ����~R��z���i��#Ǯ�O���֣���S��f�����o*����^�:J)�$�꽝f���ڼ�B<�=��~=��=T�=�P�=�6�=�e�= ��=)ſ=�=c��=B>d=:&='�<��9<�X��XvF�`��,.߼���̋�n��*#�����p�˼�   �   0ڼ���� �[��Ļ �˸`�; ���(&���鼨h�X5½,��o3J�����hۡ�������Ӿgh��羕g��վL�����|�����L�������T��I<;ʥ=��=���=���=��=���=D��=Z�=���=&��=rڹ=���=s�=8�Z=�F%=��<��<�`�;P+�� W��D����ռ����.� ��]���   �   X�XG�D�м�ԙ��[���9�&s��!ռ|+?��񟽏T���22��qq�vך�,漾��۾����ʆ�Bk���������ܾ@��������ym��f(���ҽ�H� g�Tz
=�%�=�=���=l�=B��= g�=��=0��=x'�=v��=C��=ly�=�\�=�V|=��H=`�=�j�<�8<�DB��!C�Hܱ����D�����   �   j$2�Ђ&����D�ü�S���xּ�K�ry��H½8��<�K��3���G���HҾR���z��>��N�R�������ØѾ�B���� q<���@co�X��M�<���=|Y�=Μ�=P��=(n>�m>f�>2�>�b�=P��=��=L��=j#�={��==0NL=��=u�<@�;pX�,�������p��4�/��   �   ��G�*L?��Z+������������h�=����L2ؽ����\�q!��?����<��^����c<��
�m��d��޾�
�������I�8;�ʊ���-V����<u= C�=T1�=���=�>��>�	>Z>U^>��=�'�=�h�=���=�Ȭ=�h�=��k=��.=�e�<�4< =��8ҝ��6�J@)�v�@��   �   �<��$<��(<0<`�c;(���q�Ny�g�۽�d.�1���n����|���.�B�H�(Y]���j�H"o���j��-]�^fH��".������侘���U�l�HU�4����s3�TI=�؍=b�=�=H��=?�>!�>)>��=|d�=j1�=���=�Y�=��=-��='�=��e=@=��= ��<@ʹ<�܉<�nO<آ)<�   �   Ha'<`�3< �<<�)(<�̩;��Ȼ�J׼Ԉm��Խ��)��Az����$F�9�+�E�MBY�}Jf���j��Bf��$Y�z�D�P�*�}��`qྈk����g�̄��n��`���=���=�D�=(0�=�"�=��>�>;>��=��=���=��=Ƒ�=��=T�=�#|=�V=�_2=f'= ��<��<��<��G<�h*<�   �   H�<<��[< ft<��l< e%< �ѹ�����HK���B���zh��K���X־5��n�!��:��bM�:�Y��&^�F�Y�,lM�K�9�q!�H��R`Ӿ�1��fAX�:����t��ՙ���==d��=L�=
�=`!�=��=(�=�2�=�w�=���=�ŵ=V۠=�=�(p=��J=��'=�=�v�<��< -�<�OI<��+<H)<�   �   ��T<l݉<��<���<h}�<X�<�#�N��G������L�����:���)W�G��|)���:�/`F�{jJ���F�� ;�\L)�������$��5g���@��d�*qG� �;x�+=�-�=���=:��=��=���=x�=`x�=YK�=�=2L�=�-�=�$p=BJB=��=���<��<x�v<��-<���;0b�;P��;��;x<�   �   0�_<(ʥ<�D�<���<���<��< ��;����خc�rսB�)�|u�*���OҾ�����a��U#��-�%^1��.���#�G,��6 ��Ӿ�ĥ��Ys�ZJ#�
���*��83-<\9==�!�=P\�=]J�=���=|6�=n�=���=���=gД=�o=x�2=���<�@�<0��; �5�0��H\F�HZW�8#F�0���d�� �9�L�;�   �   h�K< "�<H��<�=L=�Y=T��<��&��B�"~��Ժ�H�B��9��Q&���}Ӿ���c������'��g���	�����]�־�ְ�������G����y�� `���ܜ<&M=_O�=���=��=�`�=���=J��=`�=��=\�8=h-�<0��;(E"��!ϼ>=�$;���K�(gL��:>���#��l ��o��8�%���:�   �   ��<<��<�=�d1=`�@=��8=H~=��<0�ͻx�)��I��B���CL�|���������þ��ھ�)�>����޾@IȾ�����G���Z�Q���Ž��C��ػt�<~^X=���=$�=�4�=ʹ=l��=�u�=�[=ȓ=�)<�\g�2?��y�VE������~�н��Խ�̽`J���F��:�|���4�Hmռ0���   �    �t9���<��=�H=�[e=LMj=�QT=�� =؂�<� ��=��|�������B���v��钾6꥾����Z���﴾͇��誙�����W��?$�+�彑m����漐�;�7=�L\=y!�=m�=���=��=�=��?=@��< -�"��w���eý�+��W��u(�1�0�0���'�*�����#нob��2�E�,����   �   �kC�zn<�:=0W=�z�=+�=-t�=TGl=j@-=8��< ��91����P����4'��L��/k����|���d.����w�lS_��^?���|�ѝ���.�P^C���n<;= /W=�y�=��=Gr�=nBl=0:-=��< ���D1��������9'�r�L�\5k�������W1��1�w�TX_�$c?������՝�b�.��   �   P��`��;�6= M\=)"�=��=��=��=��=��?=T��<������(���]ý�"��R�bp(��1�>�0�:�'�����y�Ͻ^����E�쁻� &w9D�<�=��H=�Ye=Jj=jMT=*� =0u�<�= ��=�h������r�B��v��쒾��𚲾�·�m�銪��������W��B$�۲��p���   �   ��C���ػ��<P^X=��=�=N6�=�δ=���=px�=$�[=��=X0)<H,g�~1��y�L=���<�н��Խ��̽�C��HA��x�|��4�dռ��� �<L��<�=�b1=��@=T�8=�y=p�<�λ`�)��O�����HL���������þ1�ھ/-�� ���i޾?LȾ&���!J��"#Z������Ž�   �   4|���f��ٜ<�M=�O�=`��=(��=kb�=���=���=M�=�=�9=�@�<�L�;�"��ϼJ0�X�:�J�K��[L�(1>�j�#�,f �,f��ȡ%��K�:��K<� �<t��<l=r�=�U=l��<�a(��I����������B��;���(����Ӿ���&��s���)�ni�U�	�������־�ذ�L���r�G����   �   |���R��H,-<�8==�!�=�\�=%K�=Բ�=�7�=�o�=���=D��=�Ӕ=
o=�3=���<�S�<`��;`P5���X;F��=W��F����J�� �9PS�;p�_<8ȥ<�A�<$��< ��<��<���;Lá�\�c��ս�)��u� ,��HRҾN���5c��W#�ү-��_1�r.�4�#��-��7 ��ӾQƥ�-\s�"L#��   �   �f��sG���;��+=�-�=<��=���=��=��=��=z�=VM�=`�=�N�=�0�=Z+p= QB=f�=���<�+�<w<�-<��;0z�; ��;0�;X<p�T<Dۉ<��<���<�x�<�~< 2������e���L�Ð�����9Y�t���)�J�:��aF��kJ��F��!;��M)������ &��:h��l�@��   �   ��<�t��ݙ�,�=���=���=dL�=�
�="�=̋�=@�=�3�=,y�=���=�ǵ=^ݠ=;�=-p=��J=��'=B=l|�<,�<l0�<XTI<x�+< )<0�<<��[<�`t<��l<�]%< �ҹ􈟼&LK��󾽞��l|h��L���Y־���P�!��:��cM�J�Y��'^�G�Y�mM� :��q!����AaӾl2��jBX��   �   ��o��`���=Ş�=�D�=\0�= #�=�>�>�>���=���=س�=��=Ò�=��=U�=�%|=֜V="a2=�(=���<�<@�<��G< h*<�_'<��3<��<<&(<ĩ;�Ȼ�M׼Ɗm�e�Խz�)��Bz������F侬��+��E��BY�Kf�}�j�4Cf�:%Y��D���*�����q��k���g��   �   U�إ��0q3��I=�؍=�b�= �=b��=I�>,�>.>��=�d�=n1�=���=�Y�=��= ��=�&�=��e=�@=b�=���<�ɹ<X܉< nO<(�)<X<��$<P�(<�<��c;H���r꼖Ny���۽�d.�/1���n���龐��'�.�T�H�3Y]���j�I"o���j��-]�QfH��".�������t����l��   �   ��sm�����^=f��=CE�=�0�=^#�=
�>�>�>���=ж�=���=��=�=��=OU�=V&|=��V=b2=�)=���<�<��<��G<�o*<�g'<�3<H�<<X.(<pթ;P�ȻPH׼��m�r�Խ<�)��@z������E����~+�� E��AY��If�b�j�Bf�2$Y��D���*�
���p��j����g��   �   ˈ���t�и����=*��=r��=M�=
�=n"�=��=��=4�=ly�=���=ȵ=�ݠ=��=.p=��J=�'= 
=Ѐ�<<�<46�<�`I<p�+<�)<8�<<p�[<�pt<��l<Hn%< �й�~��FK��ﾽB��lyh��J���W־�����!� :��aM�6�Y��%^�6�Y�#kM�Q�9�2p!�����^Ӿ�0���?X��   �   �`�kG��;��+=r/�=w��=���=^�=���=0�=\z�=�M�=��=6O�=	1�=L,p="RB=̬=|��<�/�<Hw<�-<��;0��;�ݻ;�?�;�$<�U<�<���<��<<��<�<`�L����� �ʽL�y�������[U�7��D)���:��^F�iJ�A�F�#;�	K)��������"���e����@��   �   n���·�HK-<L>==$�=4^�=8L�=���=�8�=Tp�=8��=���=
Ԕ=�o=�3=��<�V�<��;`/5��}�0/F�(/W���E����@ �� ��9 ��;�`<8ե<�N�<���<D��<(�<0Ν;خ��Ҩc��ս�)��u�L(���MҾ����4`�`T#�f�-�e\1�
.���#��*�5 ���Ӿ�¥�8Vs�|G#��   �   �t��xO��8�<�"M=�Q�= ��=X��=Hc�=:��=0��=��=��=�9=�B�<PU�; "��ϼ|.��:���K��XL�*->���#��` ��Z����%��!�:ثK<(/�<���<�=F=l^=���< �%�<� z��>��
�B��7���#���zӾ\���������%��e���	�k���J�־�Ӱ�F����G�z��   �   �C�`sػ$'�<�dX=p��=�	�=�7�=�ϴ=f��=�x�=$�[=d�=4)<`(g�j0�t y��<����нd�Խ�̽�A���>��(�|��4�<Wռ�����<ǻ<`	=Rj1=��@=$�8=ƃ=�*�<P�ͻʯ)��D�����?L����õ��l�þ$�ھ�%�h��L��g޾�EȾx���DE��Z�h����Ž�   �   D�漐T�;Z?=,S\=k$�=3�=��=��=~�=��?=(��<�x�̦����]ý&"���Q��o(�j1���0�o�'�%�������ϽE[��ҎE��t�� ~9|�<^�=$�H=~ae=�Rj=:WT=�� =萙<���~�<�dv������B�"�v��撾�楾��������x봾O�����������
W�;$����"g���   �   �4C��n<�B=�5W=�|�=��=?u�=�Hl=�A-=,��<���081�q������s4'���L�3/k����@���.���w��R_��]?������PΝ���.��DC�ؚn<�A=*6W=f}�=��=�v�=@Ml=*G-=\�<��$-1����������/'�}�L�~)k����3��� +��b�w�M_��Y?�F����ɝ���.��   �    |�9 �<j�=�H=�_e=�Oj=�ST=�� =���<( �=�k|������B�S�v��钾꥾X���&������������F���W��>$�����j������:�;�==�R\=�$�=�=�=�=��=�?=ܥ�<���������Uý/���L��j(�F1���0���'���L����Ͻ�V��ƇE�0k���   �   ؿ<�ǻ<�=�h1=~�@=�8=�=!�<��ͻ��)��I�����CL�f���������þ��ھd)�������޾�HȾ9����G���Z�O����Ž�C���ػ�"�<�cX=���=S
�=�8�=VѴ=x��=�{�=��[=��=H[)<H�f�0#���x��4��M濽ǪнR�Խ��̽,;��$9����|�Ժ4��Lռؼ��   �   P�K<�.�<���<=�=X[=謥< �&�B��}�����"�B�w9��>&���}Ӿy��W������'��g���	������־Vְ�6����G����w��X����<�!M=�Q�=b��="��=|d�=��=Y �=w�=��=~9=U�<���;h�!���μ�!�"�:�
�K�ML��">���#��Y ��O���y%��g�:�   �   �`<ԥ<4L�<���<���<P�<ౝ;x���>�c�.ս$�)�^u�*���OҾ}����a��U#��-�^1��.���#�4,�p6 �ܴӾrĥ�$Ys��I#�������@@-<�<==�#�=j^�=�L�=���=�9�= r�=T��=:��=ה=�&o=�3=���<li�<�S�;`�4��X��F��W��E������� � :���;�   �   �U<��<���<t�<,��<X�<� �Ύ�������L�����,���W�C��v)���:�*`F�ujJ���F�� ;�NL)������$�� g��y�@��c��nG�@�;�+=!/�=~��=���=��=j��=b�=�{�=�O�=�!�=�Q�=�3�=�2p=�XB=��=0��<�<�<�'w<x�-<���;���; �;PK�;8'<�   �   0�<<��[<�lt<��l<�h%< �ѹ����nHK�e�2���zh��K���X־1��k�!��:��bM�7�Y��&^�A�Y�&lM�B�9�q!�=��6`Ӿ�1��AX����t��ə�@�=ѧ�=d��=,M�=d�=�"�=Ҍ�=x�=D5�=�z�=l��=�ɵ=�ߠ=��=z2p=\�J=J�'=�=���<��<l:�<�fI<��+<�)<�   �   (g'<ؗ3<H�<<�+(<@Щ;`�ȻJ׼��m��Խ��)�{Az����F�8�+�E�LBY�zJf���j��Bf��$Y�w�D�M�*�y��Uq�xk��{�g����tn�����n=��=*E�=�0�=t#�=(�>>�>d��=���=ȴ�=��=���=
�=kV�=�(|=��V=d2=�+=���<4�<(�<��G<pp*<�   �   �}>=�1;=�-=��=��<�U��Ă&�����$�(��f���2��]^�L�*��sS�{��"��8��`쥿-����⥿ꜿ�鎿Oz��LR�*�(��� �hr��>'v�ҧ�@)z� �����7=1��=��= ��=p��=@��=��=���=���=�M�=4��=���=�˚=Ӌ�=ܼ|=��f=#U=j�G=b�>=j�9=nG8=r�9=b�<=�   �   ~-<=�;=L�.=<b=��<�`��S������$�[G��_���� �5O'���O��v�����NE���
��h������2��Vk����u�q}N���%����������p������o�@��:E;=���=�g�=���=��=��=���=��=���=��=!��=@�=u��=^ �=��e=��P=��@=xr5=��.=��,=�.=RG2=��7=�   �    �4=0�9=ޞ3=�=���<@�D;r��Գ����	np��"��%$�x���#D��Vi��6��-G��������������1K��)��c�h��kC�j���d�ዪ��b`��n �L�Q�� �;V�D=�=�$�=X��=lM�=�@�=���=~�=�;�=��=�Ֆ=N`�=�[=�U:=� =�*=��=�x�<���<�B=Rs=RD=~�(=�   �   �{%=��5= H9=H)= ��<X�8<p����n���|�a'T�<����Dھ���)Y2�ٸT�SVs�>Ņ������F������K腿7�s���T�|2��S��׾�U���JG�a�ݽ�Z#��N<�nR=��=̾�=V�=���="<�=Z��=^=�=� �=���=��I=�=x��<�T�<8�<p��;0��;@L�;�-!<�u<�0�<�B�<0�=�   �   ��=&�+=d�<=�^9=Ty=|��<�I��zC9�Pͽ�J0�,�9���Y�����(�:��U��k��y��~��z�d7l�b�V��;�C'������3�������'������Ӽ4��<��a=㳠=�p�=@��=ii�=.X�=��=+L�=^�I=t =0�\<`I�D�����㼈� ��z���Y�f���4� �:xfL<Dw�<�   �   ���<�=2�:=��G=+8=�=pe/<hR��}������B�V�4����;�@���&�4���G���S�0X��AT�eH�r�5�B��l�C�ϾK���W����!����,��?�<\�o=�N�=�i�=rF�=(˫=$ܔ=8g=� =x�X<x4����:h�8���䳽�?½'�ý ���Ԣ�S���&aA�7�P��<�   �   ��'<�D�<Vm0=�mP=�mS=��4=d"�< 1��:H"�>��0���Pm�t
���Ͼl ��(���!�dM,�e0���,�P#���������Ӿ�R���;u���%��½B�!�@��;��=�ly=���=���=�Ĝ=ua�=BqH=�_�<��뺌t��opǽfj����#o*��[2�8�0��&��������½o ��\}��R��   �   �5���<r�=boQ=D'i=�._=�0=�ʹ<x���Q�Zbӽ�(�Z�n��8��L��>��k���:��	�ß�\����2�L�ž���.�|���6�4��~�D��h�<,E6=�a|=?6�=���=VGz=�6=�<(�5�
PE��>�����o3�`�Z�Nsz��釾�v��܉���q���%j�D�G�� �(�����<�&��   �   p�� �; ��<�H=w=�s�=�Ek=`R/=`�<��[���^�7~ҽ"e ��?Z��y��������$ž��ʾ#3Ǿe�������}&��{ql��4�ak���l������;D��<��H=4w=fr�=Bk=�L/=L�<0�[�6�^�2�ҽj �fEZ��|��h��$���T(žچʾO7ǾM���k���)���vl�>�4��q��?q���   �   ��~��M���ߕ<D6=<b|=7�=���=Lz=06=P%�<P�5�TBE��6�����bi3���Z�mlz�'懾s��W����n���j�|G�4 �@��@�����&�� �0�<��=BoQ=�%i=�+_=��0=L��<���"Q�biӽT�(���n�<���O��y���������{		��������6���ž�����|�J�6�w9��   �   �½��!� ��;n�=�ly=;��=��=�Ɯ=2d�=|xH=r�< '��f��酽gǽ8e� ��Ui*��U2���0�Ш&��������-�½����u�P�Q�x(<8I�<n0=mP=�kS=��4=��< r���P"��C����hUm�^����Ͼs$��h��!��O,��0�9�,��#�������,�ӾeU��r?u�v�%��   �   ��򡁽�,�8<�<��o=<O�=�j�=H�=]ͫ=ߔ=�g= *=x�X< �3����)h�a/���۳��6½f�ý򝸽�̢������VA�D&� ����<t��<�=@�:=v�G=�(8=��=XR/<p_��ݖ��r����V����� �;^B���g�4�d�G�[�S��2X�TDT�RgH���5��yn���ϾM��n W��   �   �'�:�� �Ӽ���<r�a= ��=dq�=p��=%k�=vZ�=��=�O�=��I=�} =�(]<�QH� u����� 	����d��8D��S���4� C:�xL<�}�<��=ع+=�<=D]9=w=�< n���I9�:TͽPM0���v���\��x���:�3�U��k�c�y�D�~�Bz��9l�O�V��;��(�܆���5��쮃��   �   LG���ݽ�]#�@}N<\nR=��=Q��=6�=4��=�=�=n�=�?�=�#�=���=��I=��=���<�g�< <`޽;���;���;�G!<8/u<H9�<�H�<.�=�|%=
�5=�G9=�F)=��<�x8<T���bq��~~��)T�Æ��uFھ����Z2�t�T�Xs�1ƅ������G������.酿ϓs��T��2��T���׾�V���   �   �c`�Zo ��Q�p�;�D=�=Y%�=��=@N�=B�=\��=(�=�=�=<��=?ؖ=c�=Ȭ[=�[:=� =�0=��=0��<���<�E=�u=F=��(=��4=,�9=L�3=��=L�< �D;x��޵��^���op��#���%�\���$D�*Xi��7���G��a���@���\����K���)��\�h��lC����e����   �   m�p�6���o�@��:&E;=���=�g�=���=���=J�=���=���=���=:��=`��=`A�=۷�=�!�=��e=P�P=8�@=�t5=��.=�,=�.=H2=`�7=�-<=�;=��.=|a=� �<�w��U�β��z$��G����� ��O'�(�O�ȇv�瘌��E��$�����$���2���k��o�u��}N��%��������   �   �&v����r(z� m���7=a��=��=F��=���=V��=0��=���=���=�M�=3��=�=�˚=̋�=ļ|=l�f=�"U=:�G=0�>=B�9=FG8=<�9=>�<=�}>=�1;=l-=L�=,�<pY��`�&����f�(�g���2��w^�i�*��sS�-{��"��A��f쥿.����⥿	ꜿ�鎿�Nz��LR��(��� �;r���   �   �p�����o��ޢ:�F;=~��=Sh�=F��=���=t�=���=���=���=V��=���=�A�=��=�!�=J�e=�P=�@=lu5=��.=�,=(.=FI2=��7=/<=H
;=h�.=6c=��<�R��R�����B$�G����U� ��N'�'�O���v�B����D��j
��
��i��52���j��L�u��|N�E�%�����
����   �   a`�<m ��Q�`<�; �D=1�=&�=v��=�N�=^B�=���=d�=�=�=r��=}ؖ=Rc�=f�[=d\:=� =�1=F�=H��<L��<�G=x=tH="�(=F�4=��9=J�3=F�=���< E;m��S������lp��!��#�����"D��Ui�j6���F������ב�������J��x(��3�h��jC����c����   �   HG���ݽU#���N<�rR=Z�=j��=��=ĵ�=0>�=��=8@�=�#�=Ԫ�=X�I=|�=���<�i�<0<P�;0�;���;�Q!<:u<L?�<8O�<��=��%=��5=�K9=hK)=|��<��8<}l��H{�z%T������Bھ����W2�g�T��Ts�Xą������E������Y煿q�s��T�2�oR�"�׾/T���   �   :�'�#��t�Ӽ`��<��a=���=�r�=a��=�k�=�Z�=�=P�=��I=�~ =�+]<`DH� s��h�㼐�6��8��$?��M��ؤ4� ):h�L<���<��=��+=�<=�b9=b}=ؚ�< $���=9��LͽBH0��@��fW��V��k:�!�U���k�ðy���~�� z�#5l�F�V�;��%�����z1�������   �   ���8�����+�TL�<��o=HQ�=,l�=I�=Ϋ=�ߔ=�g=�*=��X<��3����(h��.���ڳ�6½i�ýǜ��Nˢ�d����RA�L����@�<<��<=��:=��G=�/8=֙= {/<pE��r�������V�	���`�;�>�'����4���G�U�S�w-X�P?T��bH�*�5�2�!k�<�Ͼ�H���W��   �   ~�½��!��;�;�=�ry=\��=���=�ǜ=�d�=�yH=t�<�
��e��酽�fǽ�d�����h*�ZU2��0�:�&�I��1���_�½�����p���Q��(<�S�<�s0=dsP=sS="�4=.�< ����?"��8�����FLm����3�Ͼ�����1�!��J,��0�)�,��#��������w�Ӿ�O���6u���%��   �   d�~��/�����<,L6=h|=/9�=��=&Nz=�6=�'�<x�5�|AE�6�����*i3�íZ�&lz��凾�r�����Gn��j�\{G�V �W��(����&�P���<r�=vuQ=�,i=4_=�0=D۴<��dQ��[ӽ��(�!�n��5��aH����ݩ������	�O�������.�\�ž����Y�|���6�E,��   �   
�� �;|��<��H=~"w=|u�=�Hk=JT/=��<��[���^��}ҽ�d �d?Z�zy�����􍷾�#žg�ʾ�2Ǿ'�������'&���pl�A�4�i���j����� 5;���<J�H=�"w=Vv�=�Kk=Y/=H�<@�[�$�^�~vҽf` ��9Z�Dv����������ž ~ʾ�.Ǿ'��������"��Bkl�Ы4��b��Ge���   �   ��P&�<��=�uQ=�+i=�1_=p�0=�д<��� Q��aӽ��(�,�n��8���K��%��O���+��	����*����2��žɱ��p�|���6�M2��~��;����<HJ6=�g|=�9�=Y��=<Rz=p%6=7�<Pu5��4E�C.��
���c3���Z�gez�n⇾Lo�������j���j��uG��
 ����c���X�&��   �   H)(<�Y�<u0=XsP=�qS=��4=X&�< ���4G"��=�����Pm�`
��l�ϾX �� ���!�XM,�X0���,�<#�ߢ�������Ӿ�R���:u���%�M�½��!�`�;R=�qy=���=���=�ɜ=`g�=*�H=��<@���X��ᅽ�]ǽ�_�:��<c*��O2�W�0�Ϣ&�X�������½��lg�`�Q��   �   ���<�=v�:=�G=Z.8=@�=�k/< P�����d���V�"��� �;�@����4��G���S��/X��AT��dH�`�5�,��l��Ͼ�J���W�W������X�+��F�<��o=\Q�=�l�=`J�=Ы=J�=vg=^3=hY<��3����h�=&���ѳ��,½��ýa����â������GA�,������<�   �   V�=��+=F�<=b9=�{=���<0@���B9��OͽxJ0��+���Y�����#�:��U�ڭk��y��~��z�[7l�U�V��;�2'�c����3��^�����'������Ӽԍ�<@�a=ᵠ=$s�=T��=Fm�=�\�=��=`S�=��I=� =�V]< �G�DY�������������\(�:����4���:��L<��<�   �   *�%=��5=�K9=�J)=���<h�8<��pn���|�D'T�0���zDھ���#Y2�ָT�PVs�<Ņ������F������I腿.�s���T�o2��S���׾�U��+JG���ݽY#�X�N<HqR=*�=���=��=ȶ�=�?�=��=�B�=�&�=3��=�I=�=��<�|�<x7<5�;�S�;P��;�m!<pQu<�H�<HV�<"�=�   �   0�4=R�9=*�3=��=���<�E;�p���������mp�~"��$�t���#D��Vi��6��-G��������������/K��)��]�h��kC�`��td�ǋ���b`�gn �&�Q��+�;�D=��=$&�=҅�=BO�=JC�=���=��=�?�=���=�ږ=f�=<�[=lb:=� =�7=�=|��<$�<�K=�z=�J=��(=�   �   �/<=�
;=^�.=�b=��<�[��S�q����$�WG��\���� �3O'���O��v�����ME���
��g������2��Uk����u�m}N���%����������p�־���o�@��:�E;=L��=Eh�=^��=���=��=\��=���=���=b��=���=�B�=v��=}#�=J�e=̾P=��@=x5=��.=�,=�.=hJ2=p�7=�   �   �A�=o��=F�m=�5=D-�<��y�4����?�y�*���.]�q�7��*l��𐿛�������C�ӿ3߿㿑	߿�bӿC>��\>���B��^ij�r�5����"��(�g�@�����.��5~<J�h=氭=v0�=���=$��=���=��=��=T��=��=f�="|=��a=�JO=6�D=T�A=�E=J\O=�R]=6�m=��}=-s�=�   �   PB�=���=*Om=��7=d۵<�-Z����
��s��຾g���{4�8�g�vb���ȧ�_?��M�Ͽ�Vۿ	E߿�Qۿ'�Ͽ��_���ƍ��Af�@m2� ��Q���b�Uq��%��r�<��j=x"�=�?�=�K�=��=���=6^�=0K�=X˩=�Ĕ=��=8B_=�C=�1=�'=ڳ%=�,=P�8=�J="�]=�yq=:�=�   �   H�w=��{=�k=Tj==%�<p���j�����a�������P_*�pd[���:��&���E�ſsyп�?Կ��п��ſ����)������)Z��(����=��N�R�Tݽ��
���<�o=�=�=6C�=�9�=���=��=���=��=؈=�^=ZE/=��=���<���< �<x3�<؃�<(%�<R=�b-=d�K=b�e=�   �   ��V=�h=�{e=hwD=<_�< I:05��5ݽd�F����z��Ɩ�#�G�X�v��ґ�D���Xi��i��ÿ{��������⥿Rۑ�z]v��3G��y��߾���~w:�Dw����ü0��<,�u=LZ�=��=���=NX�=��=��=�yc=lQ =@#�<Xo<����0�_�X
���G������~*�����;!<�3�<�k	=��4=�   �   @�#=~�J=�Y=�J=�=��8<p��׸����$��+����þ ���/���X�{���̣���Ġ�Cݩ�r��j��:��������OY�</�	"�;����������&��`�:�X�=�{=u��=�Ů=ߕ�=���=��y=�-=�.�<@ﴺ`�����2��Iv�pђ�����������"�u��&8�h�� Z�(�<���<�   �   �h�<�=�D=�K=��*=�T�<  �^l�8���ŻU��Š���߾����[7�^�Z���y��H��%A��D����������z���[�uM8�-��������lOS�D�򽢝J��];��=�l|=f��=���=`�=.U= 9�<p�;��μx�f�<ڱ� 4����z|��r"�ub �������N�׽q[��j�P�ȱ�� ��:�   �   ���F�<pc#=�nD=�==�#
=�K<���q��V1���x�k&�����J� �1�WL�Ga���n�ƴs��mo��ab���M�Є3������瞳�1�|�3	!����xۼx�}<�4=ztw=��=H�v=(;=�&�<�� ���5�m��@��f-���S���r�Lȃ��	��ᅾ�:{�!:`�Je=�J��/�ٽ᱉�T]��   �   ����`O;X�<��3=qI=Z�2=(��< d�\�>��6Խ�y2�:����精�C�l4
����q�0��
<�@�a�<��02���!�pQ�X�����/��]�:�1�ὖ�Q��k��4>�<�D=�j=,�a=�-=��<�C[��a���ս#��]����(����L����Ǿ�I;��ɾFֽ�5����A���Qm��B4��[�������   �   Qp��������V<��=BL=�	S=p�+=��<�=�7d�m���3���}�틥�^W˾7J��2�.�_��������񾋯оM���p���bA� \��{k������p�V<V�=L=�S=*�+=��< �=��Cd��'�� 4��}�̏���[˾>O�5��_b���������񾿳оܦ���r��4gA��b���   �   ����Q�0����9�<��D=	j=��a=��-=���<�[���a���ս��"���]�7���䇥�H����Ǿ�D;̿ɾ�ѽ�"���>���Km� >4�ST����\��� ^O;h	�<��3=(pI=��2=h��<@�d���>��=Խ`~2�)���z벾H��6
����z�0��<�B @�}�<��32�5�!��S�V��W����1��,�:��   �   !!����T�ۼH�}<R�4=tuw=�=��v=�;=�8�< � ���5�m�����_-��S�'�r�eă����2݅��3{��3`��_=�p��I{ٽ����T� g}�O�<�e#=LoD=x�==� 
=x6<(*�����5�i�x��)��t��oL���1�ZL�>Ja���n�"�s�<qo��db���M�L�3����z����@�|��   �   XRS�O���J��.;p�=pm|=q��=Ř�=�b�=@5U=�K�< @�;t�μ��f��б�>)���lv��l"�\ ������i�׽�S��*uP����� ��:pr�<�=P�D=�K=��*=�M�<�. �fl�������U�1Ƞ���߾���.^7��Z���y�-J���B��������������z�	�[��O8�߫�Ǯ�����   �   & ��Ϯ�^)����:�*�=�{=1��=�Ʈ=���=���=.�y=ܼ-=DD�<�Y��`�����2�h8v�tȒ�������ɕ���u��8���༨5���<l�<��#=��J=ƭY=2J=�= �8<�伜���y�$��-���þ���x/�'�X�����)���)Ơ��ީ����������U������QY��/�B#�����   �   ����x:�3y����ü,��<*�u=�Z�=��=J��=XZ�=m�=2�=��c=pZ =�7�<��<pI�� �_��D/�������T*� ���H[!<�@�<�p	= �4=�V=R�h=�{e=�vD=�[�< <H:�5�99ݽ��F������������G�0�v��ӑ�k����j������Xÿ���������㥿;ܑ�_v��4G��z���߾�   �   �=��L�R�`Uݽ$�
��ߦ<�o=�=�=�C�=�:�=T��=|�=���=>�=�ڈ=��^=�L/=p�=���<�ɨ<�/�<�A�<���<�0�<8=�f-=v�K=��e=��w=|�{=�k=�i==�!�<@���j�^����a��������H`*��e[�\����:������+�ſ^zп�@Կ��п_�ſh�����������*Z���(�����   �   R��:�b��q�L�%��r�<��j=�"�=�?�=L�=x�=���=C_�=nL�=�̩=�Ɣ=��=�E_=��C=�1=Z'=H�%=,=�8=�J=��]={q=��=�B�=���=�Nm=Z�7=0ٵ<X4Z������s�zẾޥ�z|4���g��b��eɧ��?����ϿnWۿ�E߿DRۿ��Ͽ���d_�� Ǎ�HBf��m2�4��   �   �"����g�������.�P8~<��h=��=�0�=Ҙ�=<��=���=��=6��=\��=��=f�="|=��a=�JO=�D=*�A=ܓE=\O=�R]=�m=v�}=s�=�A�=G��=�m=��5=8,�<@�y������?�by�`���O]���7��*l��𐿭�������M�ӿ9߿
㿍	߿�bӿ5>��M>���B��8ij�P�5����   �   Q��ńb��o�b�%��v�<"�j=<#�=H@�=PL�=��=���=`_�=�L�=�̩=�Ɣ=��=2F_=6�C=1=�'=·%=�,=��8=�J=��]=�{q=*�=C�=���=DPm=��7=ݵ<�*Z�l����@s�m຾-���{4���g�5b���ȧ�?����Ͽ{Vۿ�D߿RQۿ��Ͽ	���^��~ƍ�8Af��l2����   �   �;����R�aQݽ��
�t�<̨o=�>�=�D�=T;�=���=��=��=x�=.ۈ=�^=�L/=��=���<�ʨ<(1�<�C�< ��<3�<�=h-=�K=f�e=��w=��{=>k=�l==D)�<p���bj�9����a���������^*��c[��]9��h���r�ſ�xп�>Կ��п��ſן��e ��W����(Z��(�����   �   p���u:��s��vü��<��u=#\�=���=���=�Z�=��=y�=N�c= [ =�8�<�< D����_�(-�� ����N*������b!<�D�<�r	=��4=��V=X�h=Re=�zD=�e�<��I:5�C3ݽ��F�㋜���⾺����G���v��ё�6���/h��.~���ÿ7���c���d᥿Gڑ��[v��1G��x��߾�   �   ���+���"���o:���=�	{=ʉ�=Ȯ=���=C��=
�y=��-=�E�<�C������2��7v��ǒ����X�����H�u��8�`��x+�� <`�<�#=4�J=��Y=4J=�=ء8<ĥ�v�����$�l*����þ֎�/��X�X�������Là��۩����������� �����}MY�d/�� ������   �   xKS�;��^�J���;��=�r|=4=���=�c�=h6U=�M�<�F�; �μ��f�:б��(����*v��l"�$\ ������F�׽�R��brP��������:�y�<*�=�D=("K=��*=$_�<x  �rVl�7���r�U��à���߾)���Y7���Z���y�G���?�����e���󻉿�z��[�K8�1����p����   �   6!�����dۼP�}<��4=�zw=��=Z�v=�;=$;�<�� ��5�������_-���S���r�Că����݅�3{�3`��^=�����yٽ)����P� z|�\W�<^j#=�tD=z�==�)
=(f<`
��:���-�
�x��#������G���1�,TL��Ca�8�n�d�s��jo��^b���M��3�l�������|��   �   �ὄ�Q���� N�<�D=(j=2�a=�-=�<�[��a�n�սS�"�P�]����ʇ���G����Ǿ�D;��ɾ�ѽ�粪��=��Km�R=4��R��9�,���@�O;��<$�3= wI=d�2=���<��c�(�>�K0Խ|u2�z���j䲾�?� 2
���t�0�g<��@�)�<��-2���!��N����V���,��u�:��   �   Pd���q��HW<�=�L=�S=��+=�<��=�
6d��㽐�3�n�}�׋��JW˾ J��2� �n_����γ����N�о����o��bA��Z���i��P�����V<t�=ZL=�S= ,=,*�<�m=��*d�����3�k�}�1���S˾FE�F0�Q��\����������оD����l��]A�)S���   �   ����`P;��<�3=�vI=|�2=ܰ�< �c��>�n6Խ�y2�$����精�C�`4
����g�0��
<�@�P�<��02�s�!�WQ� ��؋���.����:�Ǧ�`�Q��M��PG�<��D=�j=��a=��-= �<��Z�,�a�(�ս,�"��]�x�������kC����Ǿ�?;Ѻɾͽ�����:���Dm�84��J���땽�   �    �z�Ta�<Lm#=vD=�==r'
=`U<H�����1�X�x�X&�����J��1� WL�Ga�{�n���s��mo��ab���M���3����׆�����|��!�e���qۼ�}<�4=�zw=��=$�v=d";=hK�<� �t�5��
������Y-��S���r�e������"م��+{�G,`��X=����~qٽ����F��   �   ��<��=��D=�"K=��*=(Z�<h ��\l�������U��Š���߾����[7�V�Z���y��H��!A��?���������
�z���[�bM8�����ǡ���NS�*���J�@�;��=0r|=�=t��=�e�=�<U=_�<���;�μ޽f��Ʊ�^�*��&p�kf"�"V �ޫ�Ӕ���׽�J��XeP������:�   �   L�#=�J=T�Y=NJ=�
=H�8<���^�����$��+����þ���/���X�x���ɣ���Ġ�?ݩ�o��g��6��������OY�,/��!�����������%����:�r�=�{=)��=!ɮ=t��=���=��y=��-=,Z�<��������L�2��&v�������m���������u��	8��p༘��<<�<�   �   ��V=8�h=$�e=�zD=�c�<�eI:.5��5ݽE�F����p����G�T�v��ґ�C���Ui��g��ÿy��������⥿Nۑ�r]v�z3G��y��߾����.w:��v��h}ü���<6�u=D\�=���=$��=�\�=(�=�=��c=�c =�L�<p�<p䔻�p_��ՙ���,߉� #*� s��0�!<�R�<hx	=��4=�   �   ��w=��{=�k=tl==�'�<����lj������a�������M_*�md[���:��$���C�ſryп�?Կ��п��ſ����&������)Z�޲(�n��=���R��Sݽv�
���<�o=�>�=�D�=<�=���=F�= ��=��=�݈=r�^=T/=��=��<ۨ<�@�<�R�<,��<�?�<�=pl-=��K=�e=�   �   �C�=���=�Pm=��7=�ܵ<8,Z�������s��຾e���{4�6�g�ub���ȧ�_?��M�Ͽ�VۿE߿�Qۿ(�Ͽ~��_���ƍ��Af�;m2����Q��b�q�L�%�t�<��j=#�=b@�=�L�=(�=h��=A`�=�M�=6Ω=;Ȕ=~�=�I_=�C=�1=�'=z�%=,=��8=8J=��]=�}q=��=�   �   �L�=5ғ=��=��1=�5;<VJ���ݽ~�S�Lح�����7���t��u��e8����ݿ�T�����Ƨ��
���������ܿaP��)]��3Cr���4��&���O��4E��F���ݓ�'	=(�=g��=���=�=�O�=�&�=p��=p��=��~=6�U=(T3=�C=B�=B�=v�=��!=p�:=�1X=:-w=*��=�ڔ=�   �   =���=��}=��2=��M<�_�e�ֽI�N����	���'4��Mp�o������c�ٿ (��RV���^1�2��H������Mٿ�4��2���Mn�=�1��-��fģ�E<@����������=Ȯ�=�R�=���=
g�=J��=ֹ�=4I�=�L�=�G`=8�3=��=$��<p/�<��<L��<8� =�F=<�>=�a=�r�=/V�=�   �   t�=-�=�@v=�35= E�<���$½�f?�5�����
*�Xrc�4�������Ͽ��(v��$��b	�ڵ�����_꿉�οz&���!��1�a�%�'�V��	z���B2��<��Ȗ:�Ό=W �=���=n�=4�=��=��=��z=p�>=H�=4n�<`3�; �9�� ������ ���0��;4��<@b�<�� =2�N=.�t=�   �   �A[=x�p=��g=�7=`n�<��Ń����'����-�ؾ�P��VO��������,J��w=׿-��ָ��h8�������G뿘׿^���塿%%���(N�`��()վ�k��5�ꥇ��� �=FS�=@s�=z�=ȶ�=��=`wO=�=`E<�����,мH4#���K���^���Z�P�A�nY�`[��0���}?<6�<n/=�   �   �[=��@=D.O=�75=�:�<�{�h�u��	���p�(��Y���5�M�i��`���Ԩ��L���ѿ�rܿQ��O�ܿi�ѿ�ֿ�,@��^�����i��I5��|�ۄ���0j���v�J�P�;&�'=��|=6 �=�M�=��g=�7=XG~<�3�dP������/�����l<��L��D������νظ���`�@�����ߑ<�   �   ��-<LM�<x�)=v^,=H��<��;>1��Dн1g@��^��ѵ߾���$�E�J9t�
c�����������+������w7���Ϥ� ��Gu�|F����b߾�G���<�V�Ľ������i<�>.=�Df=�j=ʖB=���< 
�:���v���g޽N��9��<V�i��p��Jl���\�]DC�F�"�K��������H��߆��   �   x���{<�X�<dT=,�
=T�<����2K���`�$1m���d���o� �:�G�]m��i������N'��T;��֋�� Q��NF��`o�20I�D�!��T���6����m�ȝ��K��(�M���<n�-=�6D=�W&=PY�< :�}?�2
������qL��}���������ӓ���������q���pT���톾�Y�G�"�^6ܽx�z��   �   �;��8���H�6<Da�<.�=���<@�d;���	﻽h�)��������/��n��{�:�\FV�l��*z�L�w�z�ym��X�F�<����5����9������L�-�<��R���;��<<r#=�=�v�<��)��W��Nٽ �-���u�UĠ���ž�澒� �En	�ߪ��*
�0���&�ʾ�@�������M9�>��   �   ћ�6�^��g.���<

=0=�<��ǻ�%F�l�׽�5�ԁ���A��,羶��1�!��3��E>��hB�q?�Mk4�D�#��&����M���I����L=�@��2�^�(Q.����<H
=�=8�<�Ȼ>1F�I�׽5�.����E��1羚��l�!�3�YI>�plB�?��n4�a�#�_)�������I����Q=��   �   ��-�U��ְ�0�;D��<�s#== ��<�a)�VW��Eٽr�-���u������ž��澖� �$k	����z'
�-����z�ʾ�<������wH9�c6�d6�������6<,e�<��=��< ~d;���o�����)���d��K4��8����:��IV��l��.z�$P�n�z��|m�8"X�O�<�D��r���$=��9����   �   ��m�~��O�� N�$��<<�-=�9D=,]&=pi�<��tn?�� ������jL��y�� ��ԣ����������������� P��ꆾ�Y��"�.ܽ�z�X���X�<�_�<~U=
�
=<�<����O��(d��5m�4��h���� �/�G�`m��k�� ���g)��r=��卝�S��H���"o��2I��!�%X��d9���   �   �I��Ɣ<���Ľ������i<�>.=�Ff=Z�j=8�B=��<�}�:����]޽#y�,�9�U5V�D
i�)�p��Bl�D�\��=C�j�"�A��������H�D̆���-<�V�<��)=�^,=��< ��;�7��Iн�j@�&a����߾�����E�:<t��d�����z���"����-������_9��FѤ�����Iu�J~F�L��e߾�   �   ����"3j�>�X�J�0�;�'=X�|=�!�=cP�=\�g=~@=�s~<�X3�^@�t���m%������0��s�����8����ν*����`�Ȭ�t��D�<(a=�@=�/O=�75=�6�<@����u�r�	�#�p�l���Z�~�5���i�(b���֨��N���ѿ�tܿ9��)�ܿ&�ѿWؿ��A��������i�>K5�,~��   �   �*վ�l�����y��� ρ���=�S�=ft�=�{�==��=���=ZO=�=�KE<0����м�$#�ȷK�P�^���Z�T�A��K�(C��д�� �?<�C�<4s/=vE[=��p=��g=7=�j�<&������Ŧ'�=��%�ؾ)R�sXO��������{K���>׿���q���:��L���OI��׿5_��~桿�%���)N�\���   �   J�뾰z���C2��=����:���=� �=b��=��=�5�=��=u�=��z=��>=��=D��<@��; h�����`��� ��� �;hƅ<do�<�� =p�N=Z�t=u�=��=�@v=35=�A�<L��O&½vh?�T��y��*��sc�����宰��Ͽ��Mw������	�h������J�V�ο''��V"���a���'��   �   �-���ģ��<@��������"�=��=[S�=���=�g�=R��=&��=�J�=�N�=�K`=��3=J =ܹ�<89�<���<$��<>� =<J=>�>=��a=�s�=�V�=^��=���=��}=&�2=��M<�a�ΗֽJ�N���������'4��Np�����h����ٿ�(���V�T���1�~��`H�C����MٿK5��p����n���1��   �   |&��lO���E�LF��Xܓ��'	=F(�=���=���=&�=�O�='�=���=���=��~=D�U=&T3=�C=B�=.�=R�=��!=6�:=`1X=-w=
��=hڔ=�L�=ғ=a�=*�1=03;<$K�*�ݽ��S��ح�2��ݠ7�ĺt��u��}8��֑ݿ�T��ʟ���Ƨ��
����	�����ܿJP��]��Cr���4��   �   �,���ã�:;@��������=���=�S�=���=h�=~��=@��=�J�=�N�=�K`=��3=� =T��<�9�<@��<���<�� =�J=��>="�a=�s�=?W�=ƭ�=Y��=�}=��2=��M<_�ֽؕ�N���������&4��Mp�/�������ٿ�'��V����1����G�:���Mٿ�4��ƿ���n���1��   �   չ��x��/A2�/:��0�:���=��=$��=)	�=6�= �=��=L�z=�>=��= ��<P��; ������p��� ���@'�;8ȅ<dq�<� =��N=��t=�u�=��=Cv=�55=|I�<���"½�e?�z����Z*�pqc��ߐ�W���	Ͽ��u������	�D��r���R꿖�ο�%��!����a�*�'��   �   -'վ7j�� }��������x�=_U�=ru�=�|�=���=8��=�O==�ME<`����мF$#� �K���^���Z�V�A��J��@������0�?<�F�<u/=�G[=.�p=�g="7=xu�<(��Y����'������ؾ�O�{UO��������I��#<׿���G����6��%���SF�)~׿�\��_䡿+$���&N����   �   ����6-j���zJ��A�;��'=�|=#�=AQ�=��g=dA=�v~<@V3��?�+��� %��I��u0��:��J�����G�νi���j`��� d����<�c=�@=�3O=~<5=�C�<Hg�2�u��	��p�B ���W���5�B�i��_���Ө�SK��ѿqܿh��i�ܿ��ѿտ��>�����f�i��G5�t{��   �   ,E��Y�<���ĽX���0j<E.=$Kf=*�j=(�B=4�< ��:J�����\޽�x� �9�$5V�
i��p��Bl��\�R=C���"�$@��}���`�H�Dǆ�P�-<T]�<�)=:d,=d��<�J�;*�2@нd@��\���߾�����E��6t�xa��I���������u)����{5���ͤ�q��Du��yF����_߾�   �   �m����E�� �M�X��<��-=
>D=`&=`m�<�pm?� ��ͮ��jL��y�� ����������m�����������O���醾
Y���"��,ܽZ�z�x���h�<,h�<
[=f�
=\��<<���TF���]��,m�6������#� �x�G��Ym�h�����=%��59������O��iD���o�5-I���!��P��y3���   �   ��-������ g�;��<�y#=&=���<HZ)�W�MEٽ@�-���u������žq�澉� �k	����h'
�-�X��F�ʾ�<�������G9�*5��4��P���X�6<�o�<��=���<�Ue;T���軽B�)�I탾��>+�����d�:��BV�L
l��&z��G�g�z�.um�%X���<����j����5�������   �   ��潨�^�H&.�`��<2
=�=��< �ǻ$F���׽�5������A���+羭��'�!��3��E>��hB�c?�;k4�/�#��&�������
���jL=�����^��A.����<�
==P�< }ǻ F���׽�5��~���=��L'����
�!�#�2�B>�eB�� ?��g4���#��#���� �����jG=��   �   �.��������6<�u�<`�=��<�e;���I&�)������/��g��q�:�SFV�
l��*z�	L�i�z�ym��X�1�<��������9��p�����-��	����0A�;���<Pz#==̔�<8)���V�+=ٽ��-���u�����ž�澞� �h	���K$
�*����g�ʾw8�����lB9��,��   �    z����<�p�<]=H�
=��<諊�FJ��j`��0m����Q���f� �4�G�]m��i������J'��Q;��Ћ��Q��HF��Qo�!0I�1�!�qT���6����m�8��#J��@�M�$��<\�-=@D=�d&=�{�< � �`?�����e���cL��u��������������M~����������K���冾MY��"�$ܽ��z��   �   �-<Hh�<j�)=�e,=H��<�5�;
/�Dн�f@��^����߾����E�C9t�c����{�������+������r7���Ϥ����Fu�
|F�|��b߾vG����<�2�Ľ|��� �i<ND.=xLf=��j=��B=@�<���:��������R޽s�C�9��-V�Ei���p��:l�|�\�v6C��"��5��ځ��j�H������   �   �i=�@=�5O=F=5=LB�<pq���u�ګ	���p���Y���5�H�i��`���Ԩ��L���ѿ�rܿO��L�ܿf�ѿ�ֿ�'@��Y�����i��I5��|�����R0j�.��J� )�;��'=��|=G$�=US�=��g=�I=p�~<�"3�j0�?�����a���$��^��������"�ν\����o`�(������<�   �   �K[=�p=|�g=�7= t�<\��/�����'����"�ؾ�P��VO��������(J��t=׿,��ո��f8�������G뿕׿^��塿!%���(N�T��)վ�k���~�������B�=U�=:v�=~�=軞=��=l�O=J= yE<0.����ϼ#��K�H�^���Z�wA�x<�P'���Q����?<�U�<�z/=�   �   Iw�=��=*Dv=F65=�H�<<���#½�f?�*����*�Vrc�3�������Ͽ~�&v��"��`	�ص�����^꿇�οy&���!��*�a��'�E���y���B2�!<��ؐ:��=��=���= 
�=v7�=�	�=�=
�z=��>=��=���<@��; �η�X���Q�� ӎ�o�;P؅<X�<�� =n�N=~�t=�   �   ���=���=��}=��2=0�M<`_�8�ֽ<�N�������'4��Mp�o������c�ٿ�'��RV� ��\1�2��H������Mٿ�4��0���Kn�:�1��-��Zģ�(<@�G��L�����=���=�S�=H��=�h�=T��=e��=:L�=ZP�=�O`=�3=&=��<�C�<��<h��<=�N=<�>=�a=(u�=;X�=�   �   �W�=�7�=$�s=��=0K��/]��H ����W��ч)�V�k��K��O�ÿ��쿚P
��b��#+���4�.`8���4�h+���j�	���h5¿�ə�k�h�e�&��྿K���>�T_��w<(hL=��=���=X��=�6�=X��=y�=��h=8�5=�!=|��<Td�<�Tk<0ws<�|�<xL�<�=`88=��c=���="m�=�   �   +?�=>D�=��o==���5���7Ό����H&�"<g�ݖ��cV��X��"����T)(���1�5���1�(����J������	���1���kd�܄#���۾>���O���U��F<�K=��=��=@M�=�N�="X�=%/�=nH=Ġ=���<�S<`L�;�<;�i; f<j<�U�<=p0I=��u=B�=�   �   k��=��=�c=jz=�BV���j����;h���fӾ�����Z���������oݿ�W��z����(�j�+�0�(�@��|��)���ܿ�ʵ������xX�2���ξ��|����<��M@<�kH=)я=�"�=���=*(�=�m=t,=L��<���;���8I��l�Z`��+ ���μh�v�@T�`~\<`��<N�3=H�d=�   �   �QB=W[=.�M=n�= ΃; (>��_����i�~6��=.�fWG��d��̰��y�˿{ �:W�2��@��ܕ������`���(l˿8�����4�E�C`��S���6a����$��@}y<."A=���=v�=��{=�D=�q�<p��;@���
'�L�}���������ML½����"���匽�K�x�@_���I�<F=�   �   ��<H.=P�*=��= �<��� �ɽ��D��r��'����.��Yi�z���ݴ�5�ӿ4�f|�0�	�H!���	����8��lԿ~-���x����h���-���������Ay>�$��-˼H�<��2=$�Y=��L=�= Zp<(Y\��&;�%7���[�XL���*�3;��`A�Pc=��/�����C�����h�HNм@q;�   �   ����<$M�<$B�<rd<������U��Ru��]P;����E��/}�����1��
 ο>���#����?�����HϿ���Ǧ����}���E���?̾&؃�~����(�O�,C�<t	=T�=$+�<�?,;0����B�� ���)�-.Z��ق�B��x���Y���栾ܠ���;����b�%e3�������Lm)��   �   ƴK���N�Ȋ?<d�<P��<�E����A�a�%,M�)��Nt�Do �AO��g�ʖ��+���;���ſ>fɿ�*ƿ�-���M���䗿������P�UE!��E쾼5��pAL��ས�5�����<��<���<x�<�:��.a(������S�&bX��ӎ������Ͼ&j羶J��6������I�龼�Ҿ|䴾�m����a�#���"ɽ�   �   ��н�jH� 5���5<0L�<�9�;蠾�{���`����p�p=��:A���4"���I��o�#���H�������4������ᖿ�ˉ�,�q�w�K�q�#�����"��^s�$�P��X�����;5�<H�v<@mȻ�0�`vý��%�x�v�,�����׾��������'���2�	�6�']3��U)��h����Cܾu���S,�B�-��   �   ��(��%���� ���y�`�e<h�n< ��X�3ʶ��A$����	���<�X��e�5���P�Bf���s�Z�x���t�ߦg���R��8����2������������(������ ��Dy���e<��n<`V���*Ѷ�dF$�'��5���<A�q����5���P��f�/�s���x�<�t��g���R�\!8�����6������t����   �   $s�d�5T��������;8�<��v<@.Ȼ�0�'ný0�%�m�v�ɒ����׾���S��>�'�ӛ2��6�PY3�&R)��e����>ܾ\��%�\~-���н�`H���4���5<�K�<0�;H���ܲ��L���p�A���E��~7"�m�I���o�T���� ��g�������[��U㖿�͉���q���K��#�A����%���   �   78���DL�	��5��컺���<���<L�<햻�S(�ӈ���M�[X��ώ�̮��#Ͼd�aD���/��_���Y��Q�Ҿ�ߴ��i���a�����ɽ0�K�H�N�X�?<��<0��<pe��6B�+�`0M���6x��q � DO�6k�̖��-��S>����ſ�hɿ-ƿ@0�� P���旿J���b�P��G!��H��   �   ~A̾�ك�����
����O�dC�<=V�=x:�<`�,;~���9��|���)�}&Z��Ղ�b=������`��⠾E����7��H�b��^3�~��a���`)��r���<�S�<�C�<xkd<����ζ��L��zw��WS;z����E��2}�����<��Iο���L&��񿹱�Q��gϿ���g���O�}�"�E�����   �   ����B���L{>��&���1˼��<��2=ԺY=��L=,�=��p<#\�@;�K-��mP��E���*���:��YA�)\=��x/���#���䨷�(�h��5м`;H�<�2=��*=��=(�<����ɽ��D��t���)��Ӡ.��[i�y{��|ߴ��ӿ36ￆ}�^�	�x"���	����'�nԿ�.��z����h��-��   �   (a��T���8a�������{y<V#A=)��=��=j�{=��D=0��<R�;����(
'���}����Ȳ��7B½&���U��5݌��tK�l��`���Z�<� =0VB=Z[=~�M= �=���;,>� c���i�I8��w/��XG��e������˿� X�*��F����
�����.��O*��m˿y9��ᶃ�k�E��   �   ��c�ξ��|�S��J<� M@<rlH=ҏ=R$�=���=�*�=6�m=�{,=ܳ�<PM�;���T1��,S��S�F ���μ�v�@$��\<�<��3=r�d=Ⓛ=��=��c=�y= �V���j� ��5i��RhӾ�����Z���������!pݿyX���4��|�(�.�+��(����w*�r�ܿh˵�!����yX��   �   �#�܊۾8>���O���U�G<��K=���=j�=>N�=P�=�Y�=1�=jrH=��=p�< �S<0|�;@t<;�`i;@|<8~<�^�<ւ=�3I= �u=/�=�?�=�D�=��o=n=@��,6�����Ό��ᾐI&��<g�O����V�����z�����)(�f�1��5��1�f(�@�����J��3
�� 2��@ld��   �   >�&��ྋK���>�p_�xz<�hL=�=✴=���=�6�=l��=��=��h=^�5=�!=���<ld�<�Tk<�vs<�|�< L�<޶=&88=��c=_��=�l�=�W�=�7�=��s=�= Q���]��XH ��������)���k��K��k�ÿ�쿦P
��b��#+���4�.`8���4�`+���\�	�׌�K5¿�ə�<�h��   �   M�#���۾e=���N���U�(O<�K=���=��=sN�=4P�=�Y�=1�=�rH=ޥ=��<��S<�}�;�w<;�di;H}<�<l_�<B�= 4I=|�u=y�=%@�=E�=��o=�=`����4�����͌�]ιH&��;g�����V�������L���((���1��5�@�1��(�������S��d	��W1��3kd��   �   D~�+�ξ��|�,��|
<��\@<oH=�ҏ=�$�=8��=�*�=��m=�{,=���< P�;@���0��XR�TS�� ���μ@�v�@�(�\<��<��3=��d=���=r�=��c=�|= �U���j�®��g��	fӾV����Z�h�������:nݿ^W�|�΢���(���+�p�(������d)���ܿ�ɵ�ݟ���wX��   �   
_��Q��64a���� ����y<�&A=h��=^�=��{=��D=`��<�V�;�����	'�*�}���|����A½ą������܌��sK�<�������]�<f"=XB=f\[=��M=h�=��;~#>��\����i� 5��L-�!VG��c��ɯ��?�˿��hV�F��D��֔�
�����~��S'�Tk˿O7�������E��   �   ��������"v>�l��T˼���<��2=ֽY=|�L=��=��p< \��;�-��)P��E���*���:�XYA��[=��x/�������@�����h�t2м�$;��<|5=b�*=ґ=��<���|�ɽs�D��p���$��h�.��Wi��x��Wܴ�y�ӿ'2�P{��	� �^�	�t��"��jԿ�+��}w��t�h���-��   �   <̾�Ճ� ������O��Q�<�=��=�>�< -;�{��69���{�λ)�T&Z�rՂ�J=��w���D���ᠾ"����7����b�x^3���
���^)��h���<0\�<(O�<�d<�����������ms���M;ǲ�ӪE�-}�'���K����Ϳ���L!�n�񿹬���
Ͽ���������}�v�E�~��   �   �2���<L���߽�5��������<���<��<�ۖ�0R(�F����M��ZX��ώ�����Ͼd�FD���/��>���5��(�Ҿ�ߴ��i����a�l���ɽ��K�h�N�p�?<p��<`��<�	����A����>(M�����p��l �=>O�7d�Ȗ�Y)��9����ſ�cɿ(ƿi+���K���◿˝����P��B!��A��   �   �s��	�YI��z���\�;hF�<�v<pȻ��0�qmý��%�8�v�������׾|��J��2�'�ƛ2��6�?Y3�R)�re���\>ܾ(�m%��}-�p�н�]H�x�4�(�5<\[�< x�;����ŧ�������p�:���<���1"���I�9�o����������������w���ޖ�iɉ�(�q���K�}�#�=�������   �   h�(���� � � �x��e<��n<���f�Bɶ�>A$�w��򐵾�;�M��\�5���P�7f���s�N�x���t�Φg���R��8�����1������W����(�[��ĸ ���x���e<��n< n����1ö��<$�������(7�b����5���P�f�>�s���x�C�t���g���R�J8�j���,��m���,����   �   ��н�RH�x�4���5<P]�< h�;<���;������Z�p�W=��'A���4"��I���o����C����-������ᖿ�ˉ��q�d�K�\�#�����t"���s���aN��H���@G�;,G�<��v<P�ǻ��0�fý��%���v�������׾��������'��2�%�6�aU3�^N)�b���9ܾ�쬾t�~x-��   �   ��K� �N�x�?<@�<ī�<@����A�Y ��+M���:t�<o �	AO��g�
ʖ��+���;���ſ8fɿ�*ƿ�-���M���䗿������P�BE!�fE쾌5���@L�- �ޓ5�@������<P��<x#�<𗖻F(����`H�)TX��ˎ���Ͼ^�>��-)�����(�龔�Ҿ�ڴ�@e����a����3ɽ�   �   X@�(�<e�<S�<��d<Ħ���������4u��JP;z���E��/}�����/�� ο:���#����<�����CϿ���������}���E����>̾�׃���z����O��O�<P=��=L�< �-;�a���0��3q�v�)��Z�<т��8������K���ݠ�s���03��C�b��W3�������Q)��   �   %�<�:=��*=�=`�<~��.�ɽ��D��r��'����.��Yi�z���ݴ�2�ӿ4�d|�.�	�F!���	����4��lԿy-���x����h���-����������x>��"��<&˼��<��2=��Y=h�L=Ȑ=��p<h�[��;��#��(E罤?��*���:�RA��T=��q/�P�2���z���h�h� м��;�   �   �]B=6`[=��M=6�=@�;�%>��^��]�i�n6��:.�aWG��d��˰��u�˿x �:W�0��>��ڕ������`���(l˿{8�����)�E�7`�gS���6a���潦��p�y<,'A=D��=�=��{=��D=X��<��;4v��\�&��}�_��������7½�{��h���ӌ�&dK�������lp�<�)=�   �   X��=��=l�c=�}= �U�>�j�y��*h���fӾ�����Z���������oݿ�W��x����(�j�+�2�(�>��|��)���ܿ�ʵ������xX�*�}�ξ��|�f��v<��V@<�nH=gӏ=�%�=���='-�=T�m=��,=@��< ��;������9켸F�V ���μ�~v� ����\<x�<��3=D�d=�   �   A�=�E�=��o=�=�����4����.Ό����H&�"<g�ۖ��dV��W��"����V)(���1�5���1�(����H������	���1���kd�ل#���۾�=��pO���U��J<z�K=��= �=/O�=:Q�=![�=�2�=�vH=|�=$�<X�S<P��;��<; �i;��<P�<di�<��=�7I=��u=��=�   �   �=��=��T=T�<�ּ�ν�V�y����5�x	R��a���Լ����b���j'�td>���Q��^���c���^�R�Q��>���&�f�a��s��Q�����N�G}�ұ����L�e��h����=�{=�e�=
�=�%�=��=�_=�o%=�V�<@BZ< �D; ����޻��� dƸH]<Lڦ<�	=(�?=��p=�n�=�   �   &>�=$�=��O=p �<@P˼Ƚ\�P�b���xc��'N��֍����������$�h�:���M���Z�N)_���Z��M���:�T$�>����Q���@���BK��
������G�����(N��� =�zu=�.�=+9�=�̒=.�y=j�?=���<��}<@��:@8!�P/��l���`/��p�S���H� J<T�<X�=l�V=�S�=�   �   g=�j=(^@=$,�<
��o� LB�n���4���B�hr��7Q��g>ݿ���FC��,1��B�r[N���R��{N���B�,,1��
�p8��ܿ����&��5n@�����-�� :�Ȯ���,U�x��<��c=�-�=���=�[f=F)=�?�< ';@���4'���J�$qq�H��Px��wW�
�"��꼼�k����w<&g="�B=�   �   �:=�L5=�$=�ٮ< ��������+�A엾e��tI1�i�u�\����n˿_���X���i"� �1��0<���?�,r<��:2�P�"�4��������ʿ��9�s��q/��L�*d����$�򬎽�w���<8oD=�V=V�9=�>�<@��;p�����A�!N���̽������4��J	�3���bս�����\��ټ ��i�<�   �   ��<��<�w�<�<HY%���z�{��_쁾q�о����BX����U���w�ڿϳ���R�$���r&��)�d�&��0�t���H ��iۿ1´��ӎ��MW����L'ξu{~�A
��<c�P=��(`�<r =�)=���<�f�0�Mm���6��&%�}I�;�f��y�t`���i{��j��mN�.)+�q�����N������   �   H��� �̺�U^<�X<`���@(8�d��^�R�����z���6���s��ޚ�\b���bܿa������P���w�BQ�L-��I�ݿRB���W��St�t�6��@��"���JO���ٽ�0&� |ɹ��<�v�<���;�+��Lh��LG�m+�nf�zA��XU��%����̾�Ѿ��;z%������~��;xm�FP2����SW���   �   �i�����x� � ��;�f%�p�u����� ������Ͼ�&iG�<J�K1���s���~Ͽ�}����[�N��/����п9Ը��K��fg��6IH�et��Ͼ����
�LӞ��uڼ ^l:��<�]��L�H��(��O�MS���������0���6�{��V��z������x�Ѽ������U��F��   �   ���FD��8�(��`�A�L1��4�S�J�R�G��B��������o�I�l�x�v䒿SЦ��������\hĿ,N��o���	'���:����z�hK��*��(�%-����H���:�P�H�x��w�����h��A���T8��a�����Xؾ|���)$��<�9lP��!]���a���]�Z�Q���>��A&�.�
�6�۾�٤���f��   �   �b��L	�;s���张1� �߻��ݼ�-��S����^������羳��)=�$a�@���A1���_���]�����������d�c�UP?������ը��b�dI	��n�����P*�����ݼC3��y����^�ꛦ�ß�����=�C(a������3���b���`���㕿���P���|�c��S?�i����꾊ب��   �   �/����H�����P���x��A����0w�D���n3�bza�[���ؾR}�5&$���<��gP�Q]���a���]���Q��>�8>&�&�
�=�۾�դ���f�~��O>����0�� �A��8���S��#��G��E����侤���I���x��撿�Ҧ�Y������GkĿQ��&����)���<����z�:kK�(-�t,��   �   �Ͼ����{֞��zڼ �l:p�<��\�`A�P���	��O�O��h�����v-�u��A2����������K��&s�̼��򒾭�U��A��b��ڵ�x� �P��;�v%��"�ҝ��@� �����5�Ͼo�lG��M�o3��7v����Ͽ������ ^�I����`�п�ָ��M��i���KH�qv��   �   gB�%���MO��ٽ�3&� �ɹж�< ��< =�;|���_���<��+�&ff��<��&P��]����̾�Ѿ��;������az���pm��I2����O��Hq��@�˺Xf^<�X<0«�V-8������R�@���D��y�6���s�����yd��Xeܿ���j��������x��R��/����ݿ;D���Y���t�v�6��   �    ��1)ξ�}~��
��?c��@���c�<�$=D0=ຄ<X4�0�pc���*��T%�`uI��f�X�y�
\���`{��j�wfN��"+�Xk�y��|N�̣��ȣ<��<�}�<���<�a%� �z�����о���4EX�W�����n�ڿ����S����Lt&�r�)���&��1�����I �@kۿ�ô��Ԏ��OW��   �   s/�N�-e��3�$�1����y���<:rD=�V=:=|P�< N�;�h��Z�A��D��1�˽�y�����%��)D	����hXս�����\�p�ؼ�>��x�<�@=ZP5=|$=�ٮ<����m�����+��헾����J1�R�u�����/p˿���R���j"�>�1�2<�0�?�ps<��;2�P�"���0���
�ʿ�󠿭�s��   �   �n@�$��4.��� :������-U�d��<��c=?/�=���=�af=\M)=hQ�<�';x卼���J�Hbq��w����w�jW�8�"��Ӽ�����w<�m=�B=�g=�j=_@=<+�<(��_󶽲MB�Go��Z5�	�B�!s��R��x?ݿV��D�\-1��B�t\N���R�x|N�|�B��,1�"��8�Pܿq��''���   �   'CK�K�
�����D�G�#����M���� =�{u=�/�=T:�=XΒ=��y=��?=���<��}< N�:�!�!�����H!��(�S�@eH�P_<D]�<,�=h�V=�T�=�>�=z$�=��O=4��<PS˼mȽe�P�!����c��(N�e׍�����]��j��v�$���:�$�M�L�Z��)_��Z���M���:��$�x��Q翗���7@���   �   P�N�}�����X�L��������j�=({=+f�=*�=&�=��=N�_=p%=�V�<�BZ<��D;@����޻���� �Ƹ`\<�٦<r	=�?=\�p=�n�=���=��=p�T= �<�ּ#νV������5��	R��a��ռ�ƕ�r���j'��d>��Q��^���c���^�H�Q��>���&�T�B��V��4����   �   4BK���
�������G�T���I��\� =�|u=0�=�:�=�Β=�y=��?=8��<��}<�R�:!�� ������� ��0�S��`H��`<�]�<��=��V=�T�=A?�=�$�=��O=��<DN˼�Ƚ �P����Ec��'N��֍�����_��Ћ���$��:�(�M�6�Z��(_��Z���M�$�:��$����]��󷿘?���   �   m@����T,��D:�%����U�D��<��c=�/�=b��=Rbf=�M)=@R�<��';�䍼��p�J��aq��w���w��iW���"��Ҽ� ����w<zn=(�B=�g=zj=ba@=�1�<h���ﶽKB�Xm���3�(�B��q���P���=ݿ4���B��+1�:�B�xZN���R��zN���B�V+1��	��7�}ܿ����%���   �   zp/�iJ�b����$�m���(`� �<�tD=��V=\:=<R�< S�;�g��܄A�tD����˽Fy���������C	����XսO���\�t�ؼ����{�<dB=�R5=�$=��<���u����+�뗾���SH1��u�f����m˿����z���h"���1��/<���?��p<�f92�8�"�>��#���~�ʿ��Y�s��   �   ���$ξ�w~��
�B4c����n�<(=|2=Ľ�<h0�L0�!c���*��2%�>uI�̀f�2�y��[���`{�Qj�<fN�S"+�k�����zN������<X�<d��<Ժ�<�A%�>�z�Z���ꁾf�оq�� AX����ݹ����ڿ����pQ�Π�bq&�v�)���&�"/�0���G ��gۿ����BҎ��KW��   �   ?�K ���FO�ҋٽ|'&� TŹ���<d��<�P�;H��__��2<形+��ef��<��P��G����̾��Ѿ��;���^��:z��Cpm��I2�����N���l�� �˺hw^<0X<�{��h 8�����R�f�������6�0�s�ݚ�k`���`ܿؿ�����������u��O��*��ߝݿ4@��V��Xt��6��   �   v�ϾA����,͞�|aڼ��n:0�<�g\��>����	��O��N��T�����l-�j��52����|�����7���r��˼���H�U�\A��a������� ��ǃ;`�$�P�G���b� �̃����Ͼ��ofG��F�N/��zq��I|Ͽ�z����X�B��D���п�Ѹ��I���e��3FH�r��   �   �)���|H����P���x��:��`�黖s����3� za�B����ؾF}�+&$���<��gP�E]���a���]���Q�Ӿ>�$>&��
��۾�դ�1�f����<����8�� pA����S���ֱG��?�����;��5�I���x�9Ⓙ�ͦ�ہ��#���leĿ@K������i$��/8����z��dK��'�$��   �   Xb��D	��g��`��`�黰�߻��ݼ,�������^�闦���義�� =��#a�<���;1���_���]������������R�c�BP?�n��Ǐ��Ԩ�b��H	��l�����`���߻��ݼl'��3��a�^�`���������=��a�򌀿�.��O]��[��Oޕ��������
�c��L?�S��ˊ��Ш��   �   ��6���	��n��ZA�$��ތS����G�wB��������f�I�c�x�q䒿OЦ���������UhĿ%N��g���'���:����z��gK��*�_(��,���H���h�P���x�@/��0e��k������.�ta�Q���ؾCz��"$���<�mcP��]�C�a�J�]�~�Q���>�t:&��
���۾NѤ���f��   �   �Y������f ���;��$�L򼧗��<� �􅇾��Ͼ�iG�7J�H1���s���~Ͽ�}����[�I��+����п1Ը��K��_g��$IH�Rt��Ͼ���*
�Eў��iڼ��n:��<@\�5�N����<O��J��i�����(*�ٵ�p.�������,������l徿Ƽ�[p�U�<��   �   0T���rʺ�^<�9X<0~���#8������R�����r���6���s��ޚ�Yb���bܿ`������P���w�>Q�F-��B�ݿKB���W��Et�f�6��@��"��WJO��ٽ0,&� �Ź0ŗ<t��<���;�����W��02�V+�\^f�J8���J�������̾��Ѿ��; ��%���u��Ihm�C2�Z��F���   �   @�<@+�<\��<��<XD%���z���6쁾Z�о����BX����T���w�ڿͳ���R�"���r&��)�d�&��0�p���H ��iۿ+´��ӎ��MW����('ξ{~��
�9c�@���o�<<+=B8=�΄<��D�/��Y��U���%��mI��xf��y��W��X{���i��^N�z+�.e�
���jN������   �   I=^W5=z$=��<p�������4�+�%엾V��oI1�h�u�[����n˿^���V���i"� �1��0<���?�*r<��:2�P�"�2��������ʿ��1�s��q/�|L�d����$�����h�P�<
wD=��V=`	:=�b�<���;dM��uA�N;����˽n�������>	�*��pMս������\���ؼ $�T��<�   �   <g=�j=@c@=`3�<@�����KB�n���4���B�gr��6Q��g>ݿ���FC��,1��B�p[N���R��{N���B�*,1��
�n8��ܿ����&��.n@����r-���:������"U����<��c=1�=A��=vgf=rT)=�b�< _(;�͍���j�J�$Sq�p��8�w�>[W�h~"�亼��ĉ���w<�u=��B=�   �   a@�=�%�=�O=��<�M˼�ȽB�P�Z���uc��'N��֍� ���������$�h�:���M���Z�L)_���Z��M���:�R$�>����P���@���BK��
�������G������K���� =}u=�0�=d;�=�ϒ=6�y=��?=x��<P~< �:X!����<������x�S���G�x<(h�<��=|�V=dV�=�   �   �D�=�t=�.=�y<��C��	�����x`ྌ�,��y��ϩ���ܿ

�
E'��\E���b��|�S���,܉�`�����{��,b�>�D�PG&�0��q�ڿ/���0�u��*���۾�ځ�B��+���k<�TE=���=�c�=ߟ�=;b=�x'=8D�<8�<�,���ʊ�mȼؐ༐�м,$����`��;�]�<�=��M=V�w=�   �   �[w=�7i=�9(=`z<��=��6�W����۾�s)�q�t�>妿'ٿ���Nd$���A�\6^���v�2ۃ�.��r݃�Z�v���]�^A��#�Z���E׿I0��'�q���&�ܟ׾R~�7Z��0�%���h<�?=:�=:��=Z�u=RCD=\�=p!h< �^�H�������#���0��(��G
������什$<8��<D�/=u`=�   �   ܼB=F=Ե=h�<-�l����bt���ξ����g��i��Euο~��$�~}7�&�Q�th�@�w��}�԰w��Lh�̰Q�^;7����s ��Ϳ���e����Q�ʾ�m���J4��9]<~�+=<�[=�X=P�-= ��<��;�B����(��{�TǞ��e��,�������$��ჽ,�7��Ѻ� �����<R=�   �   <��<��=�m�<���;���۽�GZ�VX���%��5S��������á�r��0(�2?���R��_��d��#`�lS�J�?��?(�Fo����߼��-��m\Q��o��<��v�T��mн�c �XV><2L=|�=�I�<@TE<8�\��3�����PtܽBI��r"�p�1�Z;7�L�2���$�����ࡤ�"+F��㕼���;�   �   P����3<�N�<�:Y;���s���I�9�x �\����Z9�\(���a����ӿ����?�^�(�R*9��D�v*H�<�D�*�9���)����� ��ӿ����S��08��q��=j��I5��2����Ҽ���;p�<��|<`�K�j�������콬!&��U���P��(@�� I��(������\u���Y���*��w���⛽
��   �   �xX�г�� �.�`�U�pʼg搽#�xJ��;�Ҿ�)���Y�y��eᵿ2Pܿ�� �<(����k'��*���'�fT���iZ��Wݿm���6��U�Y�ş�2sѾ����n���8����� )�9 @�:����0OG�u�������G\�}����r���о9�����%U��^���p��wӾ5���j����a����}�ʽ�   �   
"彀�x���Ьg��벼Z����n~N����������1���l�����9j���ֿ�O�
&��W���������7���>ؿܦ��m~����m�4�1�z����#����L�����.Q��q����<���ʼ�Xk�Bzݽ�[3� ��|���&������R�.���9���=��i:�� 0����Do
�U^徨n��/�����7��   �   ��>�L��
Uv��H�� ������i���8�MW|��A���>
��:�Ҙo��ⒿQŬ��ÿM�տ�@Ό����E�ֿVſ�=������nq���;���
�����P�|���k��|x�����hn����|K;������ƾ�)�D$�DWD��`��gw�� ��[����l����x���b��aF�-&�:��!lɾ ����   �   j!����2��_ͽ�T�`估�⼾�Q�TT˽�#1�]ދ�
]̾��Q�5�V/a��_��J���7��'���t����#��H7��2��������jc�]�7�s�f9ξk����2��ZͽT�伸��P�Q��Z˽P(1��ዾ�a̾�!���5��3a��a������9��1�������&��&:������ߢ���nc���7��u��=ξ�   �   G�����|�������z��쮼����n�w���E;�2��� �ƾ�&�`@$�SD�b�`��bw����������i����x�#�b�d]F�z)&�R���gɾ�����>�Q��^Lv��@��,���Ԗ��m��2<��\|��E��A
�)�:�Мo��䒿�Ǭ�ܘÿ{�տ	D���a��d�ֿ5ſ%@��� ��Arq���;�?�
��   �   ���%&����L�M��2Q��p��ȳ<���ʼ�Kk�qݽ�U3�
��w��� ⾂������.�c�9�p�=�{e:���/��|��k
��X��i��p���D�7���8�x���⼰�g���<Z����p�N�����������1�,�l�����l����ֿ�R�'��Y�l ����$��3
���Aؿ"���Q�����m���1��   �   ����uѾ ���[���:��(��� ��9��:l����@G�Հ������?\�צ��mm��ٸо��� ���"N��~����꾅Ӿ���*f��N�a�έ���ʽ�kX����� r.�`nU�,ʼN鐽�%��L��>�Ҿ�+���Y�/��v㵿�Rܿ� ��)�����m'���*�j�'�V�z��[��Yݿ�n��R8����Y��   �   D28��s���k���J5�E4�� �Ҽ���;���<0�|< K����K����v��&��T��
�4K��;���C�����ҵ���p��)|Y���*�m���ٛ���� ���@�3<`U�<�CY;����g�����9�tĠ�:����\9��)��c����ӿ7���A���(�
,9��!D�V,H��D���9���)�$��� �$�ӿ����U��   �   �]Q��p�>���T�ioн�d �\><�O=�=@Y�<8}E<(V\��2����^iܽC�"l"�z�1�J47�b�2���$����%w�Ƙ�� F�t˕�@�;���<�=�q�<@��;���@۽�IZ�Z���&�O7S� �����h��n��^(��?��R���_�Ψd�<%`��	S���?��@(�p����༿�.���   �   �e�k���ʾ��m���콸4��=]<��+=ڦ[=�X=��-=���<05�;�*��ފ(��p{����I]��q����������ك��7�<��� ��0ʨ< =��B=�F=��=x�<b-������dt��ξ��E�g�nj��Kvο��%�h~7�>�Q��h���w�6}��w��Mh���Q�<7�v��t �`Ϳ|���   �   {�q���&�"�׾�~�iZ���%� �h<�?=B�=���=��u=tGD=V�=�8h<@^��0��f�#���0�z(�@
��s��@T��-$<$��<��/=�w`=`]w=�8i=:(=�w<|�=�T7�ﬂ���۾Yt)�<�t��妿�'ٿL���d$�F�A��6^���v��ۃ�����݃��v�t�]��A�0�#�����E׿�0���   �   ��u��*�n�۾�ځ����2+���k<jUE=���=�c�=��=F;b=�x'=�D�<(�<�+���ʊ��lȼА༸�м|$�����p��;t]�<ē=r�M=��w=�D�=��t=4.=w<��C�p�	�6����`྽�,�y�Щ���ܿ
�E'��\E�ʨb��|�W���,܉�\�����{�p,b�*�D�<G&���L�ڿ����   �   c�q�+�&���׾~�XX��H�%� �h<?=��=Į�=�u=�GD=��=�9h<�^�`��@�#�f�0�H(��?
�Ds��`R�/$<з�<�/=$x`=^w=�9i=L;(=8<��=�B6�"�����۾�s)��t� 妿�&ٿ���d$�^�A��5^�4�v��ڃ����݃���v�^�]��A���#� ��E׿�/���   �   �e������ʾ�m�	�콌/�XK]<��+=R�[=�X=~�-=���<8�;*����(�^p{�뾞� ]��F���٧�����nك�~�7�$��� ��˨<=>�B=BF=`�=��<�-�����{at�״ξ~���g�i���tο�N$��|7�4�Q�Ph���w��}���w�rKh���Q�|:7�(���r ��Ϳ���   �   �ZQ�jn�;��ҕT��iн\] � o><�R=��=�[�<�E<�S\�v�2�ߙ��"iܽC�l"�Z�1�&47�>�2���$�����v�\���F�hɕ�0%�;��<|�=�x�<���;"���۽�EZ��V���$�P4S�������d����&(��?�
�R�d�_�\�d��!`��S��?�h>(�Pn��m޼��,���   �   �.8��n��h��F5��-��кҼ���;`�< �|<��J�������[v콲&���T��
�"K��;���C����������p���{Y���*��l��Lٛ�J��P�����3<�]�<��Y;̊��������9����� ���Y9�J'��*`���ӿ����>���(��(9�"D��(H�d�D�t�9��)����� ���ӿ��/Q��   �   ���pѾ<�����}3��0p�� ؅9���:(���"?G�8���T���?\�¦��Zm��Ƹо���	���
N��c���Ӟ�eӾ���f�� �a�t����ʽriX�@����*.��U��ʼ␽U ��H����Ҿ(���Y�����ߵ��MܿA� ��&�:���i'�@�*���'��R�f�Y�XUݿk�� 5����Y��   �   H���� ����L���ར#Q�P]��P�<�x�ʼ�Hk�9pݽNU3��	��w��� �w������.�V�9�c�=�me:���/��|��k
�lX��i��C�����7����x�X��؆g�ڲ�z�Y���佄zN�䥧������1���l�����g��?�ֿ�L�h$�V����N�������+<ؿd���P|��N�m�v�1��   �   ����e�|�(������l��ٮ�����	n�5��fE;�����ƾ�&�U@$��RD�X�`��bw����������i��}�x��b�Q]F�h)&�>��YgɾJ����>�Ͽ��Gv��3��������7c���4�R|�g>��5<
��:��o�d����¬�	�ÿ/�տk=�X�忼���ֿTſ�:��X���jq�>�;�\�
��   �   ���J�2�qRͽ�T����Є�2�Q��R˽�"1�5ދ��\̾��H�5�M/a�_��F���7��"���l����#��?7��)���{����jc�I�7�s�79ξ,�� �2��Xͽ&T����ȁ�d�Q�)M˽�1�.ۋ��X̾����5�D+a�)]������34��!���Z���� ��S4��o������8fc���7�p��4ξ�   �   x�>��彤=v�t(������4���f���7��V|��A���>
�ޯ:�˘o��ⒿNŬ��ÿI�տ�@ῲ����=�ֿMſ�=�����~nq�{�;���
�������|�������p�Xٮ����� n�$��D@;�����N�ƾ�#��<$��ND���`��]w�/���𣅿Lg��]�x�M�b�YF��%&�(��gbɾ{����   �   ��>�x��� vg�ٲ���Y�����}N�f���������1���l�����7j��ߨֿ�O�
&��W������|��0���>ؿզ��e~����m�$�1�Q���r#����L�e��~(Q��^��P�<�h�ʼ�=k��gݽ�O3�*��Kr����������.���9��=��`:���/��x�Oh
�cR��d��C�����7��   �   4[X�P�����-���T�Hʼ�㐽S"�<J���Ҿ�)���Y�x��dᵿ0Pܿ�� �<(����k'��*���'�dT���fZ��Wݿm���6��H�Y����sѾ>������C6��xs�� ��9@8�:x���&2G�Sw�����N8\�R��� h��۲о��.���	G��x|��5��J
Ӿe��]a��G�a�>��)�ʽ�   �   �d����3<�f�<@�Y;H���������9�O �E����Z9�Z(���a����ӿ����?�`�(�R*9��D�t*H�:�D�(�9���)����� �{�ӿ����S��08��q��	j��~H5��0���ҼP��;��< �|<�bJ����C푽|k�&�2�T���`F���5���>������ް��il���sY���*� a��Л�����   �   \	�<Ԟ=$�< ��;���,۽(GZ�9X���%��5S��������ġ�r��0(�2?���R��_��d��#`�jS�H�?��?(�Do���߼��-��d\Q��o��<���T��lн�_ �0o><�T=d�=�i�<H�E<#\�X�2�ʐ���^ܽ
=�}e"�t�1�-7�F�2�,�$�Y���k�ێ��$F�|����v�;�   �   <�B=�F=��=��<h-�����vbt���ξ����g��i��Euο~��$�~}7�(�Q�rh�>�w��}�԰w��Lh�̰Q�^;7����s ��Ϳ����e����;�ʾļm�(�콖1��I]<$�+=��[=�X=T�-=���<Ѓ�;l��l}(�~a{�ֶ���T������;���~���у���7���� �t�Tܨ<�=�   �   �`w=j;i=�<(=�<v�=�`6�I����۾�s)�o�t�>妿'ٿ���Nd$���A�\6^���v�2ۃ�.��r݃�Z�v���]�\A��#�Z���E׿I0��$�q���&�ҟ׾0~��Y��܍%���h<P?=�=���=��u=HKD=�=�Nh< �]�D᜼V���#��0�(��7
�pd��`仨F$<���<R 0=�{`=�   �   (#l=�V=@�=ෙ�����=�(�x{��b��� F�	������������R�=��lb�gj���P��"7������0��\3��3%��ʑa���<�>��]���Y���5����C�x ��m��\�#��ぽ�U��X=&�c=�]y=f=�6=�$�<`�6<�Cѻt	��:����.�"P;�j�1���$�ü�T�P�<���<��*=�zY=�   �   Y=POI=�= |��)g��0%��-������ WB��-��,Ἷ�����<�4�:���]�^����
��ݟ��dg��7�������Ts��O]���9� @��:��͉��@�v#��8��: ���}� }�b�=*W=�#f=PL=؇=��< ^8��(����VdQ�Hv�0Ձ�R�x���V�Ѕ �<b���^S���<��	=<�?=�   �   �q=�"=���<p��(,|��#������ �g�7�M���Tu��	�֫���0���Q���q��ֆ��~������s���1��T�q�V=Q��W0����(��G ��`ǂ���5����.��� ��~�k� Rۺh9�<�U/=Z?+=8�<hd><'A�^z�H�~�W����ѽ~�齃:� ��Խ�j���X���V#��wo��!<�'�<�   �   ��b<�<�a�<�⻨za�~�	�� ��8پg'��4q�_����\ֿV�85"�F�>��Z���r�*���K����Ձ�DTs��F[�|4?�>"�
���տ�ɣ��|o���%�qs־�e�{���R��>n���<p��<��<��Z�0��|��-�Ͻ��L�,�dNF��W�1]��X��H���.�F����սP)���U��л�   �   �9�� 	�@=E;��0�H�D�����_�TX����pRT��ӑ�����V���3���(�
@�4�S��`���e�^ta��aT�&�@��t)��~����W���Z���=S����V����[�[� c8���@7�;��:�����Z��XŽ�g�J&K����x��L������:��h�����������N������˽��f��   �   ���P��Ȣ���e��X�,��M���7��S�����@�3�ôx�����?�Ϳ���('��"$��3��:>��B�Z�>�L�4�~%���հ�� >ο���zx�n3�;�����;�4��=��d#��"��88x�ޢ�"��l}���]>�k������Ѿ��������
��G����b�� *ӾJ��2����A��Y ��   �   	J���T�:����� �}a�����[w��gľ����K�n ��G ��ntϿ�V�<��.�jf�Tn �������$�	�,��i�п�ɫ�r�����K�{��c�þ��u�I��������4��B3�Ѳ�����V�Y���� о~t��"��5�O�H��T�YY�l�U���I�x:7������_Ҿ֙���%]��   �   ?�d�&���#���#G�t%���m�J�Խ.N9�R���Yv�Ҥ�8V�h���Ӧ���ÿgݿ3��%���u�����_���޿�ſ=����y���$W�i< �P��̕���8���ӽ��j�hE!���B��}��&�X�b�E���-�羪��c=�u�`��f��O�U�������t�������I����b��>�C1�'꾛���   �   �D��(�W�0d��y���=��*=�s㔽����V��W��(��!�`�P������ɗ�67��J����ƿcpʿ9ǿ-C��/e�������+oR���"����oA��|�W�:a�yv����=�R.=��甽b��f�V��[��-�Z�!�j�P����?̗�<:��EM���ƿ�sʿy<ǿ]F�� h��r���4����rR���"�J���   �   �ᾢΕ�7�8���ӽ4�j�rC!�R�B��w���!���b�������3��C=���`�8d��v�\�������q��짍��F��7�b��>��-��꾤����d�4�����G�d%�T�m�D�ԽJR9�b����zᾯ���V������զ���ÿ�	ݿ��)���w������b�/�޿�ſ����{��(W��> ��   �   x��.�þ��u�j�������\����2�����d��b�Y�����b	оq�����5���H��T�TY��U��I�,67������cZҾ����a]�bE�,����:�����.� �[d������_w�kľ5����K�Z"�����(wϿ�Y�����/�ph�dp �������ҙ	����п�˫�*���m�K��   �   _!3����S���j�4��?���#�����x�������r���V>��������Ѿ��%�������C�7�����$Ӿ>����D�A��T �ܧ���������b��l�,��P��
�7�V�������3�̷x�������Ϳ�����(��$$���3��<>��B���>�F�4�8%����N���,@ο�����}x��   �   C?S���<X����[�e��c8��� a�; �:�����Z�gNŽea��K���oz���F��`|���躾����b���򘾨���L�N�x���˽��f�8$�����@|E;�0���D���Ə_��Z�����TT�4Ց����y��5�d�(��@�J�S�J�`��e��va��cT���@�6v)���n�X��\���   �   ~o���%��t־|g��{�^�R��&n�X�<���<��<�;Z����������Ͻ��dy,��FF��W�)]���W�TH�$�.�N����ս� ��dH���ϻH�b<���<df�<���j}a��	����,پ�'��6q�����f^ֿD�Z6"���>���Z���r�:���_����ց�Vs�>H[��5?�2 "�ʶ�J�տ�ʣ��   �   �ǂ�q�5���쾹�������k��0ۺ@>�<�Y/=�D+=��<H�><�@�m���~�tN����ѽ�w齯0���Խ)b��jQ���I#��Mo�C<�4�<Xv=x"=���<����.|�%�����/�|�7��@v��.鿊����0�ЃQ�T�q��׆��������>������z�q�:>Q�6X0�^������ ���   �   2͉�@��#��I8��Z �Z�}� �|�І=R
W=�&f=!L=v�=��< �6���� �|[Q�v��Ё�,�x�&�V��} �HT��  S��<��	=6�?= 	Y=~PI==����h��	%�n.�������WB�.���Ἷ^���=���:�L ^�ã��W��U����g�����������s���O]�L�9�:@�s��:���   �   �5����C�N ��m���#�}ぽ��T��Y=��c=
^y=lf=d�6=0%�<`�6<�Aѻ,	������.�P;�v�1�2����ü�U�X�<��<F�*=�zY=�"l=JV=��=��������(��{�����F�*������������l�=�mb�sj���P��)7������0��S3��(%����a�h�<�(��4��{Y���   �   �̉�0@�}"��k7��2 �H}}� Y|��=,W=n'f=`!L=��=���< �6����l �P[Q��v�tЁ� �x���V��} ��S����R���<��	=��?=�	Y=jQI=t=�q���f���%��-��f����VB�t-���༿S���`<�ܕ:�0�]�����
��n����f����������r��nN]�x�9��?�r� :���   �   �Ƃ���5�X�����V��F�k���ںC�<*[/=�E+=<�<`�><p�@��l���~�QN��d�ѽ�w齉0�T�¼Խ�a��.Q��ZI#�@Ko�F<l6�<�w=>"=0��<�����(|��"�槐���ﾶ�7���t��3 �L����0�ȁQ�Ϊq�ֆ�~����������m���q�B<Q��V0�*����_���   �   �zo�K�%�fq־�b��x�V�R�@�m��<���<��<�+Z���Q���U�Ͻ��Ky,��FF��W��(]���W�4H���.�"��(�սj ��tG��ϻ8�b<���<�m�<p��4ua��	������پX'�*3q�j����[ֿ��<4"��>���Z�
�r�"���6����ԁ�TRs�E[�3?� "�"����տ�ȣ��   �   S;S���1T���[��NZ8�(��P��; � :8���ЕZ�NŽ:a�tK�Ͼ�`z���F��P|���躾u���b���򘾐����N�<����˽X�f� ��@h� �E;0�0�(�D����4�_�rV�����PT��ґ�6���s�2�p�(�R@�4�S���`�t�e�ra�n_T�V�@�Hs)�N}�w��OU���Y���   �   3��������|�4��7��6#�(�� 
x�Ĕ�9��r��NV>���������Ѿ���������C�)������#Ӿ�������A�T �Ʀ��l��,����S����,��H���7��Q������?�3��x�����-�Ϳt����%� !$��3��8>�^B�*�>�B�4��%��������;ο����wx��   �   #����þ��u�p������L��x��n�2� ������Y�n���J	оq�����5���H�
�T�TY�r�U��I�67������>ZҾt����]��D�����:����` �7\��|��#Ww��dľا�ƯK����&����qϿ�S򿎴�(,�hd�Bl �������^�	��󿩩пkǫ�������K��   �   ��ᾰȕ���8�e�ӽ�j�V9!���B��u��� ���b�������(��8=���`�4d��p�V�������q��䧍��F��&�b��>��-���t����d�q������G���$���m���Խ�I9�m���cr�2���V�V����Ц�ÿ6ݿ��"���s�*���h[򿣂޿�ſ�����w��� W�|9 ��   �   n=��|�W��\�Io��(w=��!=�t������r�V��W���'��!�W�P�����ɗ�27��J����ƿ]pʿ9ǿ%C��&e������栁�oR���"�z��3A����W�0`�Ws��Lz=�( =�3ݔ������V�bT��@#��!���P�k����Ɨ�F4���F��S�ƿ�lʿ�5ǿ�?��b��
󘿀���kR�G�"�e���   �   ��d��������G�<�$���m���Խ^M9����4v�Ƥ�1V�d���Ӧ���ÿdݿ.��%���u������^���޿�ſ6����y���$W�V< ��ᾶ˕���8�>�ӽX�j�9!�ҶB��p����ʚb��{��T�����H�<��`��a���g�������n��	���KD��]�b��>�s*�7�'���   �   �?�[����:������~ �^������Zw��gľ۩�x�K�l ��E ��ltϿ�V�<��.�hf�Pn ������� �	�$��a�п�ɫ�l�����K�j��)�þ4�u�*��|��<��Ԏ뼬�2�����D����Y�6����о�m���S�5��H�#�T�OY�|{U�I�I��17�~�P���TҾ�]��   �   ̞��:�����HM���,��J��@�7��S��{��9�3���x�����<�Ϳ���&'��"$��3��:>��B�X�>�J�4�|%���а��>ο缣��zx�_3���8���V�4� ;��#�T
�� �w�������h���O>����������о��v������?�o�������Ӿ����	����A��N ��   �   <��`��@F;��0���D����G�_�&X����lRT��ӑ�����U���3���(�@�4�S��`���e�\ta��aT�$�@��t)��~����W���Z��x=S�|�\V����[�L��\8����@��;�`":������Z�ODŽ%[�K� ��wu��4A���v���⺾���"]��|혾���^�N����2�˽F�f��   �   8c<�
�<�t�<Щ�va�Ą	�c ��پ`'��4q�_����\ֿV�85"�F�>��Z���r�*���J����Ձ�DTs��F[�z4?�<"�
���տ�ɣ��|o���%�Ns־`e�Mz���R���m��<���<�+�<��Y�������Ͻ���r,�p?F��W�� ]���W���G��.����w�ս{���8� Xϻ�   �   }="=��<����F)|�p#�r���� �d�7�M���Tu���֫���0���Q���q��ֆ��~������q���0��R�q�T=Q��W0����'��E ��_ǂ���5����
��������k���ں�E�<^/=�J+=<%�<0�><P�@��_���~��E��L�ѽn齾&��u�Խ]Y��~I���;#�Po��j<E�<�   �   �Y=�SI=�=Pk��pf���%��-������WB��-��/Ἷ�����<�4�:���]�^����
��۟��eg��7�������Ts��O]���9��?��:��͉��@�m#��8�� �}� �|�h�=VW=�)f=V$L=��=���<�25��������RQ���u��ˁ���x� �V�|u ��D��`�R���<|�	=\�?=�   �   ��S=z<=8m�<p}�VN����A�hU����.�Y�x���{ѿ¤��=*�h�P�Vp{�)�������H��u����B��y���Y���z�P�0M)����Gпߙ��W��r�!��9>���8SR��{�<&�D=<�[=�8G=�s=T4�< ѹ9�薼�A���F�,�i���v� �k�z�I���$5�� 5��Tc�<D�=��?=�   �   �E?=�b.=L&�<��~�*���V�=����y���U��Y��U�Ϳ�g��Q'�hM��Cv�6��0����/�����&3����ỏ���u�PLL��z&����u�̿cA���T���������9�髡�@�T����<@�6=�7G=I+=�X�<�6<��K������S��������菢��l������fhX� G� �c� ��;8k�<��#=�   �   �0 =l#=�R�<d����t�1�Pk��(�UJ�������ÿc���2���B�
�g�����9�������������'T�������yg���A��\������¿������H�.��Tg���b.�B��P`�L!�<<Z=��=�.�< �/:�,ɼj�T�ܭ���ӽXC����	��W��K
�Y����սu���FO[�x�ּ #��tu�<�   �   0��;`�h<8_<����L�����+���9f�a8�lW���������>|1�PNR�0�r�Nh�����ɥ���K��㪇�,s�:}R�th1����3��=��⦃��+7�<Xﾵǐ����=������'<|��<���;h�}��4=�eO��sA����#��F���b�"�t�IO{��zu���c��jH��%�����U���h�D������   �   �~�8 R���뻈-��
��4�	��p}��(Ҿ��!���i�Ϊ���пL%�p��9���S��Aj���y�d��Oz���j�bDT���9�6��
*���ϿfE����h�y� ���о@�z�4}��w�����&��H(6��s	�b������/.�$�h�{����}���'+̾�оʔ̾��������V����j��H0��
��E���   �   S���BN�p�P\���f�l��|R��^�����%F�'����ﲿ�{��������3�NwE��qQ���U���Q��3F�N�4�p2���H�࿚��pe���E��z��K��� P�z.�BC_����T��,�G��3��Y���Z����c	���p龥;�O���e���"�7���p�����꾈m��z䖾��\�_���   �   8&�ԟ̽�-u��Z2�|�X������&��⋾n5۾LP!�=``��<�����x�63��;��#�j#,�(y/���,���#����F���n�
����m�`��4!���ھcE��V%�cD���6T���-��}p�iʽ�$�#�x�?M���p���z/���H��G]��fj�zo���j��^���I�0�M�u��*���P�z��   �   *����&�q�˽�����2^�챖�����[T��k������0�ؼk�6핿v�����տ�3�~�z�
�"$���
�2��g��ֿx������Tl�a 1�_N��s^����S�����Tx����[��4���Rʽ��%� ��a#���:��A(�ܱP��w�f��󎚿]A��JZ��֏�� ������#�x���Q��6)����3#���   �   =-��bju��]�緽�Sy��<y���������t�%���^��R3�,f��I���U���`��S�ͿE�ؿ0�ܿ�Jٿ�vο`K���:�����gPg���3����)��Heu�rZ��㷽8Ry�V@y�:����"�h�t�F���%���3�0f�)L���X���c��յͿ��ؿ��ܿ.Nٿ�yο�N���=������Tg�7�3�B��   �   R��Ra���S������y����[�1��gLʽ��%���������7��=(�a�P��w����ߋ��)>��W���������.���'�x�=�Q�#3)������������&��˽����2^�j�������4`T�Ko�����4�0���k��I���ڶտK7񿞀���
�4&���
��k��ֿ�z��3�����l�,1��   �   )7!�ȹھbG��hX%�YF���5T�V�-��sp���ɽ}�$���x�UH���j�.�5/���H�bB]�eaj�	o�f�j��^���I��0������龏���N�z�$&��̽n%u�NW2���X��º�#�&�R勾9۾�R!��c`�?������{��4��=��#��%,�z{/��,���#�l������q�T���ɉ��U�`��   �   3�E�h|��M��0P��0⽖C_�\�����G��*��|��r�Z�`������1j��7�D��xa�6�"����l�q��'��	h���ߖ���\���y����N�L�hX���f���彬	R�$a����((F�˄����p~࿎��t����3��yE�tQ�f�U�z�Q� 6F�@�4�4�	���e���f���   �   �h��� �y�о~�z�R~��w�(��������6��f	�����d��(.���h��됾���������$̾)�о��̾����8���� ����j�B0�& ��=��@s�8R� ���+������	��s}�;+Ҿ��!��i�U����пx&�rq��9���S�NDj�:�y����Qz�
�j�XFT�2�9�x��+�E�Ͽ�F���   �   �����,7��YﾝȐ����P>��乀�P!'<x��<2�;h�}�%=��E���5��G�#�~�F�p�b���t��F{�jru��c�2cH���%����� ��yD�������;H�h<�i<$���`N��^������Xh�b8�rX��`������� ��}1��OR�(�r�ti���������L�������s��~R��i1����~��>���   �   ~���`�H�����g��rc.�����K`��&�<v^=��=�>�< g2: ɼ��T�����6ӽI9��>�	�,R�gF
�t����սn���xA[�t�ּ ���d��<�5 =�&=�U�<x�f���ʹ1�jl����7VJ�o�����ÿ��������	B�R�g������9���������������T��b��zg���A�N]�Ѫ��V�¿�   �   �A��T����I�����9�۫����T����<��6=�:G=M+=�b�<�N<��K������S�������؊���g�������_X�r?�@�c�P��;�s�<��#=H?=�c.=�&�<��~�.���?�=���������U�1Z����Ϳ�g�,R'� M��Dv��������g0��	����3�����9�����u��LL�{&�����̿�   �   �ޙ�F�W��r�����>����PR� }�<��D=��[=J9G=t=�4�< ��9�疼�A���F��i���v��k���I����5�� <���b�<�=F�?=&�S=�<=l�<� }��N���A��U��G��i�Y�����{ѿ֤��=*���P�tp{�)�������H��t����B��n���K��Ьz��P�M)����п�   �   �@��	T����W�����9�8���H�T�D��<Z�6=T;G=jM+=`c�<�O<��K������S� ������Ɋ���g��貉��_X�@?�X�c����;Ht�<0�#=�H?=�d.=�)�<�~�������=�ؿ��I���U��Y���Ϳfg�pQ'�M�bCv��������^/���~���2�����m���<�u��KL�\z&�^��ߧ̿�   �   8���{�H�T��f��a.�q���;`��+�<`=
�=$@�< �2:Hɼ��T�`���ӽ,9��.�	�R�TF
�H��|�ս:���A[���ּ ꈺ8��<�6 =d(= [�<4냼:���^�1��j����LTJ�$�����ÿ{������B���g�
���-8������������AS�������xg���A��[�������¿�   �   ृ��)7�V�Ɛ���� :�������/'<��<0>�;0�}�b$=�sE���5��,�#�f�F�W�b�z�t��F{�Jru�^�c�cH�z�%��������xD�D�����;`�h<�x<�����I��������d��_8��V��	���ʭ��${1��LR�^�r�9g��l������dJ������8s��{R�4g1��������;���   �   ��h��� ��о��z�bz�jw�Ě�� ױ���5��d	�����(.���h��됾����y����$̾�о��̾����#���� ����j��A0����=��<q�@�Q����8��n����	��m}��&Ҿ��!��i�����пF$��n�B9���S��?j���y����^Lz�L�j�JBT��9�Ϋ��(���Ͽ�C���   �   ��E�y��H����O�4(�h8_���꼜���G��)��(��7�Z�H������j��7�;��oa�-�"�����l�e�����g���ߖ�4�\����b��vN���I��|�e�D��,R�X\��9�v#F������y࿶������3�uE�oQ�>�U�z�Q��1F�>�4��0�0���࿏���c���   �   s2!��ھ�B���Q%��=���*T��-� op��ɽ�$�;�x�9H���j�%�+/���H�YB]�[aj��
o�Z�j��^���I��0�������i����z��&�N�̽z u��O2�2�X������&�����+2۾N!�I]`�;������u⿚1��9�� #�*!,��v/�b�,�f�#��������k㿅���څ���`��   �   �I���Z��z�S������q�� �[��-��$Jʽ��%�N�������7��=(�V�P��w����ڋ��$>��W���������'����x�/�Q�3)�������ƭ���&���˽\|���'^����#���"WT��h���	��>�0�2�k��ꕿ͎����տ>0��|�t�
�"���
�>�d���ֿ8u������V{l�9�0��   �   8%���^u��U��۷��Dy��2y���������t�����P��G3�,f��I���U���`��N�Ϳ@�ؿ+�ܿ�Jٿ�vοYK���:����YPg���3���R)���du�aY�^෽DHy�81y��������t�@���Ȅ��3� (f�G���R��h]���Ϳ��ؿw�ܿ�Fٿ�rοH���7������Kg�M�3�����   �   R���4�&�w�˽�x���%^�����]����ZT��k������0�μk�2핿r�����տ�3�~�x�
� $���
�0��g��ֿx��򍖿El�Q 1�/N��*^����S������s��֦[��*���Dʽ��%�,���;���4�`:(��P���w����׈���:���S��l������H�����x���Q�O/)�������   �   &���̽�u��J2���X�(�����&��⋾>5۾@P!�3``��<�����x�63��;��#�j#,�&y/���,���#����D���n����釔�`�`��4!���ھE���T%��@���+T�T�-��fp�'�ɽ�~$�B�x��C���d辡�/�0�H�M=]�	\j��o���j���]�*�I��0���]�����\�z��   �   �v��b�M�`��\B����e���彙R�`^�����%F�$����ﲿ�{��������3�NwE��qQ���U���Q��3F�L�4�n2���C�࿗��me���E��z�TK����O��+�|:_����D��j�G�"������Z�ș�� ����c�?4�A��:]��"�����h����b��2b��ۖ���\�����   �   Nd�0�Q�p�뻌��X��!�	�p}��(Ҿ��!���i�̪���пL%�p��9���S��Aj���y�b��Oz���j�bDT���9�6��
*���ϿcE����h�l� �r�о��z� |�w���� �����5�LY	�
���p�".���h��搾.�����̾��оB�̾������������7�j��:0�^��g4���   �   �@�;��h<`�<����tJ�����񁒾f�a8�lW���������>|1�PNR�0�r�Nh�����ɥ���K��⪇�*s�8}R�rh1����1��=��ߦ��}+7�X�{ǐ�@��p;������P:'<���<��;��}��=�O<���*����#��F�T�b���t��={��iu�3�c��[H��y%�����謽2iD��f���   �   �< =�,=X`�<郼������1�.k�� �UJ�������ÿc���2���B�
�g�����9�������������&T�������yg���A��\������¿������H�%��2g��`b.����p=`�l.�<@c=�=$N�< �4:d�ȼ��T�]���ӽF/����	��L�A
�:��)zս݅���2[�$�ּ@���䔜<�   �   �K?=g.=�,�<��~�g����=�	���u���U��Y��V�Ϳ�g��Q'�hM��Cv�6��0����/�����%3����໏���u�PLL��z&����t�̿aA���T����	�����9�+����T���<��6=�=G=�P+=�k�<e<0�K�8��F�S�f�����������b������VX�47�8�c� ��;0~�<"�#=�   �   �OC=��*=|�<���?����Q�N��ϵ��=f��i��dܿ��T�3��]�B=�����Q&��Ň��&�����������������']��3��6���ۿ�¢��4e����$���+HO��e���t����<�/=� H=��2=^�<�\U<�Zݻd�׼�{3��l�V+����������r^m�V[5��dܼp��[H<���<,\.=�   �   ��-=�A=��<Ӹ�M���.3M�V�������b�����l�ؿpY�Ly0��uY��f�� V�����R2��1¿��3��J
��r;���7����X�n�/�$��: ؿ��ha�7��>���K�����8�����<&�!=��2=�l=�w�<���:�[���c+�x�z�#�������;Ƿ���8L����|�j�-�lꪼ �}:P�<;=�   �   ���<�L�<ЈN<L���W����@�h����o� V�o���n3ο΍���'��yM���v�YK��$l��έ�����̻��{��-L����v�|1M��6'��5��Ϳ_���8U�ʵ�=���@�>�?~���N����d<-�<���<Po<�E׻^���|��!������S
�\z��t��D�
����Q]���~��;
�`���;_<�   �   �}պhZ<�a;H3ͼ������-��
��Bm ��UC��ċ�;���������� �;��j_�0������u��������؛��;��@����_�P�;����u����4��}[��L�B�l������� ,�-ٟ�L"¼ �a;8�< �,�����lCd�����H>
��a3�3X�Zeu���Nd��t:��#�u��X�f4���
�R½`�g�p
ȼ�   �   H71��䡼�Fc��t�Ԓ����I��#ྫྷ�+�{�v��x��7ۿ	��'&���C�6�`���y�����>�������tEz�2Oa�L@D��B&�<	��ۿU4��jv�N�*��߾�i��ؐ��*����0�R�\v����-�4���)y��z>�� |��������o̾�4ھ߾`ھ��̾Ur��~���>�|�<N?��H��%���   �   �Wν��q��7��x�tx����	c�З����F R�K���Ƽ���쿴���q'�$O>��Q�B�^��9c�`�^���Q�4�>���'�4/�e��7¼�l+�� �Q�K��ۺ��a�Ӱ��;c��>������n���̽:�"��sm��#����;Od���%�4��Am)���,�͌)�&���k�M����Wξ盡� En��#��   �   ��4�-�㽄|��&�T��n}���н��5��V������e+��m�����`ſC��bo�$��6,���5�
p9��'6���,�8��X���I��ſŜ���m��9+��t�ە��4��KϽΔz��yR��h��W��6-4��}���,���h��H��+:�=U�F�j�p5x�<�|�Pex���j��U���:���z���̜���ӆ��   �   q����5����=攽p����I���j���e�ь��'����;�}�y�����v����w�i_����
�������<��
�������1��z̞��z��;�>���V��=be��
�l���퀽aW��+e�,[5�~A����ɾ��	���2���]��1��87���W���`��񇯿X�����������i|�� ^��Y3�5 
�b�ɾ�   �   |�ƾ1���&��7ν���(��Naν�&��3����ƾ�I��S>�9	t�+���4ȯ�{�ƿ!�ؿm�俛�迧��gUٿ�Kǿ:1��!ڕ�}t��>�j���ƾd.����&�4ν����)��fν�&��6���ƾ�L��W>��t�∕�N˯���ƿ��ؿC��~��u��YٿJOǿ14���ܕ�l�t�u�>��l��   �   k���Y��*fe�J�
��m���쀽�S���^�V5��=��Śɾ��	���2��}]��.��84���T��Q]���������͔������y����]��U3�9
���ɾ�m���5��⽂㔽Y���[L���m�F�e�Q�������;���y� ���k����z�0c����
������>��
�p���M⿬4���Ξ��
z��;��   �   ,<+�x�!ݕ�j�4�NϽ&�z�(tR�sc��|�V'4��y���'��!b��f���&:�8U�߇j��/x���|��_x�^�j�1�U�N�:���X���󗼾�φ�*�4���$x����T��o}���нӅ5��Y����龒h+���m������cſ]��0q�4��P8,���5��r9�P*6��,�0��
��gL�l�ſǜ���m��   �   :�Q��L��ݺ�v�a�6���cc��v�����4�n���̽�"��km������;N]��"����h)�(�,�a�)�����g������Qξ$���}=n�0z#��Oν��q�:1��v��y�����uc�u�������R��L��ɼ����F���s'�^Q>���Q��^��<c��^��Q�P�>���'��0����ļ��,���   �   
lv���*��߾�j��	��W+����x�R�Xc��V�-�z��Ds�Fs>���{�����	���i̾.ھf�޾�Yھm�̾�l��������|�>G?�(C�$��+1�Tԡ��4c�Ds�2֒���DK���ྀ�+���v�:z�� 9ۿB	�&)&���C���`���y�0��������Hz�XQa�BD�*D&�L	�Kۿ�5���   �   K\��v�B���������!,��ٟ�¼�@b;`< $*�ԫ���2d�����48
��Z3�"+X��\u�����_���5����u�[�X��
4��
��½�g���Ǽ�nԺpp<��;T3ͼ!��o�-�8��^n �CWC��ŋ�����k �����~�;��l_�F���+��Կ����&ڛ��<��<���r�_�|�;�h��Ց���5���   �   �����8U�O��܄����>��~��pL����d<�5�<d��<8o<�ֻ��t�|�����뽔N
��t�f����
�p���T��Hp��/
� Y�Y_<$	�< S�<��N<l������?�@������p�VV�?���x4οt��t�'��zM�4�v�8L��#m��ܮ�����ͼ���{���L����v�V2M�`7'�6�ǔͿ�   �   I���a�f�?��K�����t���@�<��!=ƕ2=.q=쁰<���:�L��f[+��z����u����������QG���|���-��ܪ� �~:�<v>=��-=�B=��<�Ը�Z���!4M����p���b�����ؿ�Y��y0��vY�[g���V��7���2���¿�U4���
���;���7��,�X���/�X��� ؿ�   �   �¢��4e�W�������GO�e��Ts���<��/=h!H=��2=�^�<8^U< YݻԷ׼�{3�~l�M+�����������^m��[5�8eܼ����YH<,��<�[.=POC=�*=D�<�����?���Q��N�����>f��i��/dܿ*��p�3�8�]�S=�����]&��ˇ��&���������������']��3��6���ۿ�   �   � ���a���>���K�ٺ������<��!=`�2=�q=h��<���:tL��>[+���z����e����������=G��t|�N�-�tܪ��:��<�>=��-=�C=� �<0и�����2M��������b�d��� �ؿ:Y�y0��uY��f���U��1���1������>3���	���:��E7�� �X���/������׿�   �   �����6U���􂬾`�>�T{��D��X�d<,9�<���<�:o<��ֻ$� �|����ҽ뽊N
��t�X�����
�L�콹T���o�f/
�`T�\_<��<�V�<ؙN<諽�y����@�����eo�WV�倘��2οT����'��xM���v��J��;k��ͬ��� ������z��PK�� �v�j0M��5'��4��Ϳ�   �   nZ����B��������,�'՟�D¼`|b;�< �)�ĩ��D2d�D���8
��Z3�+X��\u�����_���5����u�>�X�p
4���
�Y½@�g���Ǽ�7Ժ�z< �;�'ͼ������-��	��hl �zTC�	ċ�(���S�������;�Fi_�1������!���*���sכ�X:��*���(_���;�t��Ŏ��f3���   �   �gv�q�*��߾�g�����%������R�|]����-�sy��s�s>���{�����	���i̾ .ھW�޾�Yھ]�̾�l��n�����|�G?��B�}��)1�lΡ��"c�$e��В�n�H�� �-�+�q�v�Lw��M5ۿ�	�D&&�.�C��`�R�y�J�������
����Bz��La�j>D�LA&�	��ۿ�2���   �   V�Q�"I��غ���a�F����]����������n���̽��"��km������;:]��"����h)� �,�X�)����g�m����Qξ	���:=n��y#��Nνv�q�(,�o��s������c�l���d�� �Q��I��ż����D���o'�M>��~Q���^��6c���^��Q���>��'��-��������)���   �   87+��p�ؕ���4�	EϽH�z��lR� a���z��&4��y��i'��	b��\���&:�
8U�Շj��/x��|��_x�T�j�&�U�C�:���<���җ���φ���4�G�㽛u����T��c}���н�~5�uT��_�龘c+���m�����~^ſ_�m�*���3,��5��m9�n%6�\�,�$�����iF�d�ſ��(�m��   �   ���S���\e���
��d��D瀽 P��(\�NU5��=����ɾ}�	���2��}]��.��34���T��L]����������ɔ������y����]��U3�*
���ɾ�m��J�5�����ߔ������C��
g���e����������;���y�C�������Qt��[��~�
������l:���
���������.���ɞ��z�¬;��   �   �ƾ+����&�,ν���"�� ^νޥ&�63����ƾ�I��S>�/	t�'���0ȯ�x�ƿ�ؿh�俖�迢��bUٿ�Kǿ61��ڕ�}t���>�j�_�ƾ.����&��0ν����!��^Zνk�&��0����ƾG�CP>��t�����;ů�'�ƿ��ؿ��俴����俲Qٿ�Hǿ.��eו�|xt�7�>�g��   �   �i��2�5����-ܔ�����LE��Ci���e���������;�s�y�����s����w�e_����
�������<��
�������1��u̞��z��;�(���V��Tae���
��g��!瀽AM���V��P5�N:���ɾ��	���2�ky]�Q,��J1��wQ���Y��#����~������~��w����]��Q3��
���ɾ�   �   ǭ4�y�kp��n�T�Pc}���нx�5��V������e+��m�|����`ſA��bo�$��6,���5�p9��'6���,�6��T���I��ſŜ���m��9+��t龦ڕ�ƕ4�?HϽn�z��hR��\��Js�~!4�&v���"���[�����8":�-3U���j�-*x���|�Zx���j�$�U�ĉ:�������������ˆ��   �   pEν̻q�D$�fk��s����2c��������> R�K���Ƽ���쿴���q'�$O>��Q�@�^��9c�^�^���Q�4�>���'�4/�b��5¼�i+����Q�K�Nۺ���a�ݭ���^�����X����n�T�̽�"�+dm������;uV��.����Yd)���,��)�����c�k����Kξ���<5n��s#��   �   �1������c�D`�@ђ���JI���ྡ�+�v�v��x��7ۿ	��'&���C�4�`���y�����>�������tEz�0Oa�J@D��B&�:	��ۿQ4��jv�A�*�߾>i�����`'���	��R�LM��@�-�q���m�l>�"�{������gc̾x'ھ��޾�Rھ�̾�f��I}����|��??�=�Z���   �   �Ӻ8�<�;p$ͼ�����-��
��2m ��UC��ċ�;���������� �;��j_�/������s��������؛��;��>����_�P�;����t����4��|[��D�B�L���}���L,��֟�P¼��b;�/<��'�4����"d��v��A2
��S3�N#X�1Tu��� [��l1����u�W�X�`4���
�4
½Ѐg��Ǽ�   �   ��<t_�<��N<�������Z�@�E����o�V�o���o3ο΍���'��yM���v�YK��%l��ϭ�����̻��{��-L����v�z1M��6'��5��Ϳ_���8U�µ����ƿ>��|��E��P�d<�?�<P��<�Xo<��ֻ,����|�o��K��VI
�Ao��
�X����
����K���`��"
� �@}_<�   �   ��-=VF=�#�<Lθ�����2M�F�������b�����l�ؿpY�Ly0��uY��f��!V�����R2��0¿��3��H
��r;���7����X�l�/�$��: ؿ��fa�3��>���K�໸�������<ލ!=��2=�t=P��<�a�:�>��VS+� �z� ���;�������}��1B��v|��-��ͪ� H�:'�<
C=�   �   ��<=��#=h6�<Lc̼�`ǽ1�V�34�����49j�����߿*����6��b�2��Ŧ��y�����������w��ɥ���1��xb�`�6�����߿����)j�r��濾nV���Žnżl�<,�&=�~?=��)=4�<@�*<x�h���IA��cz�Ip��>���b���<z�r4A�d��  ���&<���<�'=�   �   '=2D=��<`Gͼ	�ý,cR��g��d���f�D���2ܿ���\�3��]�cI�����R������QW��`���P����CH����]�>�3�����2ܿ@����e�5�����Q� ����}Ƽ<��<4B=T�)=�=�ߛ<�����ﾼtj9�Ԅ�?s���������X����S��x����`9�D��������)�<�
=�   �   Ȱ�<� �<@-<�TҼ����E�r���&�g�Y������ѿj���r*�lmQ��2|�õ���k��Q��� `������g��w����*|�~gQ��n*�����ѿ�
���Y�S�� ��dE��s���̼��8<�N�<��<x�C<������w7��E���>��>L����!�{v��*�J����������*;������=<�   �   `~��y�; �`84:�٩��2�E�������F�j7�����������n/?��!d��Z���+����q������/���w���d�""?����W��t���3'��h�F�K���9���2��m����ܼ �(:P�;�uh���ۼJ�s�ɵɽ��bV9�ѵ^��H|������ފ�<���
|�Sf^��9��C�fɽ��s��ܼ�   �   ��<����������������������5���.�r�{�:t���	߿&���E)���G�4�e�\����������O������<�e���G�41)�&y���޿Z���W{�2�.��u�q4��|��~R���y��2��TC��l<��7���	�=�D�,����R������]Ѿ�@߾?�h%߾�*Ѿ�p���	��0n���XD�Vt	��
���   �   �ս��~���#���&����3I���h�O̿����~V������9�����|��N�*�x7B���U��Ec�Z�g��:c���U�4B�$�*�J��������ے���U��s�Vs��`Nh�>���$����%���"�a~��;ֽ}�(�i�t�����Ӿ�Y��p��#�� -�qh0���,���"��>�����וҾ8%��t�>)(��   �   ̻9����LC���|a�QW���ؽ�:����A�i�.�uhr�3���ɿ�\� �� �,�/�4}9�J�<��q9�<�/��z �L���"���ȿ���>r�ڳ.�#��i���A:��ؽ���J�`��G������):��T���
���j��L@��F>�p�Y��Yo��}�V倿��|��'o�%�Y�	�=����)���R���G����   �   ����:��뽼����u��Dڲ��"��9l��긾|��[�?�/�~�Q���
�ĿC�忀��2A�����X�����,���3��&RĿ�z���~�I?�̏�3���Ҧk���WU���<��������j4;�|����ξ�� �6��Fb�A셿�7�����隯�u���$����d��#��q���/�a�u�6�����2ξ�   �   �G˾S��e�+��cֽbX��p����ֽ),�J͇���˾����vB�!(y�����YF�� �ʿ�
ݿ��o��M����ܿ��ʿ����[����x��B��9��C˾�|���+�	`ֽ�W��H�����ֽF,�hЇ� �˾���yzB��,y�[���I����ʿ[ݿ��c��,�迗�ܿ�ʿ���u^����x�!"B��<��   �   ��I���Ԫk�D���V���;�����Ԉ�4/;������ξ���6�Bb�酿�4������������Ć���a��,��ͺ����a���6�����-ξv���?�:�4������u���ܲ��%�W>l�2�����?�c�~�᳡��Ŀ���n��LC�2��[�$���.����z���TĿZ}����~�L?��   �   -�.�m�����C:��ؽ������`�B������#:��P�����cd��[<�YB>�W�Y�To��}�q‿,�|��"o�1}Y���=�!������d�������`�9����>���xa��W��O�ؽU�:�/����.��kr�d����!ɿ`���� ���/��9���<�<t9���/��| � ��%�A�ȿ���Zr��   �   ��U�/u��u���Ph�x���$����%���"�$T~��2ֽ8�(�F�t�v�����Ҿ�R��l�l#���,��c0��,�t�"��:�������Ҿc ��ft�q#(���ս>�~�
�#���&���K�!�h��ο����,V�[���<��/����:�*��9B��U��Hc�F�g��=c�>�U�^ B��*�������ݒ��   �   �Y{���.��w侨5������R���w��&���/��<^<�j.���	���D�����SM������gWѾ8:߾t���߾�$Ѿk������i���QD��n	�E��$�<� r��������z��� �����������.��{��u���߿d��RG)���G���e� �����RË�ʜ��D��v�e���G��2)�>z���޿_[���   �   (����F����:���2�cn����ܼ��): O�;��g��ۼ��s�s�ɽ���0O9���^�@|�񚇾�ي�����||�u^^���8��=�G\ɽ
�s�(�ܼ��}����; 0l8:⼘ک���2����������F�~8��F���� ��&���0?��#d������������As�����j���~����d�Z#?�����������   �   ����Y���)!��E��s��p̼��8<�W�<���<��C< Z�����/��[���4���F�<���!��p�^%��������Z���.� ��h�=<h��<�'�<@-<�UҼl��P�E�Cs��|'���Y�z����ѿ���s*��nQ�4|������l��e���a������h��@���(,|�bhQ�6o*����j�ѿ�   �   I@����e�d��F���Q�����{Ƽh��<�D=��)=2=�<@�ྼ�a9�Vτ�n��W�������
����N��계��X9�|{������|2�<T
=r'=�E=��<�Hͼ�ý$dR�Wh�����f��D��_3ܿ���܀3���]��I��r���R��F����W��跿��P��q���H����]���3�ޘ�3ܿ�   �   ���L)j��q��濾V���ŽXlż��<��&=^?=�)=��<��*<H�Д�IA��cz�5p��8���b���<z��4A����� ��&<��<��'=0�<=N�#=@5�<�d̼jaǽ��V�|4����r9j�����߿B����6��b�2��զ��y������������w�������1��Zb�F�6������߿�   �   �?����e����A��ĤQ�P���HwƼX��<�E=6�)=�=��<�舺�ྼ�a9�Bτ�n��H������������N��ೄ��X9�{��  3�<�
='=vF=x�<|DͼV�ý�bR�Pg��0���f��C��r2ܿd���3���]�I������Q��(����V��˶��|O��� ���G���]���3�D��"2ܿ�   �   �	����Y�j�4��|E��p���̼�9<p[�<��<8�C<�W�p���/��2����3���F�.���!��p�R%�x�������0���.������=<Ƚ�<<+�<X)-<MҼ����E�Oq��&���Y����ѿ��"r*��lQ�t1|������j��K����^�������f�������)|�dfQ��m*�x����ѿ�   �   &����F���48��s2��i��Լܼ��*:�b�;��g���ۼ��s�!�ɽ���O9���^��?|�嚇��ي�����i|�^^^���8��=� \ɽX�s� �ܼ@r}���; �{8H.�֩�R�2���������F��6������g��&��8.?�P d�腄����̏��dp��=���ᒔ�X~��(d�� ?����
������   �   1U{�N�.��r�w2��|���M��bp����*��B\<��-��ش	���D�����AM������XWѾ*:߾h�㾶߾�$Ѿk������i���QD�~n	����<�<�(l��H���Ȕ����ǟ�T����侁�.�`�{��r���߿��bD)���G���e��������9���˙��ڋ���e���G��/)��w���޿gX���   �   ��U��q�hp��Jh�������%���"��P~��1ֽۂ(��t�Z�����Ҿ�R��l�d#���,��c0��,�l�"��:������ҾK ��(t�#(���ս~~�
�#���&�"��xF�;�h��ɿ���0V����8��'������*�N5B���U� Cc�p�g�
8c��U��B�6�*������g���ْ��   �   #�.���y����<:��
ؽ������`��?�����n#:��P��d��Fd��M<�MB>�N�Y�To��}�m‿$�|�y"o�(}Y���=�������F���[���޵9����R<��qa��Q�� �ؽh�:������.�Per�3����ɿZ�B��� ��/��z9���<�<o9��/��x �t��o�'�ȿ⃟��r��   �   <��c���5�k����7N��86��(	��k��t.;����W�ξ���6��Ab�z酿�4������z������������a��(��Ⱥ����a���6�����-ξ:�����:���;��o��#Բ�4��4l�G績1��Q�?�N�~��3�Ŀ��忤��&?�����V�����*�������#OĿjx���{~��E?��   �    ?˾$y��ę+��WֽxP��<z��}�ֽ
,��̇���˾����vB�(y�����TF���ʿ�
ݿ��l��J����ܿ��ʿ����[��|�x��B��9��C˾?|��ڝ+��\ֽRR��Ty����ֽ�,�8ʇ���˾�~�sB��#y�����SC����ʿ�ݿ<��y��c��,�ܿ)�ʿ���Y��Խx��B��6��   �   ����R�:�뽆훽�n���ղ�v!��8l�\긾h��M�?�$�~�M����Ŀ>��~��0A�����X�����,���/��#RĿ�z���~��H?���������k�����P��6��_������);�,����ξ��B�6�l=b��慿�1���}���������W���Y^����	�����a���6�����(ξ�   �   �9�4��7���ka��Q��K�ؽ��:�:���Y�.�khr�.���ɿ�\��� � �*�/�2}9�F�<��q9�:�/��z �J���"���ȿ���7r�̳.�������?:��ؽJ���8�`��;������:��L��t ��^���8��=>�X�Y��No�}��߀�l�|��o�xY�
�=�&��K������T����   �   m�ս4q~��#�(�&�T���G���h�̿����vV������9�����z��N�*�x7B�~�U��Ec�Z�g��:c���U�4B�$�*�J��������ے���U�~s�s��qMh�º� ��܃%�P�"��E~�')ֽ}(�d�t��{����Ҿ�K��h�#�"�r�,�=_0���,��"��6�����ŉҾ:���s��(��   �   ��<�Y���}��Z��y��� ����������.�l�{�8t���	߿$���E)���G�2�e�Z����������O������<�e���G�41)�&y���޿Z���W{�'�.��u�4��_���N��~o��������O<�+%��5�	�v�D�D���1H��̧��QѾ�3߾���߾>Ѿ+e��N���Pe��)JD��h	�g����   �   ��|����; �8 +�}֩�U�2�
�������F�j7�����������l/?��!d��Y���,����q������/���x���d�$"?����X��t���3'��b�F�<���9��.2�Xk��мܼ�q+:���;@5g��oۼ �s�Y�ɽ�{� H9�ĥ^�Y7|�Z���KՊ������{�SV^���8��7��Qɽ��s��ܼ�   �   P��< 4�<4-<�JҼc��d�E��q���&�d�Y������ѿj���r*�jmQ��2|�ĵ���k��Q��� `������g��x����*|��gQ��n*� ����ѿ�
���Y�K�` ���E��q���̼�9<0b�<���<��C<�0�H��-(������F*��~A��~�
!�4k����������}���!��~��><�   �   >'=�H=��<�BͼA�ý�bR��g��`���f�D���2ܿ���\�3��]�cI�����R������RW��`���P��
��CH����]�>�3�����2ܿ@����e�2������Q�V����xƼ��<�F=��)==��<@1���Ҿ��Y9��ʄ�i�����.��������I�����P9�@l���%���=�<�
=�   �   �=A=��(=p�<x��� ��)�P�8���=,��ke��Ԣ��ۿL9��3��*]����xÝ���#����,�����*��`��?��ڷ]�ʜ3���=pܿ�t��
Pf�����^����Q��O��\C��4m�<��)=�GB=v�,=p��<�><������r�8���p�a3���.���ɉ��To�F�6��m߼�	 � �A<4#�<�X,=�   �   ��+=.Y=��<8|���P����L������O�Wa�B��%ؿ8����/�tY�i;���@�����:��zȿ��6��~���W��h���xY�}0�^�h�ؿ!���,b��������qEM����0H���H�<Ԅ=�,=��=T��< ��9$��t1�� �����!Ų�re���K��E2����}��/����� �:$��<�R=�   �   �f�<$��<�8H<���������b@��?����oyU����Ϳ
>�?'�0;M���v�aS��͂���®���������l��5J����v�,wM���'����i7ο�����$V��x��ǭ���@�L3��@����K<x�<���<��V<���l�х���<����8��������4���4�ﭹ����V1� �����X<�   �   ��p�<@n�:̛ϼ�3���-�Ϻ��<$ ��B��|���R��^�������;�B�_�ݱ���D���ߛ�{���Ҿ��-������D`_���;��������5���Tċ��XC��r ����T.�V��	ϼ�7�:8u<����ͼzk��Ľ���'5�g�Y���v�����Ç�jj����u���X�8�3�c�
�}½D$h�|ʼ�   �   212��Ȥ�h�i��[���M�����)��v�߾�K+���v�]��O/ۿ`-	��Z&�YD�Pga�&Zz�������������y�d�`���C��&��	�+$ۿ�l����v��~+�C ྵZ���K�cd���q���k��ᦼ�T4���� a�΅@�N"~�,������G;v�ھ�[߾Xsھݚ̾F/���:��.Q|���>��!��F���   �   �ν�s����.0�;��"����*c�l������R�?]����������L���'�.�>�h�Q���^�
>c�(~^�VrQ� ;>��['����,z쿻����9��C�Q���|����;c�_����R���������3u��^н�$��o�>Y��cϾ����w��� �O�)��-�ց)�����!�dU���;�.��3�m�Q#��   �   ƨ4���㽥O���V�B��a�ѽ&�5��:�_�+��n�\��}�ſ��ￆ��b���,��66��s9���5�0&,��n��W���O:ſ�����m�eQ+���龳h��0�5���ѽ�����W�F��q����5�`����j�������x��;��V�r4k��x��}��=x�րj��"U�:�����A���#��/����   �   �X��}�5���㽑����V¬��4�8�f�����0��$<�܅z�e���w��mF�6��(��K�(�����
��6��vJ����e����y�4{;����Y���()f����͏��~6���Ɩ�����6�+���ʾ�
���3�a�^�i���q����ģ�r���Ǖ���^���H������� M]���2��	�v�ɾ�   �   ��ƾR��� '���Ͻ�ԑ����sнz�'��䄾G�Ǿ$��D?�u�����s��Y�ǿ_�ٿ��俣�迹����ؿӺƿ*���ga��>�s�G'>�^1��ƾfO��='��Ͻ�ӑ����9xн��'��焾��Ǿ��?��u��!���v��ʊǿ�ٿ��俅�迅��t�ؿ"�ƿ ����c����s��*>�	4��   �   ���d���-f����b���~5��FÖ�
���6�v'���ʾ��
���3��{^�����p���K������b���V[��~E��,�����H]���2��	��ɾsU����5�(���������Ĭ�|7���f�;��D3�(<���z�����z���I��9��8��M�Z�����
�}:���M�͠���g��^�y�&~;��   �   �S+����j����5� �ѽV��8�W��@��=���5�c����e��Z���u�A�:��V�/k�:�x�+}�Q8x��{j��U��:�J���;�����~���l�4�p��:K��T�V�j����ѽL6�{����=���+�n�����ſ���V��t��,�.96�vv9�
�5�j(,��p�\Y�ԫ<ſ����m��   �   ��Q��������q>c�Ƶ���R��¥����&'u��UнĪ$���o�;T��YϾx������� ���)�\-�l})�c�����N��H�;?*����m�_K#��νh�r�b��.�(<������.c��������	R��^�����T �zN���'�h�>��R���^��@c�ހ^��tQ�=>�t]'�d���|쿡���';���   �   ��v�6�+�8"��[��M��d��m����j��Φ��F4�����6[�t~@�p~��&�����@A;��ھOU߾�lھ��̾�)���5���H|���>�n�9>���$2�������i�Z��O��� ��+����߾�M+��v��^��H1ۿ�.	�\&��ZD��ia��\z��������p���f�y���`�N�C��&�	��%ۿ+n���   �   %ŋ�'ZC��s ����W.��V���ϼ@��: �<�v�ܪͼ�k��
Ľ��� 5�s�Y�2�v���������e��E�u�ԮX�d�3���
��½�h��ʼ�����<@��:��ϼ25����-�A���V% ���B��}��%T��������H�;� �_����E��:��ߖ��'���^�������a_�Ζ;�r��H���I����   �   -���`%V�{y�9ȭ���@��3�������K<L�<���<h�V<�v�:_�2~���3��4����,��o��,/���G+�������P%�Д��P�X<q�<ԯ�<�>H<|������1d@��@�����zU����#�Ϳ�>��?'�B<M���v�=T��ʃ���î��������om���J����v�
xM�L�'���$8ο�   �   Z���b,b���*����EM�m���tF��L�<2�=b�,=��=���< ϡ9T���1�������ӿ��`��iF��b-����}��/�����:��<V=��+=�Z=��<�}���Q����L�>���6P��Wa�����ؿ���\ 0�Y��;��_A������;��	ɿ�s7����� X��ih��yY�L}0�<^���ؿ�   �   �t���Of�����^��.�Q�hO���A��hn�<�)=HB=��,= ��<�><x��T��8�8�X�p�N3���.���ɉ��To�p�6�n߼�
 ��A<�"�<8X,=�=A=�(=P�<���� ����P�����n,� le�բ�8�ۿb9��3��*]�����Ý���*����,�����*��Q��n?����]���3���pܿ�   �   ����V+b�R��(���DDM�����B���N�<�=��,="�=`��< �9����1�������ſ��	`��ZF��Q-����}��/����� :���<�V=��+=|[=��<dy���O��>�L�>���yO��Va����ؿ����/�Y� ;��}@�����m:���ǿ�Z6�����;W���g��xY��|0��]���ؿ�   �   Ӆ��_#V�x�Mƭ��@�R0��������K<��<d��<��V<�t��^��}���3����ט���`��/���++�g�������$�p���P Y<`s�<D��<`IH<,��������a@��>��P��xU�}��g�Ϳ�=�t>'�V:M�j�v��R��恢��������z����k��VI���v�vM�֌'���b6ο�   �   DË�_WC��q � ���.�R��8�μ@5�:8�<�[���ͼk�M
Ľz�� 5�X�Y��v�u�������e��3�u���X�L�3�r�
��½:h��ʼ�q�p�<�A�: �ϼ�0��;�-�����b# ���B��{���Q���������;���_�ఁ�kC���ޛ����t������l����^_�B�;�x��/���ڠ���   �   $�v��|+����X���H�s_���^��8�j��Ȧ�E4������Z�<~@�A~��&�����1A;��ھAU߾�lھ��̾�)���5���H|���>�;��=��#2�ز����i�PL���I����f(��U�߾4J+���v��[���-ۿP,	�4Y&�^WD�*ea��Wz�3��������~��*�y��`���C�&��	�-"ۿ<k���   �   ��Q��������7c�Ѭ���L��������#u��Tнf�$���o�T��>Ͼc���{��� ���)�U-�e})�\�����N��6�;**����m�K#��~νN�r�~���&�V6������O'c�	������R��[�����e��zK�<�'��>���Q�6�^�6;c�f{^��oQ��8>��Y'�b���w쿙����7���   �   �N+�����e����5���ѽn��l�W�Y>�����t�5�2���|e��<���u�4�:�|V��.k�3�x�#}�J8x��{j��U��:�B���;�����V����4�����H����V������ѽ��5�t����6��+�{n�e����ſ������h�f�,�L46�xq9�,�5��#,�~l��U�٥7ſ폜���m��   �   �������#f����ʈ���/���������6�4'���ʾ��
���3��{^�����k���F������^���S[��{E��)�����H]���2��	�ɋɾ:U��<�5����*��V���S���1�b�f�o���.��!<��z���(u��/C�o2��$�
�xI������Ԕ
�3��G�����b��l�y��w;��   �   ��ƾ
L��/'�!�Ͻ�̑����0pнi�'��䄾�Ǿ��7?� u�����s��U�ǿZ�ٿ��俠�迷����ؿҺƿ(���ea��7�s�>'>�Q1���ƾO��3'�̲Ͻ�Α�����lн��'��ᄾ+�Ǿh���?���t�?���p���ǿ��ٿ��俽��߅�*�ؿg�ƿ����^����s��#>�h.��   �   �Q��$�5�7�㽃��N���㽬�@3�N�f�v���0��$<�΅z�_���w��jF�6��&��K�&�����
��6��uJ����|e����y�*{;�������L(f�P��a����/��ּ��彏�6��#��\�ʾ��
��3�w^����~���������������W��DB��,��e���C]���2���	�݆ɾ�   �   �4���㽑C��N�V�����ѽ��5������9�O�+��n�W��x�ſ��ￆ��b���,��66��s9���5�0&,��n��W���M:ſ�����m�ZQ+����\h���5�0�ѽ�����W��9��X���5������`�����Uq���:���U��)k���x�p}��2x�!vj��U�B:�e��5�����`����   �   �uν��r�����"��6��)����)c�%������R�;]����������L���'�.�>�f�Q���^�>c�(~^�VrQ� ;>��['����+z쿽����9��<�Q� ��<����:c�q���N�����P���u�gLн��$�$�o�^O��vϾ�������x �e�)���,��x)������G��7�;1%����m��D#��   �   �2� ����}i�`G��&J�����)��C�߾�K+���v��\��N/ۿ`-	��Z&�YD�Pga�&Zz�������������y�d�`���C��&��	�+$ۿ�l����v��~+� �bZ���J��`��(]��h�j�d����84�s���iU�>w@��~��!��0��;;J�ھ�N߾4fھc�̾�#��q0���?|�H�>�]��4���   �   �� ���< ��:�ϼ-1��:�-�����+$ ��B��|���R��]�������;�B�_�ܱ���D���ߛ�{���Ѿ��-������D`_���;��������5���Tċ��XC��r �v���.��S��4�μ ��:H�<@���ͼ��j�� Ľ����5���Y���v�����w���fa����u�ܦX�E�3�g�
��½�h�d�ɼ�   �   ��<��<�SH< ������Rb@�f?����jyU����Ϳ
>�?'�0;M���v�bS��͂���®���������l��4J����v�,wM���'����j7ο�����$V��x�tǭ�{�@��1��������K<�!�<���<8�V<N��R��v��$+�������~�����)���
�m!���� ��R��=��� Y<�   �   ��+=�]=�	�<�w���O��d�L�p����O�Wa�B��%ؿ8����/�tY�i;���@�����:��yȿ��6��}���W��h���xY�}0�
^�h�ؿ"���,b����朸�6EM�����tC���O�<~�=L�,=��=H��< ��9H���1�������������Z��&A��M(��<�}�:�.�8��� �:̶�<�Z=�   �   �OP=v�8=H�<�L���ꪽ�@��A�����`X����l+п����W)��P�8�z����������Q��a����U��̥��0��"|{��Q��G*�į��ѿ�!����Y��������B�Dꬽ�(���q�<zQ8=�O=\;=�a=�6�<��%�ଭ�����WP�N-r�tO}�D�p��M����������ti�<�H
= O<=�   �   ��;=B+=�»<�N��Vp���<����A��T��l����̿��Ȇ&�ZYL�h�u��Ə�3����A������<����������Mv��M�TZ'�tq��ο�r��5V�fS�_)��jc>�S]��`$����<fv*=d�:=*=,��<0��; -|� ����^�^���l���$ॽ잽����jO[�L����m�P�;�o�<�� =�   �   �"�<F� =���<t���粝��1�����	j�4CI�iҏ���¿N����l��A�n�g�@͆� a���������������?��������g��B���� �����ÿc�����J��Q��բ��2�co���S���i�< ��<��<| �<`� �x 㼨�a��맽��ؽ�n�������g�����%uֽ�E���\�85ڼ@tҺ��<�   �   @�};��\<З�;`&��#��n����u��7��ރ��n���(� ��1�r�R��/s�⷇��W��M����#��/k����r�,LR�z1�����I��Gi����8�Z��𒾜� ��=��X������;��T<�Q;�f���J��b��*5 �R'��/J�/�e��w���|�"Vv�\Ad�#bH��[%�����
	��F�E�$X���   �   |U�X�\�@��Ժ���΀��
��!}�U�ѾDI!��i�
���п�F� ���9�`aT�Pk��dz����*�y�2Aj���S��9��h�� �mпݱ���i���!���Ҿp\~���
����0���x�
�8�h�f������E����12���l�3���Ё�������b;M�Ѿ��̾���Q+��Z�����i�>�/�l�񽓑���   �   �����dP��^��` ���%i�8罠kR��w����e?F�+����J��+�>*��T�L�4�hOF���Q���U�htQ�zrE��3�Ȁ�:���l�"겿a����@F��-�Dί��S��1�tk�8��&���T�n�����|_�����
�¾���ng���� ��#�����#��n�g��<}��Q/��t \�i���   �   &���ͽj�x��s6��H]��漽�'��o��T�۾#�!��a�VԔ��컿h��������#��,�&�/�%,���"��0�Z&�Za� ����6���i`��n!��۾�b��<�'��m����^���8�R|�SVн(���|�C���9*뾓��y�0�aJ�j^�=4k�[o��j��k]�I�(2/�K6�����ï�5z��   �   Ɨ��@T'���ͽ>����c�X��� �n/V����Q~���1�� m�F���,ʷ��"׿��� ���
��/�F�
�z�!񿼝տ~��������k�7�0�^��>㨾ڋU������Ι�<�d�B"��ӰϽ�(��ɂ��L�������)���R�×y�d����U��}���yz���S��V��������w���P��P(�:\�c����   �   ����v���~���5��{}���컽�w�p�w��R��t���4���g�d^��J��� ���5�ο�vٿ��ܿ^�ؿ3�ͿV��SH���>��%$f��#3���7��d
v��������5��,��4񻽿{�B�w��V��9����4���g��`��B���J�����ο�zٿ<�ܿ��ؿ��Ϳ3Y��%K��-A��=(f�3'3�����   �   4b��"樾��U����_Й�X�d����v�Ͻ;�(�/Ƃ��G�������)�	�R���y������R��E���;w���P��R�����ƛw�m�P�M(�fY���������O'�Q�ͽ������c������ ��3V�`�������)�1��$m��▿ͷ�	&׿Y��~"���
�2�J�
��{��$�͠տ����4㕿�k��0��   �   �p!��۾�d����'��o���^�V�8�Z|��Nнn(���|�U���$�ߕ�/�0�P\J�Az^��.k��Uo���j��f]���H�./��2����:���6�y��&��ͽ�x�Jp6��I]��鼽ޭ'��q����۾��!�2"a�c֔�﻿\�㿄 ���4�#�d�,�v�/�T',���"�^2��'�d�L����8���l`��   �   �BF�d/�LЯ�rS�F4��k�p4�����T����ԩ���^�:�L}¾��뾯c����� �t#�d����k�����w���*��X\��{���LZP�|R��L���'i�� ��nR��y�����AF�ʫ���L��}-Ὸ+�FV�Z�4��QF��Q�4�U��vQ��tE��3�l�����6o��벿Έ���   �   �i�Y�!�ڑҾ�^~��
���h��� �
� �h�Z��@��� ����*2�^�l�J���M|�������\;��Ѿ��̾7����%��������i���/��񽋉���I�@�\�0��$����π��
��$}���Ѿ�J!�F i������п�G������9�xcT��k�Tgz������y��Cj���S�\9��i��!�п&����   �   j����8�����𒾒� �q>��T���p��;xU< �Q;�M��l�J�1Y��U/ �MK'�o(J���e�w���|��Mv�U9d��ZH�#U%����������tE��A�� O~;��\<`��;4&���Ï�&p�9��*w𾙫7��߃��o��/*����Z�1��R��1s�����X������%��El����r��MR�.{1�� �=��R���   �   褐�U�J�(R�-֢���2��o��pQ��0o�<x��<���<$�<�������a�,㧽��ؽud���������a��y��lֽ�=��B�\�Dڼ PѺ���<-�<p� =�Ď<<���2���:1������j�YDI�-ӏ���¿�����m��A���g�Ά�b������������[@��M���g�fB��������U�ÿ�   �   �r��~V��S��)���c>�F]���"����<�x*=v�:="=$��<�;�|�ܖ���^�����`���ۥ�瞽ُ���F[�����m��2�;\x�<0� =��;=�+=�û<P��Mq���<�Ϳ���A���T�m����̿l��<�&��YL�&�u��Ə�����&B��/����<�� ��I��@Nv�" M��Z'��q�9ο�   �   e!����Y���Y�����B��鬽`'���r�<R8=x�O=�;=�a=|7�<`�%�D���b���WP�(-r�hO}�<�p�&�M����l������i�<<H
=�N<=<OP=��8=�<DN��몽s�@�
B����O`X�����+п����W)��P�V�z����������Q��`����U�� ̥��0��|{�hQ��G*�����ѿ�   �   r��{V��R��(��Ib>��[��H����<�y*=�:=�=���<��;(|������^�v���O���ۥ��枽ʏ���F[����H�m�P4�;�x�<�� =~�;=t+=xƻ<�K���o����<�۾���@���T�ul����̿����&��XL��u�1Ə�����A��!����;�����x���Lv�(M��Y'�q�Wο�   �   ����k�J��P�XԢ�D�2��l��PI���t�< ��<L��<��<�����⼢�a� 㧽h�ؽYd�����x���a��y���kֽ�=�� �\��ڼ�?ѺD��<H/�<� =�Ɏ<P�������1�Н���i�vBI��я��¿m���@l�*�A�`�g��̆�M`��������������>������D�g��B�0��������ÿ�   �   Ch����8���m9� �:���욼p��;PU<��Q;�K����J��X��2/ �,K'�R(J��e��w���|��Mv�D9d��ZH�
U%�{������� tE��?�� h~;�\<��;0��P����l�� ��ws���7��݃��m��K'�,��~1��R�,.s�϶��VV������"��	j��Ʀr��JR��x1���J������   �   ��i�/�!�h�Ҿ�X~�"�
����ܬ��X�
�X�h�j������{����*2�0�l�7���;|��|����\;�Ѿ��̾.����%��������i�}�/���� ���H� �\����ث���ʀ��
��}�N�Ѿ�G!�i����}	п�E����l�9�j_T��k�bz�@����y��>j���S�9�&g����пX����   �   9>F��+��˯��	S��+轐k�
-������T����t����^��0}¾��뾤c����� �m#�^����k���龵w���*��)\��{� �PWP� I������i��RhR�:u��
�<=F�����#I���(��(��R�X�4�&MF��Q��U��qQ�&pE��3�����j�貿�����   �   8l!�B�۾ `�� �'�Mg����^�Ԯ8�p|��Lн�(���|�/����#�ѕ�"�0�E\J�7z^��.k��Uo���j��f]���H�./��2���"�����y��&���ͽV~x�i6�t>]��༽f�'�%m���۾��!��a�tҔ�<껿���0������#�ܘ,�ց/��",���"��.��$�g^�󺿹4��xf`��   �   DY���ߨ���U�����&ș�h�d�3��$�Ͻz�(��ł��G�������)��R���y�~����R��B���8w���P��O�����w�h�P�M(�\Y�򋼾n���?O'��ͽ�����c������ ��*V�삩�z��5�1�m�ޖ�Ƿ��׿A�����
��-�<�
�(x��񿄚տF{���ޕ���k��0��   �   ����v���c���m.���x���黽�v�Ǜw��R��`����4���g�^^��E�������1�ο�vٿ��ܿ\�ؿ2�Ϳ
V��QH���>��!$f��#3������	v�Č�����(0���w��滽�s���w��N��ښ��}4�l�g��[��n���Ϗ����ο4sٿ��ܿ��ؿ��Ϳ�R��`E��%<���f�U 3�>���   �   ����hJ'�Բͽ������c����� ��.V�˅��"~�� �1�� m�@���'ʷ��"׿��� ���
��/�F�
�z�!񿼝տ~������z�k�.�0��]��㨾�U������ʙ�>�d����̢Ͻ,�(����C��Ά�F�)��{R���y����O������s��qM��>���0����w��P�NI(�WV�H����   �   �&�Տͽdtx��c6��=]��⼽��'�$o���۾�!��a�OԔ��컿c��������#��,�$�/�%,���"��0�Z&�[a� ����6���i`��n!�ږ۾lb��"�'�^j����^�N�8��{�Fн�(���|������G�� �0��WJ�%u^�~)k�7Po�4�j�oa]��H��)/�/�Ҹ�@���j�y��   �   k鸽RKP�:������i�Z罷jR�:w����[?F�'����J��+�<*��T�L�4�fOF���Q���U�jtQ�zrE��3�Ȁ�:���l�"겿a����@F��-�ί�&S�/轾k�+����$�T������l�^��엾�w¾e���_����� �$#�$��z�Kg�Q��r��&���\��u��   �   8;���\����4���?ˀ��
�!}�"�Ѿ6I!��i����п�F����9�`aT�Nk��dz����*�y�2Aj���S��9��h�� �oп߱���i���!�ҏҾ�[~���
�:��<���`�
� �h����}�������#2��l�x����v������sV;��ѾY�̾>���u ������V�i���/�d��^����   �   ��~;X�\<���;,�������m�����t��7��ރ��n���(� ��1�r�R��/s�⷇��W��M����#��0k��¨r�.LR�z1�����M��Gi����8�?���ޡ ��;���욼��;�$U<@9R;5����J��O���) ��D'�� J�ڗe�w��|�Ev�#1d�@SH�bN%��������zdE��'���   �   �:�<@ =�Ύ<<��b���r1�h��� j�/CI�iҏ���¿M����l��A�n�g�@͆� a���������������?��������g��B���������ÿd�����J��Q�qբ���2��m��0J��4w�<d��<D��<  �<`K����a��ڧ�X�ؽpZ��p��*���\��o���bֽ<5����\��ڼ к�
�<�   �   v�;=�+=Hɻ<HJ���o��ʧ<�����@� �T��l����̿��Ȇ&�ZYL�h�u��Ə�1����A������<����������Mv��M�RZ'�tq��ο�r��4V�cS�Q)��0c>��\��������<�z*=T�:=�=L��<P�;H�{�*��4�^���h����ե�➽
����=[����h�m� c�;���<h� =�   �   ګh=�R=�=�У��.��>�'�|7���� �LXD�f������� <�����T=��a�8���I��J��m0���N���d��Mz��@�b��>�����;��J��ٍ�`F��M��:���a*�������Ȼ��=`�O=��e=BzR=�N#=$��<a�;0�/�X�ռ�b���;�N�E���9�x����̼�Z�X� <�g�<b�'=�V=�   �   ��U=�
F=H��<@������l$�@�������@����L{���J�Z���9��n]�2����������	���k������:���^�(�:��O�#������Z����B�=���p�&��a���w̻���<�B=�LR=le8=��= �g<����8ȼ��)�`V`�1b���]T��>�\���$�8���H��n|<h�=I<=�   �   �E=h�=��<����0>|��h�l����d�6y6�{��_f���翖��u0��^Q�
�q�@	���������(���t��&�q�x�Q���0���+$�Ü�����~8���cm������5�� �߻�r�<rG=�C=`��<���;�҈�HF,������&��n�ٽ���e;��F��W!׽�첽�`��>%��w���<��<�   �   �W<�f�<�Ɔ<P��� �b�hL	��}���ؾ�R&��(p������տZ���A"�dX?��l[��{s�L��[���\���^�r�H�Z�6?��@"����zֿXդ��q��x'���پ�͂��*��5h� �p ~<���<P2C<x^	�6"�Ő���ڽHG��Q1��J��sZ���_��Y���H��/������սx7��2R���߻�   �   d��� �C� ,	;��?��G����r_����b��!�S�+���˨���￶��&�)���@���T�V�a�|f�*
a���S��@���(�:;�3��p���N���?�T��v��&��RDa�hW�'L�ȏO�@Q�:PƊ���ͼF0p���нGQ�-.Q� ڂ��>������tO�����t���2g��6�����f�M��$��S˽��g��   �   a��P��<������@�1��e½�d8�����mS����3�y6y�����οQ�����8%��4���>�$7B�M>���3��)$��+�R����Ϳį����x���3� ���3��o9��EĽ|)5�$��� }��h4 ��������&�D��p�����a�Ծ�\��-w��������_�������IҾ~��TE���@�� ��   �   q�3���P�?�(�P-'�s˛��C��3y�~ž�c���L�1쇿T*��:ѿ�K����	���:��>� ��v�08�*��`_�
Ͽ?���:��T�K����Cž�Ky�|���՜���)�����D�)>�������_�w��'�Ӿ���> ��7��lJ��V���Y��cU�M(I�[K6�v�������оz���*p\��   �   3�d�~��l.����N�:�-�J:w���ٽO!<�x_����㾓!�Q�W��މ��b���mſ�޿����!��,��WH��0��ݿ��ÿ�⦿�����QV����)L�>���a�;���ٽd�w�,h/���Q��������m�g�����ã����u?���c�����M���F����5���=��u��T���~:a��R=�?+�\��i����   �   rX���&Y�dP�-D���cH��	I��S���Z��Z�ʧ�(2�>�#��:S�e��]V������m����{ǿ?�ʿ��ƿ�g���N���ߗ�ᵀ��Q��)"����U���!Y�^M��@��TbH��I�X��<^�l�Z��ͧ�A7��#��>S����Y����������ǿ��ʿ��ƿ�j���Q��#◿$����Q��,"�t���   �   �O�鳖�؃;�{�ٽ>�w�nf/�J�Q�����8���g�p���-�뾜��dq?��c�R���q���L����2���:�����Æ���5a��N=��'�+��r���l�d����q)����N���-��>w���ٽY%<�}b����m	!���W����� e���pſp�޿��%����L��{3��ݿ��ÿN妿
����TV�H���   �   ���Fž�Oy�����ל�\�)�ʛ�ȰD��6�������_����}�Ӿ���: ���7�hJ��V���Y��^U��#I�G6��~�~����оA����i\�bl�ѩ��z�?���H.'�3Λ�~F�8y�d�ž�e���L��,���ѿ�N����	���D��N� ��x�:�ؽ�Rb򿒁Ͽ`��J<��
�K��   �   ��3������4��Xq9�HĽ�)5������n��4) �����H��$�D��l���|��;�Ծ�U��rs������\������e�Ѿw��2A����@�� ��Y��x�L1�������1�i½�g8�����V����3�v9y����T�ο����Z:%���4���>�^9B�*O>���3��+$�^-�Ѱ��)�Ϳs���.�x��   �   �T�Ix��(��mFa��Y��'L�p�O� ��:p���ԭͼ" p�D�н�J�j&Q�|Ղ��9��B����I����Ú���a��M�������M����I˽��g��z�� >C� l	;8�?���G�B�뽺u_������G�S���������� ������)�R�@���T���a��f�ba���S��@��(�b<���󺾿����   �   `�q��y'���پ�΂��+��6h�h�/~<��<�TC< 1	��������ڽA�K1�yzJ�lZ���_�DyY�s�H��/������ս�.���D��U߻8�W<�p�<�ˆ<p�����b��M	���~ؾOT&��*p����W�տB���B"��Y?��n[��}s�[��p���d���6�r���Z�t?��A"���|ֿM֤��   �   H��.8�����m�����5�� �߻�w�<fK=zI=���<���;P����8,������ٽ��ｉ1�����9׽�䲽�Y���
%�P�v��<��<:J=f�=Ш�<`����@|��i�h�:f�Ez6�/��Cg����D��v0��_Q�Z�q�
������^������*��T�q�h�Q���0�n��%�h����   �   [��޵B������(�&��a���q̻���<<�B=�OR=.i8=>�=H�g<0߭��)ȼ|�)�jM`��]��Eꆽ�O���{\��$�8
����(�|<`�=2L<=ʢU=:F=$��< �����:$�������1�@�]���{���K�[�4�9�Xo]�����)���������ٶ��!�������^�~�:��O��������   �   �؍��_F�vM��:��Na*�<����Ȼ0�=��O=�e=�zR=�N#=���<�c�; �/���ռ�b�\�;�8�E���9������̼�[��� <�g�<�'=PV=��h=��R=�=P֣�k/����'��7���� ��XD���������'<�����l=��a�&8�� J��J��m0���N���d��Bz��(�b��>�����;���I���   �   xZ���B�C����횾��&�`��@a̻D��<$�B=4PR=�i8=��=P�g<0ݭ�x)ȼR�)�DM`�q]��6ꆽ�O��~{\���$��	��`����|<��=�L<=T�U=F=���<����$���ǻ��H�@����{���J�lZ�`�9�Fn]�煀�Z��:��������N��ձ��v^���:�0O�w�����   �   ��g8���@l����3����߻�|�<M=�J=���<��;4���b8,�������ٽ���o1�����"׽�䲽�Y��P
%���v��<D��<BK=��=���< ����:|��g������cx6����e��5���0u0��]Q���q����뮐����Q��������q�`�Q���0�0��
#�؛���   �   �q�Xw'�u�پr̂��(��.h���@=~<`	�<[C<0,	���������ڽ�@��J1�`zJ��kZ���_�0yY�b�H��/����^�ս�.��D�`N߻ �W<u�<�҆<�q����b��J	��|��ؾ�Q&�G'p������տ����@"�.W?�\k[�,zs�F��H���M���j�r���Z��	?��?"���Iyֿ#Ԥ��   �   �T�\u��$���@a�.R�2L��mO���: m���ͼ�p���н�J�:&Q�fՂ��9��3����I���������a��B�������M���|I˽��g��w���C���	;H?��G���Ap_�������X�S�����N����ￒ��)���@���T� �a�. f��a���S�.@�$�(��9��������   �   q�3�����|0��`k9�!@ĽP5��{���e�� & ��������؀D�dl���|��$�Ծ�U��hs������\�����Z�Ѿk��!A��R�@�� ��X��� ��(��0ힼΗ1�*a½�a8������P����3��3y�&�� �ο���x��6%���4���>��4B��J>���3�($�N*�������Ϳ߭����x��   �   O�l@ž�Fy�����Ϝ���)�����D�f5��I����_����Z�Ӿ���: ���7�hJ��V���Y��^U��#I�G6��~�x����о.���yi\��k�p����?���#'�9ƛ��@�R/y�{ž�a���L�tꇿ3(���ѿ�H��0�	���8��0� ��t�F6�j��C\�R|Ͽ����8��I�K��   �   �G������{;��ٽ��w�6\/���Q�x���|����g�@����뾋��Sq?��c�M���l���G����2���:��������5a��N=��'���U����d����_'���N��-��/w�w�ٽ<��\��Ȉ��!���W��܉�`��kſ��޿ ��&��H���D��r,�ݿ��ÿ<িµ���MV�����   �   Q��Y��H��9���UH�p I��P���Y�t�Z��ɧ��1�-�#��:S�_��XV������h����{ǿ?�ʿ��ƿ�g���N���ߗ�ീ��Q��)"�����T��n!Y�oL��=��8YH���H��M���V���Z��Ƨ�\-�&�#��6S����S������8���Oxǿҡʿ>�ƿkd���K���ܗ�����Q��&"�����   �   ��d�l���!����N��-�*2w�J�ٽr <�0_����㾂!�A�W��މ�zb���mſ�޿}���!��,��WH��0��ݿ��ÿ�⦿�����QV����
L�����;��ٽn�w�\/���Q����������g�L���՘�G��_m?�mc���������U����/���7��������)1a��J=��$�������   �   �f�F����?�D�.#'�ț��B��2y��}ž�c���L�+쇿O*��6ѿ�K����	���:��>� ��v�08�,��b_�
Ͽ?���:��R�K����Cž*Ky�t��`Ҝ���)�v��d�D�/�����,�_�����ӾQ|��6 �W�7�ZcJ��V���Y��YU��I��B6��z�����о�����b\��   �    Q���������枼�1�=c½d8�|���DS��v�3�m6y����	�οN�����8%��4���>�$7B�M>���3��)$��+�U����Ϳů����x���3������2��Hn9�SCĽP!5��w��HZ��X �S������DzD�>h���w��7}ԾO���o�(�����3X�6��9��H�Ѿ4���<��k�@�N ��   �   �_�� �B�@�	;�v?��G�	��Hr_����S���S�(���Ȩ���￴��&�)���@���T�V�a�|f�*
a���S� @���(�:;�5��s���O���?�T��v��&���Ca�mU�� L��jO����:p3��\�ͼ�p���нxD��Q�т��4��ϛ���C��?
�� ���V\��A���.��D�M�d�;?˽��g��   �   `�W<̀�<�ن<pf����b��K	��}��tؾ�R&��(p������տZ���A"�dX?��l[� |s�M��\���\���^�r�J�Z�6?��@"����zֿYդ��q��x'�i�پ�͂�*�`1h���G~<$�<@yC<�	�*�=���owڽ�:�$D1� sJ�'dZ���_�`qY��H��/�����~ս�%���5���޻�   �   �P=��=L��<@���T;|�*h�I����d�1y6�y��\f���翖��u0��^Q�
�q�?	���������(���t��&�q�z�Q���0���-$�Ĝ�����|8���Bm����@4���߻T�<P=HO=��<��; ����+,�2舽t����ٽ>�ｮ'�����׽ܲ��Q���$���v��+<���<�   �   �U= F=X��<�맻���6$�0�������@����N{���J�Z���9��n]�2����������
���j������9���^�(�:��O�$������Z����B�7���cД&��`���f̻���<N�B=JRR=�l8=��=0�g<�����ȼ~�)��D`��X���冽'K���r\��$�\���䀻��|<�= P<=�   �   �<�=��t=
c.=Б<$?A�X;�rV��G޾!%+���v��f��',ۿ-	��x&���D��jb��|�ކ��������G|�z�b�r�E��m'�x3
�ݿ���(�y�I-��yΆ��������K���;��&=�m=�T�=�zo=$E=,"=�)�<��.;؉6�8����뼌^����A��������;Ȱ�< �=�wM=`�w=�   �   V:w=i=�H(=X[<Z�;����������پB�'�L�r�+�����׿�����#��SA��^���v���[
��8���^w�l^��A��$����Dnٿ�,��Pu�g*���ܾ�����F�&�E����;� =�ja=�Jo=��W=��&=�o�<@�;����˼8���-5�6�>�.{2����8�� ���`�<�=�<l�/=xV`=�   �   �qB=�E=�$=�&<� ,��.����r�x;;A��@f�=w���mͿ� ���r7���Q�d�h�L�w�B^}��w��Th���Q���7�VI��@���οt����h��� �d�Ͼ�v�Q���c5����;��=ʷ==:=�=\��< �2�LEм� C�wщ�_���8��|ý���\]���Å�B�9��.�� ��\�<�=�   �   ���<^j=TU�<���;���a�ڽ�zY�"����~��VR�����M��p����v(�ƾ?��ES�b`���d��`�\�R��@?�4(���b������kc����S� ��g���0�\�b�߽��� ��;�k�<���<(�<���;���Q� [��vu�ٲ��(��6�/�:��5��&����u����:�D�|/���n�;�   �   �� ���+<�uu<��%;���P.���:���������29��#��动��Կ�H ����)��:�n�D�_H�XOD��S9��)�_�����r�ӿ�����l����9�1������K<�$���b�� �g:@iX<0�
<pe(��%������q���.�=�\�a��.Y��Ԣ��#젾R蜾���PK����X��*�)����Κ��R��   �   �ZY��P����r� e���}ռ.˓���������Ӿr���Z�Ѱ��Z䶿X�ݿ���>@����n(��*�4�'����G�� ��ܿ����O��UZ�p���"Ծ�����1n��M�`Ļа�����Nd���н�"���d����ɶ���ԾL�N(������$���o��TҾ[���j���`�&��?ʽ�   �   ���|����dł���ü`Ec�V���5Q��<�������2��n����� ���ؿz��������*�8~��G�y��<�ֿ$���%閿��m�n2��������oQ�����^f���˼�ꌼ���ɂ����O*;�*]���1���%��Q��^ �@�0�e6;�0�>�<�:�R�/�8��ۅ	�ĭ㾚 ��FՄ�$27��   �   �>�p�z[~�H����мBL*�yg��R��j���þ��B�<�[ir�j���"�����ſ�B׿�Z⿲�� ���տ�ÿ��� !��J p��F;���
���¾�s�@��2��Ze+�H�ռ��	�h.�����0"B�Đ���E˾w��'��LG�+�c�9�y�/у�,��KV��	x��wa�[�D���$�w���PȾZ���   �   󁍾h�4�%�ҽ~�`��� �l�~rc��ս��6�?���%о�j�D�8�``d����<l��
�������|X��䯿��������¾a�+�6�����;�~��3�4���ҽ��`�� ��n��yc��ս>�6����V*о�m��8��dd����n�����������[��篿�������Z�����a���6������;�   �   �¾�x�X���5���g+�4�ռ�	�:)����콊B�򌑾�@˾`��`'��HG�e�c��y��΃�y���S��x�]sa�D�D�B�$�����KȾ�V����>�i轈R~�֠�4�м0P*��k���!�<m����þ�����<�Xmr�Ŝ��ո����ſF׿D^���h���տ��ÿ?��6#���#p��I;��
��   �   7����'sQ����.bf���˼⌼������ѧ� $;�$Y���,����AN��Z � �0��1;���>��}:�-�/�k���	�	������ф�n,7�ǣ彆�|����@���0�üBJc�(�齾9Q��?��������2�w�n�3���#���ؿ7}��N�`��z,���2I�s����ֿl���떿��m��2��   �   5��8%Ծȡ����p���M��ĻP~��褺��?d���н��"���d�"���ö�ؼԾqE�^!��������i�OҾ#��4f��,�_�V��Xʽ�MY� ?���br��V��̀ռ�͓�v��������Ӿ|��ȌZ�����e涿��ݿ����A�l��F(���*��'����"I�k� �:�ܿ���Q��vWZ��   �   y�9�{�������M<����6�� 9h:�{X<`�
<8:(�(�$�@���f���.�9�\����NT�������栾E㜾����F����X�� *�J���ƚ��E��� ��+<��u<@�%;p��� 1��:�����Ǘ���39��$��t���jԿJ �����)��:�F�D� aH�(QD�HU9�\)�V`�����#�ӿR����m���   �   �S���������\���߽X����;Dr�<���<x�<@��;蛪�Q��Q��hj꽪��(��6��:�5�2&���/k�����D�8�����;0��<�n=Z�<��;2����ڽ�|Y�Ӈ����pXR�-����N���q���x(�$�?�TGS��c`�r�d�p`�عR� B?�$5(���������Gd���   �   �h�X� �6�Ͼ�v�T��bd5����;��=L�==
$:=l
=��<�!2�8-м��B��ɉ��V���/��Xsýn���:U��l����9���� B�����<�
=�uB=ЇE=�%=h%<�,��0��M�r��<;1���f�
x���nͿ�� �����r7���Q���h���w��_}�\�w��Uh���Q�^�7��I�ZA�l�ο����   �   �u��*��ܾ����
G��E�0��;D� =�la=�Mo=8�W=��&=�y�<PI�; ����˼0���%5�Ⱥ>��r2���	���y��0�<�F�<�/=FY`=N<w=2i=ZI(=(Y<�;���������پ��'��r�����@�׿:��d�#�~TA�:^�t�v�h���
�������w��l^�p�A�*�$�����nٿ�,���   �   �y��H-�\yᾆ���B����K���;F�&=`	m=U�=L{o=rE=t"=D*�<��.;؈6�Ԥ��P�T^�����A��������;l��<�=ZwM=$�w=�<�=R�t=�b.=X�<�?A��;��V��OG޾R%+���v� g��K,ۿ,-	�y&���D��jb��|�ކ��������G|�h�b�^�E��m'�d3
��ݿ����   �   �u��*���ܾ齃��E�>�E���;t� =nma="No=��W=$�&=�z�< K�;0��<�˼
��b%5���>��r2�Ԍ�����x����<G�<>�/=�Y`=�<w=�i=�J(=0`<8�;����K���u�پ�'���r�񛥿[�׿�����#��SA�$^�,�v�����	�������
w�zk^���A�p�$�$���mٿ",���   �   �h� ���Ͼ��v�Q��_5� ��;<�=�==2%:=F=d��< 2�8,м~�B��ɉ��V���/��;sýR���!U��T���ւ9�@�� �����<V=�vB=:�E=((=�2<��+��,��X�r��:;���j f��v���lͿz� ����Vq7���Q�F�h��w��\}���w�DSh�z�Q���7��H�A@���ο�����   �   �S�߷�������\�d�߽���0)�;�x�<P��<��<��;���FQ�5Q��j꽈��� (��6��:��5�"&���k佦����D���`��;���<�p=4`�<���;����ڽ�xY�ф���}��UR�F���tL���n�̣��u(���?�PDS�d``� �d�`�ʶR�|??��2(���������Tb���   �   ��9�I�������H<�c���^����i:��X< �
<p2(���$������e���.��\����>T�������栾:㜾����F���X�� *�����Ś��D��� �X�+<0�u<�F&;T����*��!:���������i09�r"�������Կ�G �\���)�8:���D�B]H��MD��Q9�f)��]�������ӿ^���tk���   �   Z���Ծݝ������h��|:�@�û�[������=d�'�н��"���d����ö�¼Ծ\E�K!��������i�OҾ��'f���_�*���
ʽ�KY��9��@#r��%��nռ�Ɠ�,�����Ӿ�����Z�Q����⶿!�ݿN���>����(�>�*�^�'�(��F��� ���ܿ����M��`RZ��   �   z�����PkQ��꽤Sf� �˼�Ԍ�$���4���˦뽼#;��X���,��h�2N��Z ���0��1;���>��}:�'�/�f��z�	�������tф�,,7������|����в���ü�;c�{���1Q�':�������2���n�3���S��z�ؿw��������(�v|��E�`��q�ֿ����疿"�m��2��   �   ү¾n��{�U+���Y+�lwռ��	�'�����
B���l@˾N��P'�vHG�Z�c��y�΃�v���S��x�Zsa�A�D�>�$�����KȾ�V����>��g转N~����мdB*��a����g����þ���<�<��er�-���������ſ�?׿�W�T��ω���տ�ÿ������Pp�wC;�(�
��   �   n{���4�ßҽ��`�ڙ �vc��lc�� ս�6�	���%о�j�5�8�S`d����6l���������yX��䯿����������a�'�6���}�;�~����4��ҽ@�`� �&b�$gc���Խ��6�	���!о�g�ֶ8�C\d�7���i��*�������fU��᯿�|��g�������}�a���6�-����;�   �   ��>��_�PD~�����м�D*��d����Ij����þ��2�<�Nir�d��������ſ�B׿�Z⿯�����տ�ÿ���!��H p��F;���
���¾ts����/��^+�$wռh�	��"������B�C����;˾f���'�ZDG���c��y��˃�� ���P����w��na��D���$�|���FȾS���   �   ��.}|�(�4�����ü?c�C��*5Q��<�������2��n����� ���ؿz��������*�8~��G�z��<�ֿ&���%閿��m�j2����p��BoQ���꽺Xf���˼(ό�`�������|��	;�;U���'�����J��V ���0��-;�3~>�hy:���/���� 	������~̈́�&7��   �   �=Y��%��@�q�����nռ�ȓ���d���}�Ӿe���Z�Ͱ��U䶿T�ݿ���<@����l(��*�4�'����G� � ��ܿ����O��UZ�k���"Ծ柅�V���k�� >���û�2�������0d�G�н��"�V�d����K���϶Ծ�>�m���������b��HҾ����a��e�_���Nʽ�   �   � � ,<h�u<`f&;����i,���:�t���ߔ���19�|#��㊨��Կ�H ����)��:�p�D�"_H�ZOD��S9��)�_�����u�ӿ�����l����9�"������DK<�K������ �i:��X<��
<(�x�$�����Z��.�S�\�p��yO�������ᠾ+ޜ�=���}B���X��)���������r6��   �   ���<*v=�f�<���;̤�	�ڽTzY�����~��VR�����M��p����v(�ƾ?��ES�b`���d��`�\�R��@?�4(���d������kc����S���N���Ҙ\��߽d��0)�;H}�<$��<@�< 4�;�����P�H��y_꽈��b�'��6���:� 5��&���'`�@
����D�������;�   �   �{B=��E=H*=P6<8�+��-��J�r�f;;<��<f�;w���mͿ� ���r7���Q�d�h�N�w�D^}��w��Th���Q���7�VI��@���οv����h��� �V�ϾƖv����:a5����;b�=��==f):==���<��1��мB�B�(�~N��\'���jý�����L��Ĵ��Bu9����� ����<�=�   �   D?w=�i=�K(=�b<�;����p�����پ>�'�J�r�+�����׿�����#��SA��^���v���\
��9���^w�l^��A���$����Enٿ�,��Qu�g*���ܾ}����F���E�P��;Ĉ =|na=�Oo=j X=��&=p��<�u�;8��D�˼l��X5�v�>��j2���`����D����<�P�<P�/=�\`=�   �   0Ȗ=��=p#^=���<(!ƼE�ɽ�US��Ŷ�*���RP��P�������^�,n�N'��_>�PR��R_��d��Z_�v'R���>��'�:3����G���ΐ�%�R����l	����X��ҽ��L�<�XM=�S�=���=�m�=Fh=`6=d��<�F�<�!�;@nm��`���4���@�����< 6�<�=xYF=�ry=A\�=�   �   !*�=��=\�X=У�<����8)Ľ{�N��
���8�D�L��ጿ����`���%�jY$�r
;�FN�[�f�_��[��.N��I;���$����� �%��wC����N��'�p&����S�J�̽ݼ���<l'H=/L�=uS�=�cx=��M=��= ��<���;�#λp��d��@iʼ�����q���z�pA"<T�<�Z&=zQ_=J�=�   �   "�o=RFr=��G=D��<���#��V�@�6:��X\�d�A�Ʌ�����ðܿ؇�R^�6�1�.C���N�f�R���N���B��|1�F�����״ݿ����sކ�8�C�����檾E��
��X����h�<(�7=R�a=�u^=��9={�<0�M<�� �ռ�<0��Kf��	��.'����J�^��M%��غ�@�S���<�X=��K=�   �   TH=t;=�(=H?�<h}x��Л�e+�f��%�}�0��=u�e����~˿�f�����#�H�2��<�L@�؈<�F+2��"�z���o��?�˿�)��ݗv�V2�ֆ��v����.��{���p����<Jg=޿+=�}=X�< ?S��-�$[i�n����ܽ�\�Z����(��4��
Bֽm!���gX�q̼��:�V�<�   �   �b#<�E�<`��<�ș<��(�b�|�$9�<.����о��ėX��s��|`���ܿƙ ��8����v '���)���&�j��ƕ�� �Qmۿ +��C����Y�����fҾ2����������`!T���<�\�<���<��;���J�Z����.��<�.�j6R��n��� ���:~��6k�4dN��D*����̱�v�G�Ȣ���   �   �� h����Y< �K<��ѻ�`>��R���T��ޭ�����7��[u����a὿f@޿t������������]����E?��w�ܿqӼ�eN��¶t�`�7�����p���qV�@�轄�E�p�P6$<�A+<�S���;����A�����5�$=q� r��4���2þv�Ͼ;�Ӿ��ξ�b��T���̬���k��d0�j�L���   �   �<�� ���� ~;�$������멽kp$������Ҿd��q�I�����靿�q��K�ѿ�T��!�����[�S����Ͽz緿K���
��|TH�W�}|Ѿ�~��I�$�s��d����˻ ��9XS;�b$�OϬ�6�нY�����d߾�h��������2�����.E�����G���th���Ǒ�r4T�dm��   �   �R�{%�� ����J�0�̻v�� We��*�sM�Q���?���_�_�L�Q.|��Ԕ�1����1��:�����Ŀ�1��� ��KH���Z���y�؏J���֗澙`���L����e�|񩼐�黠�`���"�煭����*k������ ޾���^'��?�4�R�_���b��)^�qQ���=��4%��	�|\ھ�����kf��   �   �wc�T��q敽�x��p=�HzA�����������ڥf������ ���z@�}�d��I��r����l��t䘿�ᕿ���0���b�K>���~���ը��rc�����ᕽ�s�xk=���A�қ���������f�_ ����>��c~@�Ǻd��K�����vo��"瘿=䕿����z��� b��>����"��q٨��   �   �c��L�x��� e����������`���"�������k�����]�ݾ����Z'���?���R�g�^�E�b�=%^��lQ���=�1%��	�~Wھ�����ef�^N�U��8��P�J�P�̻�|��`^e��0�xM�������辖b�ҠL�j2|�ה������4�� �����Ŀ�4��]���J���\��ޘy��J����̛��   �   �Ѿŀ��&�$�tv��d����˻ ��9�6;��V$�kǬ����Y���5ھ�_��q����_�����fA����|D��侈c��Ñ� .T�vh�}5���h��@�;P)������墳�s$�4���P!Ҿ���d�I�`���띿Dt����ѿ�W��$�����^�%�⿂�Ͽ�鷿K������,WH�m
��   �   ��s��rtV������E���P@$<�W+<���J/�7�������1�5�5q�tm�����N-þ��Ͼ3�Ӿ��ξ]��@���Q��� xk�p^0�`������@n��`�Y<��K<@�ѻne>��V�e�T�{᭾����7��^u�����y㽿�B޿!�����N��V�z_�b���A����ܿcռ�P��d�t�n�7��   �   P���hҾ�����������H$T���<e�<�	�<�_�;����>�Z�7���@��\�.��.R�z�m�"�������~��.k��\N�:>*�E ��ñ�n�G�������#<0Q�<Щ�< ʙ<��(�4�|�D;��/����о} ��X�Pu�� b���
ܿ� �:����!'�r�)�(�&�������� �oۿ�,��u���� Y��   �   w2�p��x��ׯ.�3}��@r���
�<j=��+=`�=0%�<`�R���Ji�屫�Z~ܽ4W�T��
��"��)���7ֽC��XX��V̼ `�:tg�<ZN=x;="�(=�?�<H�x�4ӛ�I+��g��''���0�^?u������˿-h����#���2�j�<�bM@� �<�r,2���"�X��.q��p�˿�*��^�v��   �   ��C�e���窾�E����8���xj�<�7=h�a= z^=T�9=���<��M<����ռr/0�4=f�T���������6�^��@%������S�Ě�<4_=�K=��o=�Hr=,�G=؍�<���U%��ђ@�W;��&]�x�A�1ʅ�����˱ܿt��_��1�C���N�l�R���N���B�D}1���4����ݿ1°��ކ��   �   B�N��'��&��֖S���̽�ݼ���<�(H=M�=�T�=�fx=V�M=��=���<���;��ͻt�������ZʼL����q��,z�XW"<�]�<�^&=�T_=��=+�=Q�=ĭX=���<0���l*Ľr�N����C9��L�5⌿b������>&��Y$��
;��N��[���_�*[�/N��I;�@�$�
��	!�o���C���   �   ��R����0	��C�X���ҽ\~�`�<&YM=�S�=���=�m�=�h=�6=��<G�<�#�;�jm�P`�H�4���������<�5�<�=fYF=fry=*\�=Ȗ=��=#^=���<�"Ƽ��ɽ[VS�ƶ�S���RP��P�������^�>n�`'��_>�\R��R_��d��Z_�l'R�|�>���'�(3���G���ΐ��   �   F�N�	'��%��x�S���̽ ݼ���<�)H=sM�=�T�=Ngx=��M=B�=��<���;@�ͻ(������hZʼ�����q� +z��W"<�]�<�^&=�T_=��=8+�=��=ЮX=��<t����(Ľ�N��
���8���L��ጿ�����翪%� Y$�
;��N��[�ؕ_�[�.N�I;���$�p�� 鿠��	C���   �   �C����媾J
E�����p�<:�7=�a={^=:�9=��<�M< ��,�ռ/0��<f�/��t�������^��@%�,����S�p��<�_=��K=��o=
Jr="�G=���<����!��F�@�w9���[���A�Ʌ������ܿZ���]�~�1�TC���N�b�R���N���B��{1������Ƴݿ�����݆��   �   �2����`u��:�.�Rx��(e����<(m=��+= �=�'�< zR�0��Ii�����~ܽW��S��
��"�{)���7ֽ���WX��U̼�q�:�h�<�O=�y;=��(=�G�< lx�wΛ��+��d��v#�a�0�<u�u���o}˿!e�����#�"�2���<��J@���<�*2�ر"����n����˿�(����v��   �   <��_dҾ^���?��ǅ��T��)�<dl�<�< o�;���Z�������,�.��.R�Z�m�������w~��.k��\N�$>*�, �Yñ���G�����@�#<�U�<|��<ԙ<�t(�Ж|�
7��,��}�оu��X��r��_���ܿ ��7�2��'�x�)�>�&������� �^kۿv)��㈏��Y��   �   ���Hn���mV�p��4�E�`�
��W$<�g+<����F-�m��������5��4q�Ym�����9-þq�Ͼ$�Ӿ��ξ
]��6���D����wk�N^0��_������$��СY<��K<0�ѻ�X>��M彲�T��ܭ�\����7�HYu�i���t߽�*>޿����.��H��@�t\�����<���ܿXѼ��L��ʳt��7��   �   �xѾ�{��^�$�m���v���˻ ��9p&;�T$�bƬ�����Y�d�ھ�D��d����W�����^A����vD���|c��oÑ��-T�7h��4��������;�嚻<��]橽m$�j����ҾJ����I�����睿�o����ѿ�Q�������X�p��?�Ͽ巿+���:���QH����   �   <]���L�����e�Pݩ������`���"��}��g��Dk�o���:�ݾ����Z'���?���R�_�^�?�b�8%^��lQ���=� 1%��	�qWھ�����ef�N�;������lJ�p�̻|d���Le��#��nM�D���3��/]��L�n*|�hҔ�����+/��\�����Ŀ/�������E��BX���y�b�J�D��k���   �   �lc�$���ڕ�nh�hC=�h[A�N��꩘�H��o�f�X��������z@�s�d�{I��n����l��q䘿�ᕿ���0���b�J>���q���ը�rrc�4��)����n��M=� WA�~��[������K�f����N��)��w@�Z�d�.G��﨎�)j���ᘿ�ޕ��������yb��>����v���Ѩ��   �   0I�d������XJ���̻�h��jRe��(��rM�!����辺_�P�L�D.|��Ԕ�-����1��8�����Ŀ�1��� ��KH���Z���y�֏J���ė�y`���L���꽐e�d䩼 ��0�`�$�"��w����Ak�~���@�ݾ���>W'���?�]�R���^���b�� ^�YhQ���=�X-%��	�4Rھ����_f��   �   �,������@?;�ᚻ
���驽�o$������ҾU��d�I�����靿�q��I�ѿ�T��!�����[�U����Ͽ{緿L���
��yTH�R�h|Ѿt~����$�Uq���z�P�˻ �9�;�RJ$�?�����,�Y�X$վ�x����v�����ȹ��=�F��A��
�\^��0���	'T��b��   �   P�� ��ȷY<(�K<`�ѻ&\>�Q�w�T��ޭ�ؒ���7��[u����^὿e@޿s������������]����H?��y�ܿrӼ�dN��¶t�^�7�����p��*qV���$�E���
�8]$<`y+<���"����������5�2-q��h���	���'þ��Ͼ&�Ӿ��ξjW����������ok��W0�#U������   �   8�#<�b�<���<�י<�v(��|��8�.��d�о����X��s��x`���ܿƙ ��8����v '���)���&�j��ȕ�� �Rmۿ!+��D����Y�����fҾ���i��I����T��*�<�r�<4�<��;�ڣ��Z�R���\����.�'R�/�m�fw�?}����}�^&k�UN�b7*�W�������G� q���   �   *V=z~;=��(= J�<�nx��ϛ��+��e���$�u�0��=u�c����~˿�f�����#�H�2��<�L@�؈<�H+2���"�z���o��?�˿�)��ޗv�U2�ˆ��v��.�.��z��Xi����<
o=��+=ԋ=�7�<��Q���(:i�i����sܽvQ�N����� ��-ֽ���fGX��:̼@֝:�z�<�   �   �o=Mr= �G=X��<L	���"���@�$:��R\�]�A�|Ʌ�����ðܿ؇�R^�6�1�.C���N�f�R� �N���B��|1�H�����״ݿ����tކ�8�C�����檾�E��	����(p�<<�7=B�a=�~^=R�9=,��<��M<�w�\�ռ<"0��.f����� ��,��q^��3%������pR�Ĭ�<�f=6�K=�   �   P,�=u�=ЯX=@��<@����(Ľ^�N��
���8�A�L��ጿޏ��`���%�jY$�r
;�FN�[�f�_��[��.N��I;���$����� �'��wC����N��'�k&��t�S���̽�ݼ��<�)H=�M�=�U�=�ix=��M=�=L��<&�;�ͻ ����4Lʼ�����q�`�y��n"<�g�<�b&=dX_=�=�   �   `��=7�=}�=HJ)= $��x���u�#>����㾻n(��Fj������ÿxs�pS
����&�+�dx5���8�5��+�&����
�ԑ��XĿ�W�l�\�*�K�羼����#�s�����$A	=8n=Բ�=�ӗ=���=b��=�\= �.=m=L�<Pft<��+<�c<x�B<�g�<|%�<�B=¼J=�O|=2?�=QX�=�   �   �$�=���=��=ƥ(= �T:p�w��{��+���M߾�R%��*f�����翿2��Z�D�ԡ(��I2�Ъ5��G2�@�(�4��o�@���	���:��.gh��X'�a��Pz��k�������ɻ�N	=�j=`��=���=�=o=�A=��= ;�<��H<�O�; �_�����n:p�;H�<���<��*=�a=%�=I��=�   �   r�=��=8}=t&= �b;�8]�z���B��jJҾ�H�+4Z��z��_�����ݿr������< ��2)��J,�T)�:" ��������/޿'l��}Z����[����JYվ($�� ��]u���D���=b]=�=b�|=��]=��+=4��<X<2<pt𗼜j�D��4������#ؼ �j��;B:H��<��=��M=J��=�   �   �[=��r=n�b=8�=P��;�5������h������!�1jG���������I̿�￪� a��`�v�X1���T����+T̿^��_��$�H� H��=���Nm� ���@�I� V�:>�=:rE=�[S=�J:=ԛ=�*_<p������Y�����9���uǽ�̽6�ýᲭ��ǋ�F�B��sǼ�H<��د<ĩ$=�   �    ��<B�,=x�9=(�=��5<lw��)ʽ��E�f0��&;��7d/��yj�mL�����tJտQ��JU��H
���
�p��𿣏Կ(���@%���j���/��q��F�����H��Iѽ� � ��;���<|Q =�=��< ,��@缂ju�\���& �5B�@4�%JB�ԦF���@���0����e����8��JUX�Б�����;�   �   �a��|x�<���<(��<pZg<�I���>������2��P�Ͼz��~G����w���ٷ���Ͽެ⿿���l�7������ο�ζ�������~���F������Ͼ�Ƈ�rW ���o���+<|Y�< ��<�U<p 5�Fu6�<����g��Y7�N�f�����`
��Ht��Ǹ�������7����ĥ`�|~0�B����������   �   P�D�0q=��SD<�'�<((z<��p
P�����R��J��\R�r�"�� R�2g��寘���������ƿ�2ʿDhƿw����竿ƀ���e��r�P�k�!�E�����,:R����F�T�� "�`�O<Ǔ<��<߅���Z�X�н��#�t3f����� A��Oվ���ZD������J ��\V��#ҾWѳ�����_��$�nĽ�   �   ۞н.K� 7M� <��`<���:8��z�������x�����*���4`%�2M��vs�{�������ܟ����)Z��S���)i��wq��K���#�������<v�V7�܃��L�� �~:HuH<���;�-~�XaZ�5�ٽ�2��쁾�`����޾�]������*��4���7�44��c)�z��k�8�ھZ����`}�	�,��   �   \*���½>.����<X�<����5��mȽ�.�u7������*����B���9�?T�\i�5v��hz�!Yu�ʄg�*6R��U7�,�s4�������т��W*�n�½L�-���h <��<x���5�qtȽF.��:������U����E�0�9� CT��i��9v�'mz��]u���g�:R�/Y7��.�N9�������Ԃ��   �   �@v��:�]�����輀+~:HyH<@��;~�VZ�.�ٽ�
2�遾B\��6�޾�Z�J��ӯ*��4���7�\	4��_)�$���h�2�ھ6���Z}��},�o�н��J��M��%<x�`<���:p�輑�������x�:�������c%�x5M��zs�����t���ߟ������\������Gk��:q�K�i�#�������   �   �����=R�����T�+"�(�O<͓<@�<�̅���Z���н��#�\,f�����<���վ~z��=��p������hP꾇Ҿ�̳������^�N�-wĽ$�D�HO=��hD<P,�<`&z<(�TP�����R�eM��2V���"��#R� i������P�� ��d�ƿg5ʿ�jƿ� ��+꫿�����g��@�P���!����   �   '�Ͼ�ȇ��Y ����t��p+<�]�<��<�V<0�4�|g6�X�b�4S7���f�F|�����Zo��ȳ���}��D3��pQ�`� x0��t�������������<���<���< Vg<@Q��}B������4��6�Ͼg���G�����x���۷��ϿG��D��~o�������ο�ж�����t�~��F�����   �   t��ꚥ�,�H�<Lѽ��p��;���<�T =d!=�ʰ< ���|�Zu�z���R  ��;�R�3��BB�z�F�^�@���0�N��U���/��xEX�tx�����;���<6�,=J�9=��=��5<\{�8-ʽ^�E�`2���=��f/��{j��M��l��PLտc��jV��I
�����
�����_�Կ����&���j��/��   �   I�?���Pm�\�����I��?�:
�=�tE=�_S=tP:=>�=xP_<��p����Y���������e�ƽ�̽C�ýi�������{B�hYǼ�y9��<��$=�[=��r=@�b=n�=p��;6!5�Ă��P�h������"��kG��������<K̿Hￌ�b��a�~�X2���&�����eU̿_��2��i�H��   �   ���/Zվ�$��۸��^u� �D�:�=�]=��=�|=��]=��+=��<�_2<����ڗ�pR＠��j����(ؼP�j���D:@��<��=��M=���=�=��=&9}=L&= �b;�;]�����C���KҾ�I�W5Z��{��B�����ݿ�����p= �Z3)��K,�)��" �D��l���0޿�l��[��`�[��   �   �X'���⾉z�����*����ɻ$O	=nj=��=���=L �=.o=t!A=&�=�D�<�I<�~�;�'^��B� �:p1�;��<,��<Љ*=N	a=�=Z��=�%�=i��=��=x�(= �T:z�w�d|�o,���N߾QS%��+f�H��;迿ʩ述���:�(�J2�<�5�H2���(�\4�p����)
���:���gh��   �   4�*��羌���?#�	����A	=x8n=���=ԗ=���=���=�\=j�.=Pm=��<gt<0�+<�d<��B<�g�<�%�<�B=��J=�O|=*?�=FX�=P��=�=�|�=�I)= ���x��v�U>�����n(��Fj�����ÿ�s�~S
����.�+�lx5���8� 5��+�����
�����XĿ�(�l��   �   �W'���⾰y��������`�ɻ�P	=zj=u��=发=� �=�o=�!A=z�=�E�<�I<���;�^��?���:p2�;�<d��<�*=|	a=��=x��=�%�=���=\�=̦(=�U:r�w�F{��+��~M߾�R%��*f����m翿Ԩ� ���~�(�RI2�j�5�NG2�ح(��3��o����S	��:��tfh��   �   ���Wվ&#������Xu��KD��=�]=&�=8�|=��]=~�+=���<@b2< ���,ٗ��Q�F�� ��ʦ��ؼX�j� �D:Ԧ�<
�=��M=ԣ�=z�=Z�=�:}=�&= c;6]�����A���IҾH�V3Z�tz��������ݿ���h��< ��1)�J,��)��! ���R���.޿Bk���Y��P�[��   �   �F��;��CLm�C���B�I� ��:�=pwE=�aS=R:=��= U_<ؠ�����<Y�Q���X���)�ƽ��̽�ýA�����{B��XǼ _9��<��$=�[=��r=��b=�=���;&5��|����h������ ��hG���������H̿O���8`��_�r�V0���p������R̿�\��b����H��   �   �n��0�����H��Dѽ������;L��<:X =�#=�ΰ< (�����Xu�����  ��;�*�3��BB�^�F�D�@���0�8��&����.��EX�,w�����;T��<(�,=@�9=>�=��5<�q�&ʽ4�E��.���8���b/��wj�3K��R���Hտa��8T��G
����R
�N��� �ōԿ�����#����j���/��   �   ��Ͼ�ć�,T ��락�^���8+<4h�<���<�V<��4��e6��쮽�a��R7�W�f�,|�����Fo�������}��63��d6�`�x0�pt���������	����<P��<���<�rg<�;���:�����0����Ͼ��P|G�:��gu���׷���Ͽ���G��kj���6�Ῥ�ο�̶�-�����~�h�F�����   �   ����5R�8���T���!�P�O<�ד<Ȫ<ǅ���Z���н��#�,f������;���վhz��=��a������\P�|Ҿ̳�s����^�&��vĽ��D��F=�0vD<6�<�Cz<����P�F���R��G���N�,�"�R��e��𭘿���D���T�ƿE0ʿ�eƿ����嫿�~��d��b�P���!�X��   �   z6v�3�s}���輀m�:@�H<@!�;P~�PSZ�)�ٽ
2��聾\���޾�Z�=��ȯ*��4���7�W	4��_)�!���h�%�ھ(����Y}��},�Ėн��J��M�p8<��`<���: �輺��'��~�x�A���ͻ��}]%��.M��rs�[���Ƣ��&ڟ��}���W�������f���q�j
K�ԛ#����%���   �   �R*���½V�-� ��HC< <�z�·5��lȽ.�G7��^�������B���9�?T�Ui�5v��hz�Yu�Ǆg�(6R��U7�	,�i4�������т�hW*���½j�-�����:<p<�j�6�5��fȽ�.�b4������8����?� �9�8;T�i��0v�dz��Tu���g�02R�1R7��(�F/��u����΂��   �   ��н@�J���L��I<�`<@��:�����o��6�x�|���
���&`%��1M��vs�x�������ܟ����'Z��S���)i��uq��K���#��������;v��6�����̬� �:X�H<09�;@�}�TIZ���ٽ&2��偾�W���޾�W���&�*�@�4� �7�z4�-\)�����e���ھα���R}�^x,��   �   ��D� !=���D<�<�<�Ez<����P���콋�R�`J��<R�e�"�� R�.g��ᯘ���������ƿ�2ʿChƿx����竿ŀ���e��o�P�h�!�7�认��9R����0�T�x"�(�O<�ۓ<P�<Զ����Z���нG�#�X%f�t���7��,վvt쾦7���������XJ��Ҿ�ǳ�6����^�|��mĽ�   �   ൙�Ę�<���<@��<�rg<0A��|=��4��g2��1�Ͼl�|~G���w���ٷ���Ͽݬ⿿���l�9������ο�ζ�������~���F������Ͼ�Ƈ�W ��<g��P3+<|j�<���<�/V<��4�Y6�T䮽�\��L7���f��w��� ��kj��®���x���.��ꅾ��`�pq0��i��皠�Ľ��   �   ��<��,=��9=��=`�5<0t��(ʽJ�E�F0��;��-d/��yj�iL�����sJտQ��JU��H
�ė��
�p��𿥏Կ)���@%���j���/��q��5�����H��Hѽ�����; ��<�Z =�(=|ܰ< k�����HIu����� �l5�f�3��;B��F��@���0������'%���4X��\��p2�;�   �   l[=��r=&�b=�=0��;H5��~����h������!�)jG���������I̿�￪� a��`�v�Z1���V����,T̿^��`��$�H�H��=���Nm����&�I�@��:�=�xE=�dS=�V:=T�=�w_<Pu�d����X��w������T�ƽ��̽/�ýϟ��.����kB�D=Ǽ�~6���<��$=�   �   H�=��=�<}=�&= c;l7]�:���B��[JҾ�H�'4Z��z��`�����ݿr������< ��2)��J,�V)�<" ��������/޿)l��}Z����[����EYվ$�����[u�`eD���=�]=�=:�|=� ^=�,=@�<��2< N���×�x:�v����~���׼��j� 3G:(��<`�=��M=8��=�   �   �&�=d��=��=V�(= (U:ʯw�{{��+���M߾�R%��*f�����翿2��Z�D�ԡ(��I2�Ҫ5��G2�@�(�4��o�@���	���:��.gh��X'�]��Kz��T�������ɻ.P	=�j=Ӕ�=���=�!�=" o= %A=J�=�N�<�I<P��; �\� ���s:�_�;��<���<,�*=
a=�=���=�   �   ���=�<�=�ϡ=X�l=�.�<�会Ͻ��N���d��~57���t�愛�����c(޿'?���9	����a����L	�Z����޿�B��e��ev��9�#�������UW����t� �P')<��/=H�=f��=���=8ٔ=XT�=��s=�|R=�2=(=Xg=|X�<а�<� =�=,�6=h^]=��=2�=�ɫ=�b�=�   �   d*�=�s�=���=D>l=�N�<ּ[�Ƚ��I�Br�������3��Cp�昿e��C�ڿo(��(��*Z�����Y�d�of��?ۿ���ங���q�՞5�)��2��T!R���۽����N:<�0=��|=��=���=*�=���=@@^=��8=�G=���<h��<p��<��<�ӵ<�=�<��=��>=�)m=���=_n�=���=�   �   �@�=�ݨ=JG�=��i=`!�<x��݅��k�;����8�B'*�d�c�B�� P��c
пpI�p �e���	�W�T` ��F��8п`���T̑��e���+�//�BM���C�`�ǽ����=j<,?1=��s=�Q�=ǅ=@�r=քK=B�=\��< c< �g;�	��`%��M�ϻ �::@�4<X'�<�=6V=�=Um�=�   �   �<�=ٔ=K͍=8�c=@b�<�X��C���%��ۍ�Y�پK���NP��<��B��A�����ؿ���];������ ���1��eؿ^��=��.s��� Q�e��o�۾2Y���+����0Ӵ� }�<�1=�c=��l=��W=�C+=@�<@#<�<�ͼ�#��'S��o�Zv���e���?���$����sg;xi�<��)=0�i=�   �   �A=��n=�x=6�W=�=�]|��m�L�	���r�����"��X7���k�3����\�� ����ҿ��ݿ��῅�ݿ�,ҿ�g��6ߩ��Y��hgk��p7�(���Ͻ���u����v��X25� -�<J{,=��G=��9=�
=Т�<��ϻV@�pl��Ω��8׽Sr��������V��ɽ	����A�|נ�@T�;|��<�   �   X�<
�=�G=C=t�=@j�;�����ԽopD�'��$<����qtH��Mw���W䥿�S��{��[M¿Ǵ��N�������d���#v��G�^��6��Z��N�E�%ڽ.�/� �':`T�<V\ =8=\��< k<���V�T�.���]���&��H���a��"r�w�v��o���]�\�A�ڒ��,��U���G&�Y���   �   \̈́��h[<=�#=��=�6y<�6��C�X���u��������ʗ#�1K��q��G��5Y��d����I��4��`���\m��<Uo�0�I�oY"����}����s��b�vq��������@<�i�<N�	=�/�< ;�;�dм,���G���&�8�]��h�����Đ���:��8�¾W���[��;ޝ��x��)�T�����Ͻ��a��   �   �w�����D<�U�<\�=��<��8�/�Q�ͽl4����8q��!��ĝ�Ж>��Y��ao���|�8���(|�i
n��>X���<����L���'ž�0����0�&ɽ��*�`��Pp�<8X�<�|�< ��;Ǽ� ���P��T	>��7������;�������m�LA������`�ɾg����}���5��u��   �   ��(#c���S� u<���<�i�<�eT<<݃�fgt��b�<�B��ˌ��Ἶ����L%�-6���@�XED�x+@���4���#�[��r�F%��^��̩<�t��*c���S� u<T��<g�<�UT<X냼rt�Ij�N�B��Ό��弾���p���O%��06���@�ID�/@�-�4���#� ��-�,)��!a����<��   �   f�0�,ɽ:�*�@��l�<dY�<��<���;mǼ���:H���>�-4��a騾ԃ;�	�����Vj�1>������꾢�ɾ[���[�}�R�5��m齌w�ؙ��*D<�[�<̞=��<�a�V�/�Y�ͽ�4������t��&������>���Y��eo���|�B���,|�.n�DBX��<�%�������Ⱦ�ׇ���   �   �s�|e�iu��`���P�@<�i�<��	=�8�<Pu�; Pм1y��8��a�&�b�]��d��}��狳��5���¾H���V���ٝ�u����T�/
�$�Ͻ&�a�H���P�[<�=,�#=f�=@,y<�A���������Qu�µ�����?�#� K�`q��I��<[������K���6��Y���)o��qXo��I��["����M����   �    \��6�E�)ڽ&�/� N':PS�<�] =�=��<��<�훼$�T�X��xX���&� H�M�a�r�v�v�5�o�"�]���A�،��"�;M���9&� ��T��<��=G=bC=��= R�;T��9�Խ�sD�m)��<?�� ��vH�hPw�� ��/楿�U�����oO¿ж��9����!���f���&v�\�G�,������   �   �ѽ�'�u����x��P<5��+�<"|,=�G=��9=D�
=h��<�]ϻ3�&`l��ũ��.׽0g�����>��K��ɽ��~�A�p������;��<�A=��n=\�x=�W=�= �|���m�v�	�"�r���������Y7�Ȥk�����[^��������ҿ��ݿz��a�ݿD.ҿ1i���੿+[��sik�*r7�k���   �   ��۾EZ����+�r��x״�l{�<*1=�c=��l= �W=�I+=x��<�3#< �<�̼��#�XS��po��v���e�Z�?����w���"h;|�<(*=�i=�>�=�ڔ=΍=t�c=�_�<�Y�F����%� ݍ�@�پ����PP��=��f�������ؿ9���<��%������	3�Kgؿ;_��@��t��Q�n���   �   60��M���C���ǽ���H;j<v?1=��s=�R�=vȅ=�r=̉K=R�=���<�1c<@Xh;���� ���#��λ =:`�4<�7�<�=0V=q�=;o�=B�=�ި=�G�=��i= �<��Շ���;���l:�6(*���c��B���P��Wп}J뿕p ��e�f�	��W��` ��G��9п����̑�qe�A�+��   �   <)��2���!R�E�۽h��`N:<*0=B�|=��=H��=*�=đ�=NC^=��8= L=���<(��<���<H��<�ݵ<LG�<b�=��>=*-m=��=�o�=���=+�=Xt�=���=>l=HM�<Lּ��Ƚ��I��r��k����3�aDp�s昿�e��͌ڿ)��x��|Z�4��Z����f���ۿ��#���N�q�"�5��   �   ������hUW�O��܋ �))<6�/=��=���=���=Xٔ=wT�=��s=D}R=2=v=�g=�X�<0��<@� =�=B�6=v^]=��=5�=�ɫ=�b�=���=�<�=�ϡ= �l=�-�<\��Ͻ�N�9������57�(�t�����ւ��w(޿;?���9	����a����L	�I���	�޿�B��e���dv��9��   �   �(�2��T R�W�۽���8V:<�0=X�|=��=���=w�=
��=�C^=�8=`L=@��<���<��<���<@޵<�G�<��=��>=X-m=2��=�o�=���=@+�=�t�='��=4?l=�P�<@ּ��ȽH�I��q��!���8�3�JCp��嘿�d���ڿ�'������Y����hY���e��� ۿ5��r���0�q�@�5��   �   �-�%L���	C���ǽL��� Jj<&B1=��s=vS�=%Ʌ=@�r=ЊK=B�=p��<�4c<�ah;උ�P��0"�`�λ�,=:p�4<8�<T�=�V=��=�o�=pB�=bߨ=�H�=�i=�%�<���Y���`�;�S���7�&*���c��A��uO���	п�H뿂o ��d�<�	��V��_ ��E��7п�����ˑ�Ne���+��   �   z�۾�W���+�_��ɴ����< 1=j
c=��l=ީW=`K+=D��<�8#<��X�̼��#��S��oo�Xv�&�e��?�$�w���(h;�|�<�*=ސi=B?�=T۔=3ύ=��c= i�<��X�)A��v�%��ڍ�րپG���MP��;��H�����_�ؿ?���9�����n���0쿆dؿ�\����2r���P����   �   �ͽ�$�u�g��r��5��7�<��,=��G=��9=|�
=H��<PPϻ�1��^l�ũ�(.׽�f������ ���J񽺜ɽ����A�t������;�
�<J�A=��n=�x=��W=@=�|���m�B�	�:�r�������{V7�~�k�����l[��l���/�ҿ��ݿ��ῡ�ݿ�*ҿ�e���ݩ��X��ek��n7�����   �   �W����E��ڽ��/� �):�`�<�b =l
=��<x�<�雼T�T����X�<�&���G��a��r�P�v��o��]�w�A����h"��L��L9&��������<��=�G=�C=ʳ=���;����ԽVmD�%��[9�+��6rH��Jw����⥿�Q��x��JK¿����T�����Lc��� v���G�Z��
���   �   %�s��^��k��`����A<�w�<��	=�@�<@��;(Kм%x��N����&��]��d��]��̋���5����¾9���V���ٝ�u��t�T�
���ϽF�a������[<|	=l�#=��=�Py<x'��h"��ru�5���F����#�pK��q��E��BW��T����G��g2��_���}k���Qo�=�I��V"���Zz���   �   �0��ɽ�*� >�d�<�f�<̌�<P��;XgǼ`��=G��U>��3��9騾��;�	�����Oj�*>������꾗�ɾN���;�}�*�5�Wm�Bw�8���@5D<�c�<ܤ=<��<�����/���ͽ<	4�^����m��������>���Y��]o���|�0���$|��n�<;X�ƶ<��������`���:����   �   7��pc��iS�01u<<�<,v�<�wT<�փ��dt��a���B�tˌ��Ἶ�����|L%��,6���@�RED�u+@���4��#�W��h�8%���]����<����~c�؇S�u<l�<dw�<P�T<�ʃ��[t�[�6�B�mȌ��ݼ�4���]I%��)6�_�@��AD��'@�D�4�J�#�x��t�!���Z��z�<��   �   (�v�\���xND<,k�<�=���<���L�/�5�ͽ�4��q��[!�����Ŗ>�
�Y��ao���|�6���(|�g
n��>X���<����A���ž����B�0��%ɽ��*�@��$z�<�f�<`��<p�;�WǼ���i?��1�=��0��<娾 ;���u��'g�;����8�꾸�ɾ���?�}���5��d��   �   ������[<�=,�#=(�=�Iy<�/������hu�龵�������#�'K��q��G��5Y��c����I��~4��a���[m��<Uo�-�I�kY"�
��s}��˘s�Jb��p��,���(	A<�u�<�	=DH�< ��;x8м�q����㽭�&���]�a��
 ������0����¾-��
R��b՝�q����T�`���Ͻ�a��   �   �<��=�G=xC=ʳ= ��;�����ԽpD��&��<����htH�yMw���W䥿�S��{��]M¿ʴ��N�������d���#v��G�\��.��Z���E�e$ڽ�/���(:D^�<|c =0=T�<��<t՛�2|T�H��S�U�&��G���a�"r�j�v�D�o��|]���A������D���*&�����   �   ��A=B�n=Ԙx=�W=�= .|��m��	���r�i�����X7�|�k�2����\������ҿ��ݿ��ῇ�ݿ�,ҿ�g��7ߩ��Y��igk��p7�%���Ͻ�[�u����u��(5��4�<ڀ,=Z�G=�9=��
=Dƃ<�ϻF%��Ol�b���J$׽�[��&���\���?񽌒ɽ����:qA�ء�� �;��<�   �   �A�=�ܔ=-Ѝ=r�c=Lh�<x�X��B��͕%��ۍ�G�پD���NP��<��A��A�����ؿ���_;������	 ���1��eؿ^��?��-s��� Q�c��h�۾$Y���+����ϴ����<�
1=zc=F�l=��W=�P+= ��<�[#<�� ���̼�#��S�2`o�6�u�2�e���?�����]����h;Џ�<z	*=
�i=�   �   �C�=~�=0I�=v�i=@%�<���f���@�;�����8�='*�b�c�B��!P��c
пrI�p �e���	�W�U` ��F��8пa���Ȗ��e���+�,/�:M��pC�
�ǽ� ��xDj<�A1=��s=+T�=Lʅ=��r=&�K=��=|��<0Sc<��h;�k��������plλ��?:5<DH�<v�=�#V=�=|q�=�   �   �+�=1u�=���=�?l=�P�<�ּ"�Ƚ��I�;r������}�3��Cp�昿e��C�ڿp(��(��,Z�����Y�d�pf��Aۿ���ᮙ���q�՞5�)��2��F!R���۽`��0R:<00=l�|=;�=$��=6�=��=NF^=�8=�O=<��<p��<\��<@��<��<�P�<��=��>=�0m=���=�p�=���=�   �   :��=(�=ꆹ=�=��9=p�;��\�,6�5s�2����g���8�rGm������ʫ�O�¿6տM��{�俺���(տ�ÿ�$��t8��*rn��9�
�����YC}�,-��_��@3��p9�<:@;=Z�u=�\�=�?�=�=.��=vMr=�v^=�?L=`�==��4=��2=�8=��F=�]=�z=��=fZ�=�;�=��=(*�=�   �   ��=t��=���=
��=F<=�c�;>dS�2|���m�[ӹ����[45��i��?���稿y���	�ѿ�ݿ����ݿ�ѿſ��0�������%j��x6�
V�����6aw��	�۳����d�Dθ<��<=��t=Iq�=t�=�<�=�Vx=��a=�J=,-5=b�#=
�=�=TN=�(=�@=�_=�Ӂ=���=< �=�?�=.�=�   �   �=j/�=�+�=08�=��A=H�<x�7��I��]�⚮��t��)h+�E�\�����;��/���@ǿ�,ҿ`�տwҿ�-ǿ'-��y���X7���]��],�����ݱ��Rf�	�x�r�`B�p��<ރ@=X�p=�f�=t9=:�l=�P=P�/=$�=l��<�O�<ȥ�<\f<0bs<HY�<�X�<�==�8=�Ki=`�=��=Ȓ�=�   �   ��=h{�=�R�=H�=��I=P^x<Tq�Wxѽk�D�����侫���I�"y��H��_���%��s4����Ŀ�����*��m+��f y�� J� ���p�󅟾��K���\�?��iT�X��<��D=bh=(�l=��Z=ԁ8=R]=�<`<`QH�ЅY� P���G˼�~˼�D����K� �@��^<�)�<H9=\�v=:��=�   �   OW�=� �=�[�=b�=�fQ= h�<pe��Ѧ�\\%��놾��ƾ�����1���[��\���g��k������=����W���5����K���m[��K1�ԙ�oǾ�T��`'*��e��T}�� �<"�=��F=|BX=f�J=$$=���<P�<��!�R�p�B�&��M隽4V��,ӫ�D¡�����V�V�P���6�H�4<�F=2|N=�   �   ڷ+=��i=�c�=���=��U=�w�<0�޻d�n�B�@\����!�Z��s�:�)^�n�}���_䒿�|��7���즊�t�|�E]�2�9� <�Z$侮����\��Z��V���jc��N�<\h =�C=&}>=��=h�< �<8\ϼHVY� ���"߽!#�v���&�q�)�*R#�@q��[����Ľ_A��,"� �����<�   �   ��T< �=�NQ=��g=�ST=��=�+�;��]�����(�0/���������X���5�z&P���d�}�q�,Lv��oq���c�y�N��f4�����)�s��D~��J�&�@k���6� ar;���<�.=X{7=*=@ĩ< �_���5����`�����B�Z�e������Y��Oڋ�臾j�{��]�`�6��|��½��]��9���   �   ������.<�a=lA=��J=
:'=�ȧ<��F�H/l���*4A�����_�����"S���#��l4��?�D�B��}>�4_3�F9"�����
龃����,����:��/� �\�8�%�0�<�C=ha5=܇!=į�<��4�l�����hu���8�5�r�-����c����;�hѾ�U̾�ؾ��=��s��zg�v�,�
��؃��   �   a��$`��(�\<�$=�58=�3=>8 =���; �ܼ�锽J�.�F�lj���ٮ�S)Ծ�V�����F��,���]�V����*о�Y�������C=����u[���O��8�\<�'=78=@3=n5 = e�; 	ݼZ&	�4�F��m���ݮ��-Ծ�[�����"����x`�����W.оQ]�� ����H=�2#���   �   �5��\��	&�\(�<�A=�a5=��!=0��< �2�zb��)q���8�r�T)��bﭾk^��Θ;�cѾ�P̾ Ծ�k9��ao���sg�A�,���w҃�$�����.<Jf=A=T�J=�8'=���<��F�n8l�Y�8A������!��F�쾤U�X�#��o4�?�|�B��>�.b3� <"�����厷�3/����:��   �   ��&��o��$=��r;8��<��.=�|7=R!=�Ω< /_����L���?Xི���B�y�e������U��Q֋�.䇾�{�]�^�6��w�)����]� $����T<��=�RQ=��g=�ST=�= �;���[���R�(��1���������
�x�5�p)P���d���q��Ov�sq���c�T�N�i4�$��8-�v��s����   �   �\�F]�Z���{c��I�<�g =�C=r>=��=h�< �]8�ϼ�HY�_��c߽����t�&�<�)�L#�wk��P��;�Ľ@9��~��]��d&�<j�+=��i=4e�=G��=`�U=(s�<��޻R�n����\�0��$�D����:��+^�_�}����撿�~��֦��u���D�|��]�U�9��=�('�ה���   �   @V��y)*��h��4�����< �=ؘF=DX=R�J=�$=D�<��< �!��9�4�B�&������M���ɫ�1���뢋�^�V�z��`6�0�4<�O=�N=�Y�=��=�\�=hb�=fQ=�c�<�m��RԦ��^%�d톾%�ƾ&���1���[��]��Ui��ߏ��������qY��e7��T��n���o[�TM1���qǾ�   �   $���L�K�v�佒�?���T�l��<��D=Xh=6�l= �Z=D�8=c=|!�<�4<��G��XY��7��T.˼�d˼P+����K�  >��H^<�;�<̆9=��v=���=��=�|�=]S�=x�=��I=�Ux<u�>{ѽ��D�������t�I��y��I��8`���&���5��ܝĿ��9�+��],�� "y��!J����r��   �   �ݱ�Tf��	���r� H���<ʃ@=��p=Ng�=�;=
�l=ԎP=��/=��=t��<\^�<`��<�|f<h�s<�i�<th�<�D=��8=pQi=��=��=e��=D�=60�=8,�=:8�=�A=`�<z�7��K󽨳]����bv��i+�l�\���������/���Aǿ�-ҿM�տ[ҿ�.ǿ�-��!����7��ۨ]�n^,������   �   �����aw�>
�Q�����d��͸<��<=�t=�q�=��=�=�=�Xx=��a=�J=|05=�#=��=
=�R=�(=�@=�_=-Ձ=��=r�=�@�=��=���=���=���=���=�<=�Y�;0fS��|���m�Թ�b���45�di��?��/訿���ѿ'ݿ���IݿR�ѿwſ�1��:���&j�y6�FV��   �   ����C}��,��_��|2���9�<r@;=��u=�\�=�?�=�=L��=�Mr=w^=@L=��== �4=��2=V�8=�F=&]=�z=��=pZ�=�;�=��=**�=;��=�=؆�=�=�9=@�;��\�l6��s�h���h���8��Gm�ž���ʫ�^�¿@տS��z�俶���(տ}ÿ�$��d8��rn���9��
��   �   �,`w�(	�������d�@Ѹ<�<="�t="r�=k�=�=�=dYx=��a=|�J=�05=��#=Z�=Z=�R=D�(=�@=�_=CՁ=2��=��=�@�=�=���=��=��=y��=<=�j�;JcS��{���m�ӹ����45�Ti�R?��u稿�����ѿ6ݿ��Uݿk�ѿ�Ŀ�C0�������$j�:x6��U��   �   �۱�:Qf�����r�6����<~�@=(�p=Ah�=*==��l=,�P=:�/=��=\��<`�<Ķ�<f<��s<�j�<0i�<PE=��8=�Qi=��=6�=���=��=�0�=�,�=(9�=��A=�<�7��G�ܰ]�����s��wg+�b�\�c����~��M.���?ǿ�+ҿz�տ�ҿ�,ǿS,�������6��ɦ]��\,�:����   �   l���N�K����(�?��ZS����<F�D=nh=��l=f�Z=Z�8=
e=�$�<H;<��G� TY��5���,˼Lc˼ *��șK� �=�PJ^<l<�<N�9=�v=���=�=H}�=LT�=� �=��I=xkx<Fm��uѽ��D�o��y�侤���I��y��G��
^��a$��;3��T�Ŀ����붿�)��c*���y�J�����n��   �   S���$*��a���p����<ؼ=b�F=�GX=v�J=h $=P�<��<��!��5Ｄ�B�v������L���ɫ�ܸ������ރV��y��^6�p�4<.P=��N=_Z�=R�=�]�=�c�=�jQ=�p�<[���ͦ�$Z%�5ꆾ��ƾl���1���[��[���f�������������tV���4�������rk[��I1�X���lǾ�   �   �\�X�pR��HOc�dZ�<�m =�$C=~�>=d�=��< �h8��μ�FY�]���߽n�Z�6�&��)��K#�Tk��P����Ľ�8�����W��((�<��+=V�i=pf�=��=h�U=���< t޻�}n����\����2得��V�:��&^���}�����ⒿN{������Y����|��]���9�,:�3!�7����   �   ��&�xe���-�`�r;(��<
�.=��7=|%=�թ<��^�������W�4��QB� �e�ִ���U��9֋�䇾�{��]�=�6��w�����h�]�@"���U<��=*UQ=�g=$YT=��= `�;Ё����`�(��,��Γ����*�G�5��#P�j�d�7�q��Hv�glq���c���N��c4�����%�p���{���   �   P(�ܔ\�(�%��>�<J=�g5=֎!=8��<�2��_���p��8�M�r�&)��:ﭾK^����;�cѾ�P̾Ծ�]9��Ro���sg��,�Y�҃�ȏ����.<�h=v	A=`�J=�?'=\֧<��F��$l����/A�ᔋ����ϙ쾶P�˦#��i4��	?��B��z>�+\3�x6"�*����އ���)��&�:��   �   �T��<;��h�\<�.=p=8=�3=�< =��;$�ܼ[蔽����F�4j���ٮ�,)Ծ�V����=��$���]�Q�����)о�Y��棃��C=�M���Z���L�� �\<&+=�;8=�3=�> =���;(�ܼM㔽<��F�Jg���ծ��$Ծ�Q��F��n��F���Z������%о�U������f>=�G���   �   �z��/<�m=�A=��J=2?'=�Ч<�F��,l�ü3A�r���0��ѝ�S�}�#��l4��?�@�B��}>�1_3�D9"�����
�u���r,����:�/佲�\���%��5�<�G=hg5=N�!=0��< �0��V��靽�l�"�8�<�r��%��#뭾�Y���;�^Ѿ�K̾xϾ�5���k��/mg���,���.˃��   �   0%U<ޑ=\YQ=~�g=�YT=j�= G�;J��P���b�(� /���������I���5�q&P���d�|�q�,Lv��oq���c�v�N��f4�����)�s��4~���&��j��5� �r;���<�.=��7= (=ߩ<@�^�<������O�L���B���e�4����Q��Hҋ�5���m�{�]��6�Qr�����]�����   �   ��+=V�i=h�=���=��U=�~�<P�޻J�n����\����� �M��k�:�)^�l�}���_䒿�|��7���즊�s�|�D]�0�9�<�O$侢�����\��Z�*V��Xcc�HT�<|l =�$C=L�>=��=*�< D�84�μ:Y�����߽P���B�&��y)��E#��e�F��i�Ľ�0����p���P:�<�   �   ]�=>�=_�=�d�=�jQ=�m�<0a��7Ц�\%��놾��ƾ�����1���[��\���g��k������?����W���5����K���m[��K1�љ�oǾ�T��:'*�*e���z����<\�=.�F=�HX=��J=L$$=@�<(<xt!�0�L�B�����ך��C������믡�����sV�Dk�x,6��5<�X=��N=�   �   ��=�~�= U�=%!�=��I=xfx<�o��wѽ0�D�����侥���I� y��H��_���%��u4����Ŀ�����*��m+��e y�� J� ���p�ꅟ�z�K�ì�^�?� T����<ؼD=�h=^�l= �Z=(�8=j=�1�<�Z< G��)Y����@˼(J˼8���iK��;��r^<0N�<Ў9=N�v=���=�   �   ��=�1�=p-�=f9�=��A=��<z�7�GI�ޱ]�՚���t��&h+�C�\�����;��/���@ǿ�,ҿa�տyҿ�-ǿ)-��x���W7���]��],������ܱ��Rf�	�؎r��>�T��<�@=^�p=�h�=�>=�l=Z�P=D�/=��=���<(m�<<Ń<��f<Фs<z�<4x�<ZL=^�8=fWi=d�=8�=;��=�   �   n��=���=^��=���=(<=�h�;�cS�|��m�Uӹ����[45��i��?���稿z����ѿ�ݿ����ݿ�ѿſ��0�������%j��x6�	V�����0aw��	����� �d��ϸ<��<=$�t=Mr�=��=t>�=�Zx=f�a=��J=�35=��#=��=�=lV=�(=F@=

_=�ց=���=��=�A�=��=�   �    �=0q�=gT�=���=�M�=�=0�T�y͖��t�z���俾�@�9F,���U���}��ʐ�^ڞ�{ݧ�����j৿�枿n萿pV~��fV��+-�i���þ����M,��½"w&���(�T�<=�&B=��R=j�V=��S=hdN=�&I=�E=B�D=�0G=��M=�PX=<�g=R�{=�~�= �=�Ѩ=���=�:�=�J�=Ȋ�=�   �   �=�=l��=޿�=zD�=��=ʌ=h�8�%X��ti��:}�� ��Ƶ��)�8�Q�Yty�:G�����S������]����"��][��V�y�JxR��)���Q������`�'�ko������j��w�<�� =C=fQ=�WS=�.N=F%F=�>=��7=� 4=�4=�|8=H�A=,�P=D�d=t�~=}}�=8�=�q�=���=�.�=���=�   �   2��=���=0��=���=W��=nh=@Sһ����P��x�l�������������F�Wsl�����A(��ژ��;|������D���񆿽�l�;G��c �B����ɳ�0v�&��4����ก;�~�<�(=�LE=��M=jI=��<=�,=Z=,=�=42�<��<8��<,�	=	=�*:=H�\=���=���= ��=���=���=�   �   �_�=��=�E�=T-�=���=��"=�Ԋ:PR������R�s*��ñݾoa��I5��X��w�����v������^��z�����v���W�<;5�	���޾�M��g1Z�����*��dm��;<��=��3=Z�F=~E=^�5=F�=���<\��<$�<�� <ԝ;���:�B�:�=g;�<,ه<PP�<�w=�}T=���=��=�\�=�   �   �G�=܀�=YA�=d8�=��= /5= �'<����Vǽk2�u�������(��G�J'>���Y�t�o��m}����%}��o�^1Y���=����;���!���,艾q�6��׽�H����� -�<"�=l�>=�E=D�5=�= r�<�l< 7�:��2�8b����H��,�$�'���|bԼ8�P� (K;89�<>l=p_=،=�   �   f�{=<"�="%�=��=oq�=RRG=@��<�΢�x����;���`�")���վ���� �ӭ8��uK��lW��j[��W���J��7�
��?�E1Ӿ����j%_�����������;�w�<�3=J�F=�<=ĸ=L&�<��<X��0��ʑF�xi���!���½�н� ѽ%�ĽR����n��|�9�Ԣ��@�;<>�<8}8=�   �   �=@jd=rg�=�|�=c!�=V�U= �< ]�ֵA�ҽ��-��}������pؾ�t�wC���%���/�m3�W/���$���� ��-վ�R���w��|(�!˽��=��Uû��<�C&=��H=�H=c+=�=�<�<��`���$����Y�Ƚ�� ������,�� 8�8�:��3��#�\���<ݽ�O����3� nR���u<�   �   �J&<6!=�U=4{=bh~=،^=�U=��A<�T���������=���������$"ʾ��龮Y�>	�A��F��9 �n���ƾ�̡�ӄy�6�2��b�N�s�,G��Хz<�=H�J=~�W=��B=�= *t<P�;���1������m��l�$�A�L��~p�������P����Ό�nh���}e�|>�" ��~ͽ�q�� ���   �   |��,<��=V�M=V�h= q_="3=���<��!����`���گ�z1:���r�0���o⬾�鿾��˾˂Ͼ�hʾz����������ee��Q+��罆����۹���,<X�=^�M=�h= q_=�}3=���<�)"����代���6:�O�r�|���(款����˾!�Ͼmʾ���5������ke��V+����U����   �   t��U���z<j�=L�J=��W=� C=��=�;t<j;�L�1����e����$���L��xp����b��������ʌ�e���we��v>�^�wͽ�q�h��j&<'=�U=�{=di~=L�^=�S=(�A<�a�����;���=�<���蘦��%ʾ ���[�n@	�������L; ���澜ƾ�ϡ���y�J�2�5i��   �   &˽X�=�p�û���<NA&=�H=B�H=�d+=�D�<��<x�`���$�������ȽY� ����&�,��8�?�:���3�[#�<���3ݽH��P�3��BR�0v<x�=od=i�=�}�=�!�=^�U=���<�Y]��A�"�ҽN�-�g�}�g����sؾ�v��E���%�>�/�3��Y/�%�B��� ��0վ�U���"w�R�(��   �   o�[������0h�;�r�<��3=
�F=��<=�=�-�<��<������F�xb�����w½��Ͻ��н��Ľ�����f���9�Љ����;�O�<&�8=¡{=7$�=s&�=��=sq�=�PG=l��<�آ�#���Y>�t�`�f+��uվd��� ��8�xK�4oW�hm[�W��J�-�7�������3Ӿܶ���(_��   �   ��6�p�׽�H���@(�<��=֏>=ZE=��5=��=z�<()l<@�: �2�<M����.;��+��'��� HԼ8cP�`�K;|L�<�t=:_=�ڌ= J�=\��=PB�=�8�=��=�-5=8�'<j��tZǽ�m2�
������V+����))>���Y���o��o}����]'}��o�X3Y���=�w����������鉾�   �   B3Z�����,��Hs���;<��=ڒ3=l�F=�~E=&�5= =|��<���<��<`� <`�;���:�{�:��g;p�<�<�a�<�=x�T=���=	�=�^�='a�=*��=�F�=�-�=y��=
�"=�~�:�R��
���R��+����ݾ�b�K5�<X�ew�����w������_��b�����v�i�W�t<5�����޾�N���   �   vv����5�������;�|�<x�(=�LE=�M=�I=n�<=��,=�=P=�=,=�<���<���<��	=z=1:=�\=9��=ڒ�=���=C��=��=1��=q��=���=���=��=6g=`dһZ�������l�.�����������F��tl������(�������|��m������$���l�G��d �_����ʳ��   �   V�����'�p������0j��v�<<� =C=�Q=FXS=�/N=�&F=x>=�7=�#4=�!4=�8=��A=r�P=��d=��~=�~�=L9�=�r�=���=x/�=���=>�=���=��=vD�=��=�=(�8�4Y��4j�<}�;��3��^)���Q�uy��G��S������T������I#���[����y��xR���)�P�������   �   ���jM,��½�v&���(�l�<"=�&B=�R=��V=��S=�dN=�&I=v�E=��D=@1G=�M=HQX=��g=��{=�~�="�=�Ѩ=���=�:�=�J�=Њ�="�=6q�=^T�=z��=bM�=��=��T��͖��t�*z���俾�@�VF,���U���}��ʐ�hڞ��ݧ�����g৿�枿e萿\V~��fV��+-�S���þ�   �   ������'�Hn��N����i�z�<�� =tC=�Q=~YS=�0N=�'F=t >=��7=H$4=�"4=��8=�A=֌P=��d=М~=�=j9�=�r�=���=�/�=̡�=0>�=���=R��=�D�=o��=��=�8��W��i��:}�7 ������)���Q��sy��F�����������������"��[����y��wR���)���������   �   rv�׊�2��p�Ṕ;t��<`�(=~OE=|�M=�I=��<=��,=�==2!=�?�<��<���<\�	==�1:=l�\=i��=��=(��=w��=.��=���=Ա�=(��=h��=/��=Nj=pAһA���b��8�l�@�������&����F�\rl�n����'��.����{��	������������l�2G�c �ђ���ȳ��   �   /Z����8(���d���;<:�=�3=�F=h�E=N�5==��<���<T�<�� < %�; ��:���: �g;� <l�<�b�<.�=��T=ϲ�=T�=$_�=�a�=���=PG�=�.�=��=h�"=�B�:�R�����R�:)��/�ݾr`�uH5�:X� w�2����u������]������;�v�`�W��95�ݎ�1�޾L���   �   ��6��׽8H�����6�<Z�=��>=�E=��5=t�=H��<H6l< �:�2�|H����~9���+��'� ���FԼx`P���K;�M�<u=�_=*ی=�J�=��=CC�= :�=��=�25=�(<��VSǽ�h2��������3&�����%>���Y�R�o�Kk}�p���"}��o�H/Y��=�X��|������l找�   �   
�,{������;$��<Ү3=p�F=��<=��=<6�<@�<Ѓ�4���F�:a�����@v½��Ͻ�нz�Ľ,���|f��d�9�t�����;0Q�<�8=ܢ{=�$�=z'�=�=�s�=�VG=ȧ�<����\���9���`��&���վ
�� ���8�[sK�0jW�Oh[�W�Q�J���7���~�U.Ӿ[����!_��   �   *˽��=�@û@��<(I&=X�H=��H=�i+=�M�<��<��`�,�$����G�Ƚ�� �����,�v8���:�e�3�*#���i3ݽ�G����3��?R��v<��=�pd=1j�=V�=�#�=h�U=��<@�\��A��yҽW�-�s�}�ԭ��/mؾ�r�IA�'�%�.�/��3��T/�4�$��	��� �*վ�O���w�8y(��   �   �s�\5����z<�=��J=2�W=.C=^�=�Lt<�Y;���1��ad���$�#�L�9xp�p��:��������ʌ��d��nwe�hv>�5��vͽq��
���n&<�(=�U=�{=�m~=0�^=�[=@B<C����������=���������uʾ���jW��;	����ݧ��6 �.��- ƾpɡ�Ry���2��[��   �   �ƹ���,<F=Z�M=��h=�v_=$�3=H��<��!�(���������0:��r�󟔾>⬾�鿾��˾��Ͼ�hʾk��x������`ee��Q+�Π� ����ٹ� �,<H�=�M=��h=~v_=6�3=���<`I!�0��ԯ��ԫ��,:��r�؜���ެ��忾^�˾j~Ͼ|dʾ\ ������W���_e� M+��������   �    �&<�.=N�U=R{=�n~=
�^=LZ=�B<�M���	�����P�=�X���~����!ʾ��龠Y��=	�:��?��9 �b���ƾ�̡���y��2�vb�h�s��D����z<J�=��J=X�W=�C=Z�=�[t<�B;�t�1��ꣽU]����$���L�<rp�#����������Nǌ�a��qe��p>�O��nͽ�q������   �   n�=�ud=�k�=k��=)$�=��U=��<@�\���A��}ҽP�-�n�}�]���Qpؾ�t�jC�~�%���/�j3�W/���$���� ��-վ�R��|w��|(�� ˽��=��Jû��<�F&=�H=��H=�j+= S�<x< r`�^�$�g���@�Ƚ�� �M��h�,��8�":��z3��y#����-*ݽ�?��"�3�`R�(9v<�   �   V�{=�&�=�(�=��=�s�=VG=h��<�ɢ�Y���F;���`��(��pվ���� �̭8��uK��lW��j[��W���J��7���<�;1Ӿ����O%_���F����㼰��;�|�<B�3= �F=��<=d�=�<�<��<�h����<xF��Z��E��n½�Ͻ�н��Ľ��p^����9�o�� >;�b�<(�8=�   �   �L�=���=BD�=�:�=��=
25=��'<���Vǽ�j2�N��f����(��=�D'>���Y�t�o��m}����%}��o�^1Y���=����6������#艾V�6�ʗ׽�H�P����0�<��=�>=�E=��5=��=,��<�Il<�I�:0�2��5����J-���+���'��r��,Լp0P�@�L;�`�<>}=�_=�݌=�   �   c�=���=�G�= /�=��=��"=�
�:�R�>����R�[*����ݾfa��I5��X��w�����v������^��}�����v���W�:;5����޾|M��R1Z�v���*���k��;<��=.�3=��F=��E=��5=V=���<T��<4�<�� <�a�;��: ¬:��h;&<x��<t�<�=؋T=���=��=a�=�   �   x��=���=���=���=.��=�i=pJһ:�����N�l�������������F�Usl�����B(��ܘ��<|������E���񆿼�l�9G��c �@����ɳ�#v����3�� �о�;��<��(=@OE=��M=�I=�<=��,=" =>=*%=�H�<t��<���<&�	=�=27:=��\=���=8��=��=	��=m��=�   �   �>�=P��=���=E�=y��=t�=X�8��W��^i��:}�� ��ĵ��)�9�Q�Xty�:G�����T������_����"��][��V�y�KxR�}�)���N������X�'�To�������i��x�<T� =BC=�Q=�YS=X1N=x(F=�!>=L�7=&4=�$4=�8=��A=x�P=��d=p�~=J��=�:�=�s�=���=V0�=d��=�   �   �P�=�u�=�6�=:~�=�ޤ=�b=��<�rʼ�֪��� ��>{��H���}����+2���L�Rya���n�g�s�+�n�\~a�=�L�gp2��+�I��K���q�����2��K��<x�Xlռ� \��x&<�4�<�Ţ<�9�<�b�<�[�<���<�Q�<p|�<� =x�%=0�@=@<]=��z=+ތ=�˜=��=�
�=�B�=���=���=��=�   �   .>�=5�=>��=���=0�=Pe=�X�<$���mD��\����u�ץ��O�������.�$�H�e]�0�j�o�=�j�D`]�|�H��/��G���6��+���$H.�'&ٽ.+m��ü �Ӻ@Y><L�<�^�< #�<�!�<�b�<hn�<`�<X��<2�=�-=<?2=�dM=�Cj=�i�=��=��=�µ=���=�3�=�5�=��=�   �   t��=�^�=�G�=���=�>�=6�j=�R�<�����@�����O�e��$��4�ھ��	��K%�N�=�׋Q��^�'`b�� ^�lQ���=��M%�o�	�p�۾�禾�o�<� �qaĽ�L� ���@�a;,g�<\�<�v�<R�<�ͫ<�ş<��<ट<��<`[�<���<�=��=�87=N"U=�[v=1�=���=��=z �=���=`��=�   �   &,�=���=�U�=�o�=�="�r= p�<8�#��ly��t���VM�䓾��ž?����c�5-�0?���J��vN�sdJ���>�/�,�������8ƾ�y��(MT����㣽 �������8<0��<H0�<$\�<�<$��<̲�<xf<`�?<x*<�V'<��8<�`<�s�<HR�<�g�<�=��G=qs=m(�==��=Ⱦ�=�   �   h�=�t�=�^�=���=�)�=�{=��= �	���<�[Cҽ��.��\׫��ھ������b�'���1��05�>�1�f'�x�����o�ؾLʪ���~�J�1���὞�t�����`�;`�<,d�<p�=lp�<�Y�<,l�<�[S<@m�;�],���ϻHE1�HJ`��@n�p;U����L ����;�<&H=�>=�(w=p��=��=�   �   �!�=�`�=�ݴ=G;�=*�=Y�=��$=hI<�����á����z�Q��玾�o��F�ܾ*J���8�������t��k�b��U&ھ@b���싾�M��j
�������P*��8)�<|+=��=$�=�)=j�<�Ƈ<@A�;@�ݻ�ޙ�����y%���F��[��b�b�W�<�;�Z��&���km��eo<��=4�M=g��=�   �   >p=��=x�=��=^�=�р=��6=$��<8�h���b�c�ս�$���b���������E�;S�C�چ�����Υ��\ʾ�9��ތ���W�BS�ýL�I�`�P���l<H=�"0=�n==dr2=�{=��<x7$<dܻ�k̼�3��K��ڣ�����i�׽���z<��ҽ�M��5+��4�L�$�ռ@��D��<4>+=�   �   �D=rV[=��=�ʏ=�x�=�|=ƙB=���< ��Nr	�P���S��q�*�s|^��/��0R��8������a���T˸��H��,U��촁���N����ͽ�je�X;��8�5<�<=*?=��Y=�}Y=ڀ@=��=\��< Cѹ� ¼��J����h2ֽ���<3�4�.��9���:���2�x�"�)�
��۽����`y4���_�pR]<�   �   �(<�	=zL=��r=~=��n=$F=��=�4:<0�u��<��:��"��� ���E�~�f�P6��|���� ����&w���X�G�3�p:
�8��6,_�Dd��X!(<V	=� L=��r=*~=��n=F=H�=�):<H�u��<��?��e���# �B�E���f�59���������2����,w�Y�
�3��>
�	��r7_�Lv���   �   �J���5<48=�?=*�Y= |Y=:�@=b�=P��< vϹ����»J�؀���+ֽ����.�T�.���8�V~:��2�~�"���
���۽����hm4���_�Pr]<K=T[[=��=@̏=�y�=:|=$�B=|��< ���x	�w����
�*��^�u2��.U�����G���尽��θ��K��*X������m O�Ԓ�
�ͽ�te��   �   V�I�X�P��l<z= 0=�l==<q2=�{=��<hA$<�Bܻt_̼��3��F���ӣ�������׽a���3Ὄ�ҽ�E���#����L�|sռ ����<E+=�p=��=�y�=��=��=�р=��6=���<��h�J�b���ս�$���b�Z�������{�;���򾞊�����I���_ʾ�<��k�����W�xV�%ý�   �   ����(���P���!�<�(=r�=��=8)=�j�<�ɇ< X�;�^ݻ�ҙ�<���2p%��F���[�^b��W�̳;�l�������l���o<.�=�M=)��=$�=�b�=ߴ=<�=�*�=�X�=�$=�=<l���Wǡ�����Q��鎾+r��+�ܾmM��O:��������u�Mm��
�� )ھ�d����M�)m
��   �   <��,�t�`���Ə;��<�_�<��=�n�<HY�<�m�<�bS<���; C+� �ϻ�(1��(`��n��U�h��@Q�� ��;���<�P=~�>=>/w=��=��=�i�=*v�=�_�=��=*�=�{= �=�p
�^�<��FҽD�.��I٫�Aھ>�����'���1�c25���1�'��������ؾ̪���~���1��   �   ���1棽���x��(�8<4��<-�<Z�<0�<���<��<�f<��?<�$*<�j'<x9<��`<쁐< a�<@v�<�=>�G= ws= +�=J��=��=h��=h-�=��=SV�=�o�=�=b�r=�l�<h $��py��w���XM�l哾��žE����d��-��?�r�J�gxN��eJ�L�>�g�,���ƫ���9ƾ{��OT��   �   A� �cĽ� M�d ���ba;d�<��<�t�<(Q�<�ͫ<ǟ<H�<訟<@�<b�<���<d�=p�=�=7=4'U=>`v=g�=���=v�=�=��=x��=F��=H_�= H�=��=�>�=��j=P�<t���<B�������e��%��z�ھw�	��L%�D >��Q��^�8ab��^�mQ���=��N%��	�z�۾~覾8�o��   �   �H.��&ٽ�,m���ü@�Ӻ�U><��<�]�<x"�<�!�<�c�< p�<`b�<t��<�=�/=�A2=�gM=fFj='k�=�=��=�õ=���=n4�=t6�=���=�>�=t5�=t��=���=�=�e=�V�< »�|E������u�v�����d�� �.���H��e]�Öj��o�Əj��`]���H�/��G��龘��z����   �   ��2��Kཾ<x��lռ�\�x&<D4�<�Ţ<�9�<�b�< \�<x��<�R�<�}�<2!=�%=��@=�<]=
�z=aތ="̜=��=�
�=�B�=���=���=��=�P�=�u�=�6�=2~�=�ޤ=��b=<��<�sʼ�֪��� �8?{�I���}�'���+2���L�cya���n�k�s�(�n�W~a�1�L�[p2�v+�,��/���\����   �   lG.�%ٽ�)m���ü@\ӺH]><x�<\a�< &�<D%�<g�<4s�<\e�<��<>�=�0=nB2=2hM=�Fj=_k�=��=��=�õ=ɾ�=�4�=�6�=ȱ�=�>�=�5�=���=���=��=
e=(Z�<<����C�����9�u�������羫��H�.���H��d]���j��o���j��_]���H�=/�BG�G�龝�������   �   �� �_Ľ�L����� �a;�k�<��<�{�<�W�<�ԫ<�͟<T�<���<\�<�f�<L��<��=��=�>7=
(U=�`v=��=١�=��=B�=F��=���=���=�_�=|H�=���=�?�=��j=�V�<���	?������e��#��4�ھ�	�@K%�w�=��Q��^�_b���]�kQ���=�M%���	�)�۾�榾F�o��   �   T��7᣽��� ���9<���<7�<�c�<��<��<���<P*f<�?<�2*<�v'<�9<�`<p��<�c�<�x�<�=��G=�ws=i+�=���=�=���=�-�=n��=W�=�p�=B�=��r=\v�<0�#�hy��q���TM��⓾~�žx����b�-��
?���J�{uN�cJ���>��,�r����[6ƾ�x���JT��   �   ���2�t� �����;�'�<<l�<��= z�<�d�<�x�< xS<��; *� �ϻ(1��`��n��U�����&��`��;H��<TQ=2�>=�/w=t��=b�=4j�=�v�=|`�=$��=�+�=*	{=�= s���<��?ҽ��.�
��ի��ھ�����͖'�5�1��.5��~1��'����]���ؾMȪ���~���1��   �   ?����������@3�<(0=h�=2�=�/=,w�<�Շ< ��;@3ݻtș�0���bl%��}F��[�,b��W�`�;�J�����@�l��o<��=΢M=���=�$�=,c�=�ߴ=D=�=v,�= [�=\�$=``<����������&�Q��厾Lm��{�ܾ G���6����ִ�.r��i���d#ھ�_���ꋾJ	M��g
��   �   @�I�0nP� �l<�$=(0=t==�w2=�=��<�Y$<�ܻ�T̼��3�pD���ѣ�7���2�׽K��3���ҽ�D��,#��νL��qռ |庘��<�E+=�p=��=�z�=��=� �=JԀ=>�6=��<Ȳh�n�b��սn$���b�w���؛���;�侓����%��>��~Yʾ�6��zی���W��O�cý�   �   �)����5<�B=�?=��Y=�Y=ʆ@=��=X��< �̹������J�|~���)ֽ���.���.�7�8��}:�1�2�>�"�\�
�O�۽'����l4�X�_��u]<L=�\[=��=o͏=g{�=�|=��B=�
�< H���h	�����w��X�*��w^�-��O��᥯�N|��ͩ���Ǹ�'E��R��&����N����2�ͽ�_e��   �   HB(<.	=�&L=�r=\~=4�n=:F=V�=K:<�zu��<�m8����� ��E���f�6��H���������&w�|�X��3�H:
�����+_��b��@%(<�	=f"L=�r=H~=�n=F=P�=`T:<ku��<�64��|��r ���E���f�K3��S��{�������� w��X�J�3�6
������_�,P���   �   nR=�a[=��=�Ώ=5|�=�|=0�B=��< d���m	�-���`���*��{^��/���Q��������A���:˸�rH��U��ܴ����N�����ͽje��9����5<V>=*?=��Y=v�Y=�@=��=h��< ˹���ЯJ��y��$ֽ:���)��.�D�8��x:��2�S�"���
��۽�����`4�hw_� �]<�   �   
p=� �=|�=��=0!�=jԀ=r�6=��<�h��b���ս$�0�b�����v����;0�*�ǆ�������᾽\ʾ�9���݌���W�#S��
ý��I���P�x�l<� =R%0=.r==�v2=ց=�<�a$<`�ۻ`J̼��3��?��f̣������׽V�⽿*ὐ�ҽ=�����L�L�8Zռ�9�Tͮ<�L+=�   �   �&�=�d�=�=>�=�,�=[�=L�$=pW<p���a¡������Q��玾}o���ܾ
J��~8�������t��k�Z��M&ھ6b���싾�M��j
�_���N��@"���+�<\-=Z�=��=�.=Pw�<؇<���;�ݻL��������c%��sF���[���a�T�W���;����H��� l���o<=��M=Z��=�   �   �k�=x�=Za�=���=�+�=�{=�= 	�@�<�<Bҽx�.���.׫��ھҍ�}��]�'���1��05�?�1�f'�v�����h�ؾDʪ���~�4�1�s���t������;H"�<<h�<@�=x�<�c�<\y�<0}S<0��; >)��dϻX1���_���m���T��� ���,�;�
�<XY=^�>=6w=
��=�=�   �   �.�=T��=�W�=0q�=b�=��r=pt�<��#�ky�t��\VM��㓾��ž*����c�1-�.?���J��vN�tdJ���>�/�,������8ƾ�y��MT�����㣽~����� �8<��<T4�<�a�<t�<ش�<��<�/f<��?<�>*<��'<$9<�	a<���<�p�<ԅ�<$=2�G=�}s=�-�=���=��=:��=�   �   N��=8`�=�H�=Ū�=�?�=��j=�U�<����@��j���e��$��#�ھ��	��K%�L�=�؋Q��^�(`b�� ^�lQ���=��M%�o�	�k�۾�禾�o�0� �PaĽ��L������a;�h�< �<8z�<�V�<ԫ<�͟<l�<���<��<�j�<���<H�=n�=�B7=,U=�dv=��=���=C��=��=k��=���=�   �   ?�=�5�=���=��=��=e=�Y�<����,D��?����u�ͥ��I�������.�"�H�e]�0�j�o�=�j�F`]�|�H��/��G���4��(���H.�&ٽ�*m���ü�uӺ[><��<�`�<T%�<�$�<�f�<Hs�<�e�<��<�=�1=�C2=�iM=�Hj=@l�=���=��=�ĵ=���=,5�=7�=4��=�   �   f��=�z�=�}�=�t�=R��=ZX�=JWB=�O_<<��t^�������]�&���}%¾,���o��5�+� ���#�� �+��|��K�}�þ���`Yj��f(���彁I���#<��l��h����ְ��ȼ��D���\)�H�ݼ�g�� t ���;���<F�=ȓ7=Plj=��=�=�
�=�+�=�=$1�=�D�=`��=�   �   fG�=Z��=X�=�{�=t@�=�{�=�.D=��n<\��Fh���c�&Y�����K���B��.S�ŧ��� �@���>����a��i���<���]�d�O�#���޽UX��$�1�DI�Ў�� a���q���~ܼ8���`����aؼ���X&��gu;d�<8&�<@�-=��_=�8�=� �=�k�=���=�/�=*��=���=���=�   �   ��=�p�=(y�=p^�=#��=v��=I=<�<�v���,��4��<K�є��-�� �پ�t�����������d��������%�پ�泾AӍ�6�T����h�ɽ|��x�����@ll�pta����H8��p�Ӽ��������ɼ�n��H�� �
:��@<��<��=X?>=�ik=7z�=�H�=�ʳ=z��=���=J`�=B6�=�   �   ��=���=�d�=Π�=j^�=�;�=�aO=`J�<����9}��L�6�D�{�����Sž���2����%�	�����&�����%?ľ�q��s�|��};�G��������E��D̼H�5����з���_�@![�X���0w����¼����͚�rV�L�� l?; �H<Ļ�<��=.=T�Y=�ׂ=�E�=H��=�="o�=�L�=�   �   ٠�=���=@V�=��=8��=AR�=��T=x��<�J��9I��>ǽ����RY�P�������kǾ`ݾ#\�������۾t3ž_��W���U�8���wѽ�a}�\d ��R+�@��:���;�9�;�F;�k���#� ��0!���ۯ��
��XG��8�����4��(�� c ; �3<
�<�{ =��/=�`=E��=�<�=�C�=�q�=�   �   ~��=�=O��=��=^�=���=8zV=8��< J��������b���:�3���i��8��5���1����ľ�&Ⱦ�Aþma���Ԣ�������_�L�)�`��J���Ҩ�x�D�Х�;���<���<���<0vc<��;�ͺ`���Ɖ��*�� �޼ �������� ����l�̼�햼�w�@��:Xo<,�<�0= mj=�P�=�6�=�   �   ��=�@�=*�=Ro�=���=�-�=VR=���<���;\¼J�n��ǽ�j�o:� �d��/��pӓ�Hߜ� T���ۚ��ُ��~���U��#)�L���n!����1���b�xr
<�:�<d�=�;=L� =,��<0��<���;0���$V��\��z����?�`�^��|t��1�>N|��j�H��� ���@h9\<� =�mD=8�~=�   �   �a=-�=�F�=؏�=�%�=B�x=N/E=8x =��-<|c��I+��Ӕ�f	ؽ��$�.�tK�3�`���m�Hgp��h��rU�-:����6�{��:L1��R^�@�.<���<L�&=*�>=�@=�/=F�=$G�<��(<п��L���^�H�]�����Fխ�IƽA�ֽ2�ݽ�fٽ1(ɽfŭ�z���;�`ź� t�8�߯<�$=�   �   ��
=J�D=B�h=Njw=�Gq=�bX=��.=��<��E<�1�xU�b�V�SR��O�ν{}������j!�p)���)��!�ֿ�����J����Å����P[��Bo<x�
=R�D=�i=�mw=�Jq=eX=l�.=���<�E< >��[�V�V��'Ͻq���q���n!�Ht)��)�\�!����S�������Ʌ����}� &o<�   �   ��.<��<��&=(�>=��@=�/=ҵ=�C�<�(<��� H���Z���]���dЭ�@Cƽ��ֽ'�ݽ~_ٽ� ɽc��������;����� `�8��<�#$=�a=;/�=vH�=g��=�&�= �x=l0E=bx =��-<0�c�4N+�ה��ؽ� ���.�wK���`�R�m�.lp��h�qwU�:1:�R�������U1��q^��   �   ��b� \
<�0�<"�= 8=� =\��<���<P|�;�����T�����`����?��{^��st�'��B|��j��G�N��D粼�����\\<�� =ltD=��~="�=�B�=��=�p�=���='.�=�R=ؓ�<P��;¼� o��ǽlm��r:���d�$2���Փ��᜾�V��_ޚ�"܏���~���U�')����=&����1��   �   B��H�D���;(��<���<��< ic<���; Vͺ���0ǉ�(����޼����>���� ���４�̼�ږ��Q� ��:X'o<$/�< �0=Bsj=�S�=9�=\��=��=���=��=�=V�=*zV=��< q��������i�����3�1�i��:��r���� ����ľ*)Ⱦ=Dþ�c���֢������_�(�)���,����   �   �g}�Ti �xd+��R�: ��;��;@;�?k���#� ���"���گ�����A��z��8�4�0����� ;��3<��<ނ =V�/=8�`=��=v?�=�E�=�s�=\��=̣�=:W�=Ӷ�=���=fR�=>�T=���<�T��=I��Aǽ���NUY�䗌�����@mǾ^bݾ�^�S�ﾋ��S�۾�5ž4�������U�a��_{ѽ�   �   %�����E�dL̼�5�P���`Л�Pk��+[�����Pz��@�¼����˚�`jV�05�� �?;��H<�Ŵ<*�=�.=�Z=Hڂ=FH�=T��=��=�p�=(N�= ��=f��=Te�=I��=�^�=�;�=\aO=�G�<|���=}�zO�d6���{���]Už���.���	�2�	�����(��k�㾮@ľ�r����|�t;�����   �   )�ɽ.|��{�����`vl�~a�`��P<����Ӽx��h����ɼhm���� n:A<���<�=�B>=mk=�{�=6J�=m̳=��=��=Xa�=,7�=؛�=rq�=�y�=�^�=B��=j��=~I=��<�z��h.��5��=K�����!.��V�پv��������}��#��\�� ��<�پ糾ԍ�{�T�����   �   ��޽0Y��� 2��L�����0d���t��0�ܼ0����X���`ؼ����"� }u;��<�)�<8�-=��_=�9�=�!�=�l�=���=�0�=���=D��=B��=�G�=���=��=|�=~@�=�{�=@.D=x�n< ��9i��Hd� Y�����L���羦���S�1��;� ����Z?�F��������������d���#��   �   ��彟I��$<��m��p����װ���ȼ��X���)�P�ݼ�f���p � ��;T��<�=��7=�lj=�=T�=&�=�+�=:�=N1�=�D�=x��=~��=�z�=�}�=u�=M��=DX�=WB=8N_<H���^��&���]�F����%¾M���o��5�2� ���#�� �+��|��K�n�þ���OYj��f(��   �   ��޽�W���1��G� ���P_���o�� |ܼ����d �8���[ؼ0��P�@�u;�!�<\,�<:�-=��_=�9�=�!�=�l�=���=�0�= ��=h��=b��=�G�=ހ�=��=\|�=�@�=|�=�/D=��n<�Ἓg��8c��Y�����K��������R�j��o� �ݘ��>�������ֿ��������d���#��   �   ��ɽ0|�pv�8���cl�pka��	��x2���|Ӽh�缈�弐�ɼ�d��`���E:�A<l��<�=jD>=Vnk=v|�=�J�=�̳=*��=T��=�a�=l7�=��=�q�=z�=@_�=���=b��=I=�!�<dq��G+��3�b;K����/,���پ�s��A�����������������پ�峾^ҍ�åT�����   �   "�����E��=̼0�5�Pn�������P�@[�����hl����¼�������� UV����@�?;��H<�ʴ<>�=��.=�Z=�ڂ=�H�=���=@�=q�=�N�=���=���=�e�= ��=�_�=�<�=�dO=lQ�<X���4}��I��6��{�l��<RžI��Q�����	�����$����㾂=ľp��
�|��{;�����   �   �[}�,_ ��@+��V�:��;�\�;��;��j���#��m�H���˯�`����4��o����4�Pٟ�� !;��3<��<l� =��/=0�`=���=�?�=,F�=t�=ɢ�=X��=�W�=���=׻�=	T�=��T=���<5�83I��:ǽ���PY�����ƥ��iǾ�]ݾ�Y�c�ﾲ�꾹�۾J1žo�����8�U���tѽ�   �   ���XmD�p��;8��<T	�<�<(�c<`8�;�4̺ت�����`��h�޼���P���� �<����̼�Ֆ�I��,�:�,o<l1�<�0=&tj=�S�=�9�=���=@ �=V��=��=b�="�= V=<��< �V��.�������3�N�i��6��땦�����g�ľ�#Ⱦ?þ�^��LҢ�������_�>�)�O�� ����   �   8�b���
<`E�<v�=�@=ĉ =8��<ȗ�<�ŵ;�K���B����⼤�� �?��u^��nt��"��?|�<j���G�����䲼 ���h`\<�� =NuD=��~=�"�=(C�=��=�q�=��=0�=�R=p��<���;������n�&ǽ�g��k:���d��-���Г��ܜ�qQ��'ٚ�)׏�g�~���U� )����I��b�1��   �   @�.<���<µ&=X�>=DA=��/=|�=XU�<0�(<v��\7�� S�L�]��񏽛ͭ��@ƽ��ֽ��ݽB^ٽ�ɽ����O����;�Ȯ�� �8��<�$$=�a=�/�=BI�=^��="(�=½x=N5E=�~ =X�-<(Yc��?+�Δ��ؽ��.��
K�Y�`���m�+bp��h�nU��(:����C轋��@B1��1^��   �   $�
=�D=�i=�rw=Pq=�jX=��.=8��<ЯE<���DF�H�V�O��m�ν{�����i!�jo)��)���!����0���ڸ��oÅ���0X��Eo<t�
=r�D=�i=�ow=`Mq=thX=��.=(��<�E< ��A�(�V�L��D�ν�u�����@f!�|k)���)���!�����������}������P6��ao<�   �   �a=�1�=�J�=Ɠ�=>)�=x�x=r6E=P =�-<x`c�NC+��Д��ؽ~��.��K���`��m��fp�]h��rU��,:�\����!���K1� P^���.<���<��&=��>=@�@=�/=D�= R�<P�(<Pv���4��XP���]��fɭ��;ƽ��ֽ�ݽaWٽ�ɽ۶����0;�L��� ��8\��<�*$=�   �   �$�=�D�=��=�r�=䛝=�0�=j	R=��<@��;� ¼��n�Fǽ�i��n:�L�d��/��,ӓ�ߜ��S���ۚ��ُ��~���U��#)����&!��J�1���b��u
<�<�<��=�==Ԇ = ��<`��<���;�R���B���⼾��r�?��o^��ft���25|�Pj���G�����ϲ��J��`�\<ڏ =�{D=��~=�   �   ���=�!�=x��=��=�=��=0V=��< ��F��}���j���X�3�)�i�R8����������ľj&Ⱦ�Aþ]a���Ԣ������_�0�)�$��	���>����D� ��;䨆<��<��<(�c<�$�; w̺ �� ������p�޼4�����8� ����p�̼�Ė��&��=�: Mo<p@�<��0=zj=tV�=�;�=�   �   ��=j��=�X�=b��=K��=DT�=��T=��< <�,6I�=ǽB��RY����k����jǾ�_ݾ\�������۾l3žW��N����U� ���wѽHa}��c ��O+����:P�;�F�;�i; �j�p�#�Pu�����̯������1���i��Ț4������X!;��3<8)�<�� =��/=ڿ`=��=B�=H�=�u�=�   �   n��=���=�f�=r��=�_�= =�=�dO=�O�<`��d7}��K�%6�֔{�����Sž��� ���� �	�����&�����!?ľq��f�|��};�4������Z�E��C̼ؕ5���������xY��[�ଗ�p����¼����(���SV�P���@;`�H<�Ѵ<@�=��.=$
Z=�܂=�J�=���=��=hr�=�O�=�   �   ���=Br�=Zz�=�_�="��=q��=�I=� �<xs��%,���3�M<K������,���پ�t�����������d��������!�پ�泾<Ӎ�,�T����I�ɽ�|��x�����8jl��qa�����5���Ӽx��(�张�ɼf�� ���_:0A<l��<ک=�F>=�pk=�}�=�K�=�ͳ=B��=L��=lb�=8�=�   �   ,H�=��=��=v|�=�@�=|�=�/D=p�n<����g��vc�Y�쉔�tK��
�@��-S�ħ��� �?���>����a��h���:���U�d�G�#���޽CX����1��H�8���``��q���}ܼ����4�����]ؼ���x���u;�!�<�,�<��-=H�_=Y:�=\"�=qm�=H��=D1�=b��=���=���=�   �   �=>�=j��=\�=-I�= �=l;�=B�*= �4<�3ռ[V���h�b�0�3j�,됾�䩾����yʾ�ξ�Tʾ����������%p�� =��	�Z�ҽMʛ�T�t���[�vmf�^k���!��x��w�۽�_��$����� ٽ�b���̎�ܹ?�@仼 �9��<��-=��u=!p�=�\�=B��=�<�=Xm�=��=�t�=�   �   ���=�1�=��=��=G�=�"�=tÇ=bT+=�d=<�0̼�������
-��He�m���Rx��3繾�aƾ��ʾ}-ƾ���by���ڎ��j�,48���
�N�˽������i���P��[� ���������4�ԽL�罜��;�!
ԽNh��Z��8�<�0k�� @���<0(=�eo=�ݖ=x��=�N�=v��=�F�=ȭ�=���=�   �   E�=K�=���=���=��=�$�=�"�=��+=PzT<�������J޽$g"��zW�������߮�z���au���&���*��u꛾Jo��Q$Z�lD*�ci��\ɷ��1���I�\2��8<��~`��y���R��}h���Խ��۽�׽9�Žg:��������5��Q��@����<��=T[=&ދ=r�=$P�=�o�=Z��=��=^b�=�   �   D��=��= ��=8��=r�=Œ�=���=�*=�q<�k����`�o�ƽ0"�T_B�� q�rh���ܝ�yM������z|��X��F|���m��@����ٽ#Y���KQ��O�`f��r�,��(^�tf��̏���O�����q��!)������u��.��"ż����p�J<�<�*7=�Zq=g�=p�=���=>��=���=�x�=�   �   �,�=�=f�=��=|A�=X��=<�x=��%=��< U�΢=����������(��Q��u�����`s���������ᅾ�vm�ddH�dF ���� ���M`�h�
��U���I��hR��H�ּ��^nL�}��ɑ�9�������^��&e���a��n+� �߼(�I��+.;���<:� =f08=4�l=��=�	�=�/�=x��=���=�   �   z*�=�:�=���=n�=�"�=~�=��c=n=P�<������o� �ӽ���dV.��K�"�b��Mp���s�ܹk�6�Y�Z�>�8�������󲽞9j��r��wg�`\J���}:@斺P���~������<,�t�T�Ȅq� ���~�Tp�~�V���4�|��x�����D� x�8�oP<hf�<��=��S=ݳ�=��=��=~2�=�   �   ?��=�K�=�=w�=�*�=|�|=E=�=��Q<xM�Tr�|Nm������w佪'���"��t3��=�>�46�J�%�n��=���m��X�b��Q�H-� �;(��<`/�<�h�< -< 6\:��-�����5���,�PhG�TjW�Hu]�Z�Z�(�O��4>�8�%��.��J����H� ?�9��g<�
�<�W.=Td=Z2�=zn�=�   �   k��=ރ�=�0�=�2�=~:v=��M=�[=�ؼ<���;�|4�Ĺ����J�bC��t��d�ڽ�:���{�����A�6�>���#���x��T�A� "¼�{��av<?�<|J=<�=��=Ԏ�<xC�<�<�����Q�:#�^�?� �\�4\s�R��K����,��Z�w���\�\t4�h� ��~��  ���<��=�9?=H�m=�   �   �NC=<�Z=�s`=��T=�B:=�U=\p�<(�3<@�J��׎�����;���q�?�����D�� ½��ýꂻ����ؕ���-X��b	��5\����;X?�<@�=�SC=>�Z=Bx`=*�T=<G:=
Z=�x�<��3<�dJ��ӎ�.���;�v�q���𢧽�H���$½�ý����ͣ��m���n8X�hl	�0X\����;�1�<T�=�   �   �3�<E=�=��=���<|9�<h�<0?�������W�%���?���\�Ys��O������(����w�}\��j4�Ҍ �Xl�� @�6,'�<��=�??=��m=���=��=�2�=�4�=L>v=<�M=,_=@޼<P�;8y4���� �J�hE��z��\�ڽe?���~�����D�n
�v���)��~����A��2¼���XHv<�   �   ���;��<�$�<^�<` -< �Z:`.�x����:���,�.kG��kW�6u]���Z���O��/>�&�%��'��;���uH� 6�9بg<��<8^.=,d=�4�=�p�=P��=�M�=��=�x�=,�=R�|=�E=�=P�Q<PN��s��Qm�4��� {��)�z�"��w3�D
=��>��76�� &����ű潪r���b��`�hG��   �   ��g� �J��h|:����`���������<B,���T�6�q�����~�8p��V���4���d����|D� 8 9(�P<$s�<�=p�S=|��=: �=��=f4�=1,�= <�=���=��=�#�=�=l�c=h=�<�����t��ӽ����X.���K�S�b��Pp��s�V�k���Y�l�>����q��������@j�Dy��   �   ƺ
�`���S���\����ּ<��sL�r"}�C̑�s������`���e��(�a��m+�x�߼0�I� m.;���<� =^58=�l=8�=��=�1�=*��=(��=J.�=B�=��=��=ZB�=��=:�x=`�%=,��<8U���=�5���������(�%Q�eu���� u��L��H��dㅾ�ym��fH��H �Ϋ�s����R`��   �   fPQ��S��j����,�R-^��h��1���;R�������r��P*��w���u�:.�Pż�봻`�J<��<X.7=�^q=6�=�q�=��=���=ʙ�=�y�=L��=��=З�=���=�=<��=٪�=��*=�q<�n��� a�n�ƽ�#�aB��"q��i���ݝ��N��h����}��eY��{}��6�m�Ң@�|���ٽ�[���   �   a3��b�I��
2�f<<�R�`�u{���T��Tj��fԽD�۽�׽�Ž�:��������5��N�����P�<�=�[=pߋ=Zs�=[Q�=�p�=^��=p �=(c�=�E�=�K�=J��=��=�=%�=�"�=^�+=(wT<������kL޽:h"��{W�����k����ா����lv���'���+��R뛾p���%Z��E*�jk��2˷��   �   �����i�� Q�N�[�4���������L�ԽB��a����e
ԽVh����L�<��h�� ���@�<�(=�go=Zޖ=B��=�O�=��=�G�=L��=\��=0��=J2�=�=P��=r�=�"�=rÇ=T+=�b=<3̼|������-��Ie������x���繾Obƾ�ʾ
.ƾ�����y��`ێ�΁j��48�~�
�Z�˽�   �   �ʛ��t�Ơ[�hnf��k��["���x����۽�_��$��`�e ٽqb��e̎���?��Ỽ�
 :��<��-=��u=�p�=�\�=���==�=�m�=��=�t�=B�=\�=���=j�=0I�=��=S;�=��*=��4<�4ռ�V��i��0�jj�H됾�䩾����yʾ�ξ�Tʾ����������%p�� =��	���ҽ�   �   %���.�i���P�n�[�����N�����_�ԽD��\���轂Խ�f�������<�Pd�� @l�D�<(=�ho=�ޖ=���=�O�=H��=�G�=l��=|��=P��=r2�=.�=���=��=W#�=�Ç=rU+=�i=<`.̼�������-�He�����w���湾?aƾ�ʾ�,ƾ�����x���ڎ�[�j��38�s�
���˽�   �   a0��ԻI�N2��6<�p|`�Dx��,Q���f���Խi�۽�׽k�Ž7��������5�HF�� K� !�<^�=�[=!��=�s�=�Q�=.q�=���=� �=hc�=F�=�K�=���=���=��=�%�=�#�= �+=ȄT<��������H޽f"�1yW�/��������ޮ����\t��%���)���雾{n���"Z�<C*�ig���Ƿ��   �   �GQ�L�c���
���,�r$^�d������L��C|��om��Q%�������t�.�Xż�Ĵ�8�J<$�<�07=v`q=��=Mr�=���=��= ��=6z�=���=$�=R��=���=��=B��=<��=��*=.q<xb����`�o�ƽ| �^]B�]q�;g��V۝�L������{���V��{��Ԅm���@�4~�N�ٽ�V���   �   ��
�M��,A���I����ּ� �nhL�P}��ő���K���/Z��Z`��n�a�"e+�@�߼�I���.;��<�� =�78=��l=��=k�=,2�=���=���=�.�=��= �=���=JC�=P��=��x=Ĳ%=���< �T���=�5���o����(�Q��u������q��������=����sm��aH�D ������^G`��   �   �ag� J���~: G�����r������5,���T�t{q�0u�.~~�lp�d~V���4�l��؞���hD� >9ؕP<�w�<��=�S=��=� �=r�=�4�=�,�=�<�=���=��=�$�=u��=�c=L=0�<�������쎽�ӽ
��LS.���K���b��Ip�׆s�.�k���Y�$�>�V���}��(ﲽ(2j��l��   �   �2�;亃<�9�<�s�<--< �]:��-��x���,� �,��]G� _W�di]�"�Z���O�,(>�ڕ%��"��3��HiH� o�9��g<��<|_.=@d=m5�=Eq�=Ҳ�=cN�=��=�y�=$-�=.�|=LE=�=h�Q<�,�Di�zDm�"{���q�h$�>�"�#q3�"=�P>�X06���%�-��c�潗h��b�b�XB����   �   �J�<�O=��=^=���<�P�<@�<@َ��܇�@=�H���?���\�$Os�^K��n����%����w�Fy\��g4��� ��h�� ��6�)�<ƾ=�@?=��m=Q��=���=�3�=x5�=l@v=�M=�b= �< 9�;hX4�@���V�J��=��M��͟ڽ�3��Fx�����=���x�轹��(s��T�A��¼ ��{v<�   �   �YC=n�Z=l}`=~�T=�L:=^`=��<��3< �I�����<���;���q��鑽ڛ��hA��p½��ý;���Ü��ڔ��Z,X��a	��1\�P�;A�<�=�TC=B�Z=�y`=��T=4I:=�\=��<��3< J��Ď�����;�L�q�4葽[���>��K½ߍý|��w�������b"X�\X	��\��:�;�M�<z�=�   �   c��=���=C5�=!7�=�Cv=&�M=�e=\�<�J�;�R4�����|�J�?������ڽ�7���z�Ħ��@���f��P#��Bx��j�A�T ¼�n� ev<�@�<dK=X�=B�=X��<H�<��<����䇼(D����?���\��Ms��I�������"��,�w��p\��^4�Ɓ ��W�� �Y7�7�<�=�E?=F�m=�   �   ���=P�=��=�z�=t.�=��|=�E=�=��Q<�*��i��Fm�}��ht�T&���"��s3�5=��>��36���%�,��ӫ�cm����b�PP�*��	�;ı�<D1�<$k�<�-<��\:��-�H���x1�F�,�HaG��aW��j]��Z�&�O�%>�b�%�,��&���MH� ��9��g<�(�<be.=zd=�7�=Fs�=�   �   .�=�=�=���=��=&�=j��=��c=�=h�<؟����VT�ӽ���XU.�>�K�v�b�Mp�*�s���k���Y�,�>���L���8�9j�Rr�0ug�`RJ� �}: ɖ�����{������9,���T�@�q�fy���~��p��V�T�4����d����YD� �9��P<p��<4�=�S=m��=�"�=J�=�6�=�   �   �/�=��=�=���=D�=���=��x=t�%=ܘ�< �T�ĝ=�����������(�Q�u�X���2s���������ᅾ�vm�NdH�HF ����撪��L`��
��T��HH���P��p�ּ���lL��}�]ȑ�u������\���a��n�a�f+���߼x�I�`�.;��<r� =X;8=��l=��=*�=�3�=���=���=�   �   l��=��=��=��=\�=���=���=��*=�-q<d��H�`���ƽw!��^B� q�>h���ܝ�ZM��桫�j|��
X��;|�� �m��@����ٽ�X���KQ�0O��e�� ���,��'^��e��	���O��[~��to��/'��m����t��.��ż�´�@�J<l�<�27=�bq=,�=�s�=���=*��=��={�=�   �   |F�=VL�=���=���=��=&�=�#�=0�+=p�T<����k���I޽�f"�!zW�ƈ��c����߮�k���Tu��x&���*��n꛾Fo��E$Z�bD*�Mi��Gɷ��1��ҽI�2��8<�8~`�Ny��[R��h��Խ��۽�׽��Ž�8��砄���5�hH��@X�H!�<��=�[=���=�t�=sR�=�q�=L��=F!�=�c�=�   �   t��=�2�=R�=���=��=|#�=ć=�U+=�i=<�.̼)���'���-��He�Z���Dx��(繾�aƾ��ʾz-ƾ���]y���ڎ��j�)48���
�B�˽������i�p�P�Ԡ[�ཀ����U����Խ ��6��|	Խ�g��v��0�<��f�� `z�(�<�(=�ho=�ޖ=���=�O�=���=�G�=���=���=�   �   ~�=�"�= ��=��=�G�=n��=t�=Z�v=r<=(P<@���·K�E7�������/ �&@��gY���i�R�n�z&i�Z0Y�jIA��$����~�ֽy��^u������������޴�2�t�/�8wN��(h��2y�.��y�hbg���K��C)�e���k���P��م�P�k<ZP'=�#�=�p�=�?�=^?�=��=�`�=���=�   �   &�=��=�e�=~��=�=�c�=Nu�=�[s=p=��M<����G��Ϊ�M������%<��T�Rud�t�i�Y�c�*	T��|<��> ������Ͻ�ʤ�`����e���5��-9����۽v��*��bI�d�b�>�s��zy��s��eb�`�G���%�E������&aL��M��(;j<�E%=�=�u�=T�=���=l��=^5�=�{�=�   �   8��=@��=���=��=I�=S��=C�=i=4�=��C<�z��<�FE����a���0�DvG�:�U��>Z�E_T�F E��.�L���ｍ���Ԣ��trq�>�a�`"x�B���W�ƽA�������:���R��c��i���c�FT��);�Л��e�:���a@�hqs��Db<{=v�t=wP�=�\�=m�=��=p��=��=�   �   `��=i�=�X�=BK�=�/�=Z�=�A�=PV=�=0�(<�Du�~�.�]���Z�н���.�,3��\?���B���<��.���������˽u��DFl��H<�$�-��SB�P�x������ٽ���d�#�vY:���I���O�a�K�-;>��Z(��h���ٽA9��Ns0�X>d��"J<��=D<b=`c�=ʩ�={=�=h]�=V6�=���=�   �   ���=�I�='��=9�==�d�=v�x=�8=�n�<pa�; I���"�����6���6��D
��,�֜#�|?%�L����0��
�ͽkŞ��g��O#�@3��ռ4����J.���x��ڪ�Cݽ�����*���0�7.���#�`��b�������-��j7"���i�H�<���<�D=���=�6�="ƴ="M�=���=���=�   �   }�=���=Dƹ=P�=���=zF�=ޢI=�'=�y�< ��`���j-�f=r��᡽c�ǽ�������n��������:��!���O��ΕW�����ϟ�8�'��O�X:�X������Bl�[k��Źͽ�"��1��:�
���Vm��ϽN����
u�T>�@׌���%;�*�<r6=D{V=|8�=��=�i�=Ӡ�=Pb�=�   �   u%�=o7�=��=F�=
s=<�A=�a
=䰞<0�;�o2�tS׼�J*��Eg��L������载m˽>Ͻ`]ɽR(�������J~�8�5��$ڼ �-���;p7$<�VL<|< ��8`��w��vK�q����㭽�Ƚ�ؽ-�ܽ��ֽ��ƽpo��$����f�2�$��xļ8�����;�Ժ<N=�N= �}=<t�=R��=L��=�   �   �֌=�i�=4�y=�6V=�S(=�3�<HKg< ̛���b�-ۼ4���9I��o�Ie��Ҡ���X��P��]�� \����t�j�A� &��p��@���5P<`��<F�<��=�]�<4��<�&%<`5��Z����މX��$��tʘ�Qa������{������
���k��@�����:��p$�@x;Ñ<j� =d�3=��^=��=��=�   �   �lR=.8H=&�-=�t=ܣ�<�ͩ;�� ���Ƽ���D��g���ݫ���h��}���ł�j�r�XW���2���b��6��x�<Tƹ<&=��3=@bK=FrR=�=H=��-={=$��<��;�� ���Ƽ:z��D��g�"�檆��h��T��eǂ�.�r�^W���2�$��pp���n����<���<4�=�3=�\K=�   �   2�=�Q�<���<�%<�p���i����.�X��(��(Θ�}d�����J}��{���
���k���@�T���/����#� �x;Lϑ<L� =�3=��^=��=�=;ٌ=l�=R�y=H<V=�Y(=�?�<0cg<  ��H�b��#ۼ����7I�Ro��e��P���8[��Q�������_��ڹt���A��-����@l���P<d��<�:�<�   �    ?L<c< �|80"`������~K�����|譽Ƚ�ؽڽܽ��ֽ��ƽ�p������J�f���$��qļ��@ �;�޺<`=�N=ұ}=�v�=���=^��=�'�=�9�=��=OH�=�s=�A=Lf
=ܹ�<@(�;c2�$O׼�I*��Fg�N�������꽽�
˽BϽ�aɽ�,�����>S~���5�(3ڼx	.� ;�$<�   �   �(:�������Xl��o��g�ͽd'�L4��<������o�.�Ͻ����
u�=��Ҍ� )&;2�<�:=lV=�:�=��=mk�=���=d�=�~�=r��=ȹ=�Q�=���=XH�=��I=+=��< �������-�F?r�3㡽؜ǽ��������p� �a������H���S��ڜW����۟���'��   �   ��ռ����(Q.���x��ު�JGݽF��8��/*�0��8.�F�#�����������o���6"��i�ؙ<T��<4�D=+��=i8�=�Ǵ=�N�=���=R��= ��="K�=���=v:�=`��=f�=�x=�!8=8r�<pi�;�H��>�"������������
�j.�؞#��A%�j����4����ͽ�Ȟ��g�jU#� >��   �   �-��XB���x�����ٽq��Z�#�t[:��I���O���K��<>��[(�Ai�Q�ٽ~9���r0�@9d��)J<2=�>b=�d�=	��=�>�=�^�=t7�=���=j��=j�=�Y�=HL�=�0�=R�=�B�=�V=�=��(<�Fu���.�����)�нL��A0��3��^?�U�B�ϐ<�B.����������˽ ��Kl�|M<��   �   �a�x&x�����٪ƽ������r�:�T�R�bc��i���c�0T��*;�>���e�:���`@��ls��Jb<�|=^�t=kQ�=z]�=H�=��=:��=��=��=���=r��=L�=��=���=�C�=�i=��=��C<�}���<�bF�����P���0��wG���U��?Z��`T��!E�M�.�j����s�������vq��   �   g��	7���:��c�۽b��*�|cI�Q�b��s��{y�|�s�!fb���G���%�������� `L�K���@j<�F%==Tv�=��=���=���=�5�="|�=��=6�=:f�=���=p�=;d�=�u�=�[s=�=x�M<L���6�G��Ϫ�C��h��F&<���T�vd�5�i��c��	T�P}<��? �`����Ͻ	̤������   �   ?��9��y������z2�Ճ/��wN��(h�3y�.��y� bg���K�EC)�����j��X�P��օ���k<�Q'=$�=<q�=X@�=�?�=��=�`�=ԕ�=��=#�=D��=��=�G�=t��=�s�=,�v=2<=�P<@���d�K��7�������/ �/&@�hY���i�m�n��&i�j0Y�tIA��$������ֽ����u���   �   �e��5��9����۽P���*�$bI�ٯb���s��yy��s��db�4�G�U�%���������:]L��F���Gj<LH%==�v�=B�=���=&��=6�=>|�=��=b�=bf�=��=��=�d�=�u�=�\s=�=�M<(�����G�Ϊ�d��R��
%<�y�T��td�Și���c��T�|<�^> �\����Ͻjʤ�����   �   T�a�� x�G���>�ƽ������ߧ:���R�uc��i���c�eT��';����b��6���[@��[s��Wb<H=H�t=&R�=^�=��=�=���=��=2��=8��=ʾ�=��=e�=���=\D�=�i==X�C<�m���<�\C�����:����0��tG���U�E=Z��]T��E��.�@�����������Bpq��   �   �-��PB���x����w�ٽ?����#��W:�ڳI���O���K��8>�X(�f��ٽ�4���k0��!d�<J<�=dAb=�e�=ҫ�=D?�=_�=�7�=���=ȗ�=�j�=6Z�=�L�=G1�=�=�C�=jV=>= �(<x0u��.�i���,�нj��-�F3��Z?���B��<��.�g������O�˽+��TBl�TE<��   �   ��ռ����PF.���x��ת��?ݽ�����f*��0�.4.��}#�j������-�����."�P�i���<���<l�D=a��=V9�=fȴ=:O�=v��=���=p��=�K�=��=;�=��=g�=��x=%8=�z�<@��;�;���"�����!���ݓ� 
�7*�p�#�=%����k�,��g�ͽ8�<�g��J#�l*��   �    )���9�ț��ί��l�rg��A�ͽ��!/��7�������f�6�Ͻ:���p�t��3�xÌ���&;@;�<�==�V=�;�=t �=l�=*��=�d�=R�=���=�ȹ=�R�=X��=kI�=:�I=�.=���< pܷБ���$�:4r��ܡ�_�ǽg�罺���)l�C������j�Ὦ���K����W�J��dğ��'��   �   �kL<0�< �8��_�Hi���mK������ޭ��ȽE�׽��ܽ�yֽ��ƽ�h���풽��f���$��bļH��`E�;��<=�N=|�}=-w�=��=屩=(�=:�=N�=I�=zs=<�A= i
=P��<`N�;K2� @׼�@*�^;g�G�����o⽽�˽z8Ͻ�Wɽ#�������A~���5��ڼ��-���;@M$<�   �   @�=|h�<Ĥ�<x@%<�����I��b�ZX����:Ę��Z�������t��������k���@����$����#��y;xԑ<J� =~�3=@�^=��=��=�ٌ=�l�=��y=�=V=F[(=D�<ng< �� �b�ۼd���.I�� o��_�����&S���y������V��@�t���A���`������XOP<,��<�P�<�   �   ZwR=�BH=��-=D�=�<pD�; � ���ƼBo�4�D�g�0�~�@���b���������V�r��QW���2����[���#���<(ɹ<F=��3=*cK=*sR=�>H=�-=X|=8��<�;x� ���Ƽ�u���D��	g��������b��������:�r�@MW�Z�2� ���O��p� <0Թ<^=T�3=�gK=�   �   �ی=|n�=��y=�AV=�_(=,N�<�g< �{�8�b�ۼ���+I���n�o_��ě���T���{������Y��R�t�ԢA�$��m���i�� 9P<��<�G�<̝=�_�<,��<p+%<�*���V���
���X��"��Ș�d^������Mw���
������k��@�B�������#�`gy;�ޑ<<� =0�3=�_=�=��=�   �   �)�=�;�=�=�J�=ds=v�A=~m
=$ʞ<�o�;@<2�L:׼�>*��:g�H��q����佽�˽�;Ͻ�[ɽ�&������\I~��5��"ڼ��-�`�;8:$<�YL< < `�8H`�`u���tK��􋽲⭽�Ƚ�ؽ��ܽ�}ֽݲƽ&k��E@�f�v�$��_ļ���@_�;X�<=�N=X�}= y�=���=���=�   �   ���=B��=ʹ=�S�=���=K�=��I=�1=Ď�< `ȷX����#��4r��ݡ��ǽ܉������m�:������u�Ὀ��5O���W����\Ο���'�PK�  :�ؤ�����Tl��j��	�ͽ�!�V1��9�	����`j��ϽX���&u��4�XÌ� �&;(?�<v@=܄V= =�=�!�=ym�=���=�e�=�   �   h��=�L�=$��=/<�=L��=Th�=y=n'8=�~�<��;�9����"�N���U������=
��+�0�#��>%����S��/����ͽ'Ş�h�g�\O#�\2��ռ0���<J.��x�Nڪ��Bݽ������x*��0�R6.��#�<�������������0"���i���<���<ܧD=J��=R:�=xɴ=BP�=|��=���=�   �   v��=8k�=�Z�=�M�=2�=��=�D�=V=�= �(</u�h�.����P�нA��.��3�t\?�*�B���<�T.����Y�����˽G���El�pH<�Ο-�hSB���x����q�ٽn��/�#�4Y:���I�x�O���K�~:>��Y(��g�T�ٽ�6��n0��'d��9J<�=�Ab=f�=d��=�?�=�_�=�8�=���=�   �   ���=���=0��=$�=��=��=�D�=�i=�=��C<�l���<��C��Ɇ�Փ�|�0��uG���U�o>Z�"_T�- E��.�<����r�������@rq�
�a�&"x����1�ƽ���t��ʨ:���R��c�@i�Z�c��T�K);�3��-d�8��^@� cs�XSb<�~=.�t=BR�=D^�=�=n�=��=V	�=�   �   ��=x�=�f�=@��=��=�d�=1v�=`]s=R=��M<������G�Ϊ������d%<���T�3ud�[�i�F�c�	T��|<��> ������Ͻ�ʤ�N����e���5��9����۽j��*�vbI�N�b�"�s��zy�Ŝs��eb��G�3�%�����Y���p_L�,J��xBj<hG%=n=�v�=&�=���=(��=6�=T|�=�   �   x��=0�=N��=lW�=޻�=@-�=p��=!�=�^=��=`�<��|�(iּ8WG�8z���󵽇�ӽ�潪��k����ӽ7q���g���Q���i�Fe�x���ܧ������ǗL�G����%������;�ھm|߾�ھj�̾DT���B���'|��Y>�V��I��@���<��)=��=�q�=���=,�=t��=d�=�   �   �s�=���=�=8�=,>�=�~�=$�=zi�=2�W=�5=���<P9��Բּ�E�[���N���9Ͻ�(�d|�@D߽�\ͽ4��҂�����'_�4_Z�~�y�������ܽ���G�&�}������1��2�Ⱦ�L־j�ھ�O־W�Ⱦ����P����v�nQ:�|$ �%H���j漀�%<R/*=E��=�}�="[�=|�=��=��=�   �   В�=8�=�D�=0\�=O��=�C�=�h�=>)�=r$C=���<�T<�Nһ�ټPK?�Vm��G������5ѽ��Խv�̽Խ���(��e���(_��@��Z;�
=Y�֩��0�ǽ�7
���8�*�l�점��訾d����mɾB�;Ţɾ,Ἶ��������h�.�.��n��^˼��><z�*=��=�o�=�R�=���=���=��=�   �   P��=���=lc�=���=@��=���=n��=V�X=-=Dý<p��;8F,�8"�ک9�T{��T���孽�/�������a������5��"gY��z,�6��
�@&���f��V��S��P�!��yQ����*[������q��'ɹ��������~������1RQ��A�?1ֽ �t� B��H�]<�*=_�=��=��=�V�=P<�=`~�=�   �   ���=+��=T�=��=$G�=�σ=�uT=$L=4,�<p�1<�b��ّ�л�2�9���j�KA��$ۖ�:����\������u�vXF�J��4�׼LW��D ���ȼ~c��e{�j���@���//�=tZ��5���~���P��lw������&˓�d\��A�a���5�h!��_��P�N��I{�Ht<x�$=v�y=h��=�
�=>��=�_�= 1�=�   �   �O�=��=���=�-�=@Kp=t�;=2g=�<�F�;��؂��8��`"���E�"�b� 4w�7���O~�T�m�ƱO��'��!�@���
���� n����ɻ`���n����|ǽb��.���P�h_m�fV���\���c���hu��Z\�V/<�B����#J��j*+���>���p<�7=��d=�"�=���=]��=���=j��=�   �   vA�=*L�=�:�=�JP=��=ܑ�<���;���Tॼ*b ���%��eB��;W�lmd�hj���g��h]���I��C,�`���5���%� �z: P&<ذ�<4-�<8�Z<��D;��`���|ӂ�f/���Z ����*v6��G���O�g�M�zC��90����������� �����1)�رD<�8=&xE=Ff}=�-�=Ϣ=pD�=�a�=�   �   G݁=ܫ_=X-=8�<��'<`���l�ʼ>r%���Z��v���T��7$��6���W����S��8�j�b�H�<M!��������:���<���<��<=DE=��=�	�<��-<p8������cf�8���ٽ����2�����f�K!����+���ĽVA���AZ��F��0K����;xj�<��=4�M=lsu=6�=r�=���=�   �   ƃ7=��	=�e�< ԇ�h�����-��w������\���޿ҽ��ٽr�ֽ�Qʽȯ��؝����~OG���	�|����d� �2<$��<�=�8=��Q=p�Z=8�R=��7=��	=�t�< ����諼V�-�r������y���?�ҽ��ٽ�ֽ-NʽH����֝�����PG�ޖ	���� �d���2<��<4=T�8=»Q=V�Z=��R=�   �   ���<0�-<�Y�����nf�6#����ٽT��,6�Ɖ��i��#���/���Ľ}B���BZ��E��'K� ��;�q�<r�=B�M=�wu=_�=��=l�=�߁=α_=�^-=8�<`(<�9��@�ʼdh%���Z�6r���P��� �����������R��h�j��H�2P!���!���b��p�<8�<L
�<�=�?=�=�   �    3D;�a��#��؂�45��^ �H���y6���G�*�O���M�V	C�P<0��������N���������,)���D<d;=N{E=�i}=p/�=�Т=lF�=�c�=�C�=�N�=Y=�=QP=��=䠳<`��; ���Х�[ �z�%��`B�D8W��kd�6j��g�`k]�v�I��H,����@��8&� *y: :&<Х�<�!�<ȀZ<�   �   ����v�����ǽY��`!.�O�P�$cm�IX���^��me���ku�2]\�I1<������K���*+���>�8�p<�9=&�d=&$�=r��=켸=W��=*��=�Q�=.��=Ҷ�=d0�=�Pp=T�;=Tm=P�<�u�;0l�z�����l"��E��b�06w�퍀�\S~�R�m�*�O��!'��,�K����
� ��@#����ɻ�   �   �i�m{���������2/�nwZ�;7������ZR��$y��F����̓��]���a��5�G"��`���N��G{� t<0�$=��y=���=�=���=�`�=�2�=*��=���=(�=��=EI�=�у=dzT=�P=�4�<�1<@�a�֑������9�6�j��B��ݖ�n���!_��;���b#u��]F�z��t�׼�a���
����ȼ�   �   ��f��Y��-���!�[|Q�t����\������Ds���ʹ�@
��ݘ��r�������>SQ�~B��1ֽP�t� A��`�]<r*=�_�=��=��=�W�=V=�=t�=t��=4��=�d�=���=ͅ�=x��=��=n�X=�/=�ǽ<p�;�B,�$"漶�9�0{�6V���筽�1�����d��$!��C8���kY��~,�~:���
�X&��   �   *�����ǽa9
�n�8�9�l�	����騾�����nɾT�;��ɾ�Ἶ\��X���Th�}�.�%oｕx\˼�><��*=��=rp�=eS�=h��=t��=��=���= �=zE�=*]�=T��=�D�=�i�=2*�= &C=<��<��T<�Lһ��ټXL?�+n��m��c���7ѽ>�Խ7�̽����P*���f��,_�v@�\^;�"AY��   �   ;�����ܽ;��6�G���}������2����Ⱦ.M־��ھNP־��Ⱦƣ��f����v�FQ:�>$ ��G�� h� �%<�0*==:~�=�[�=�|�=�=�=Rt�=(��=��=��=�>�=R�=��=�i�=��W=b6=��< ;���ּ�E����hO��b:Ͻ�)�f}�HE߽�]ͽ5��܃��<��*_��aZ�V�y��   �   �ݧ��㽮��p�L�����&������;�ھm|߾��ھ6�̾�S��2B��'|��X>����H��`���<�)=l�=|r�=ݥ�=��=���=��=���=f�=x��=�W�=���=P-�=r��=�=�^=^�=��<`�|�<jּ�WG��z������ӽV���콚��+�ӽpq���g��
R����i�je��x���   �   �����ܽ ���G� �}�Э���1����ȾL־��ھ"O־��Ⱦ������2�v�P:�9# ��E��0c�X�%<2*=p��=�~�=�[�=�|�=L�=(�=xt�=P��=��=��=�>�=��=��=Hj�=��W=�7= ��<�,����ּ E�|���M���8Ͻ�'ὂ{�hC߽�[ͽh3��>���@��D'_��^Z�n�y��   �   ���`�ǽF7
���8�D�l�U����稾z����lɾ�;�ɾ�߼�l ������fh��.�:k｀늽 S˼p?<��*=��=6q�=�S�=ػ�=ƫ�=��=��=V �=�E�=z]�=���=E�=Dj�=�*�=�'C=���<��T< 1һ��ټ�G?�jk��P��
����3ѽ��Խ��̽"���'���c��F&_��	@��X;��;Y��   �   ��f��T��U���!�FxQ����Z������8p���ǹ�3������ǥ��m���3OQ�#?��,ֽЀt��3��H�]<**=Xa�=��=u�=HX�=�=�=��=���=���=&e�=b��=N��=��=ω�=ZY=^2=<ν<P!�;x/,����9�r{��Q��㭽�,�����_��^���3��,cY��v,��2�2�
�|&��   �   �_�a{���������-/��qZ�4��}���N��vu������ɓ�gZ���a�K�5�M�*Z����N��({� 1t<��$=��y=ǔ�=�=6��=�a�=3�=���=C��=��=r�=�I�=�҃=0|T=�R=�:�<8�1<��a��ʑ���v�9��j�=��hז�����(Y��K����u��RF�<���׼O��������ȼ�   �   ����i�����yǽ��U.���P��[m�hT���Z���a��$du�tV\�L+<����>�'D���+���>�X�p<�>=��d=�%�=y��=���=���=���=TR�=���=V��=�0�=Rp=�;=Zo=x�<Џ�;0K��o�����"��E��b�+w�ڇ���F~�Z�m�4�O��'���4��H�
�@[��܉��oɻ�   �   ��D;��`���uς��*���W ����vr6���G�L�O���M�C��50����sy�������։� 
)��D<^@=E=~l}=0�=�Ѣ=G�=hd�=CD�=8O�=�=�=>RP=�=,��<��;���$ʥ��V �B�%�ZZB��0W��bd��j���g�_]�|�I�Z;,�Z��'��H�%� |:0f&<$��<�6�<ЬZ<�   �   t�<@�-<��Ķ��*Zf������ٽ^���.�_���b������#�B�Ľ^:��T5Z�d;�K��.�;{�<�=�M=�yu='�=V�=��=l��=Ĳ_=�_-=X�<�(<�,��8�ʼ�e%���Z�&p��N�����䒓�H���N��t�j�@�H��C!�`t鼘��p���<��<��<J =:J=��=�   �   �7=@�	=$��< P�׫��v-�l�����?�����ҽ��ٽ �ֽTFʽ����Vϝ�1����CG�V�	�����^d�p3<���<T=��8=�Q=� [=,�R=��7=h�	=�v�< ����櫼�-�q����������^�ҽ8�ٽ8�ֽ�JʽJ���ҝ�직�:EG�j�	�(�� <d��3<(��<� =x�8=��Q=:[=�R=�   �   R�=�_=�d-=0"�<�-(<�����ʼ�\%�&�Z�ek���I�����{�������7L����j��H��D!�y�������P<���<��<V=FF=��=��<з-<�4������bf����P�ٽp��$2�����e� �f��E(�ʿĽ�<��r8Z��<�K�@7�;�~�<r�=��M=�|u=��=��=��=�   �   �E�=Q�=@�=<WP=�=��<��;`j�̺��TO �D%�JTB��+W��^d�j�F�g�`]���I��>,�<���/����%� �z:HU&<䲃<�.�<@�Z<��D;�`���ӂ��.���Z �r���u6�d�G��O���M�fC��80�@���}������������)�H�D<HA=��E=vn}=�1�=
Ӣ=bH�=�e�=�   �   �S�=*��=��=�2�=�Vp=�;=�t=4(�< ��;�㻄e��p��"�
�E�B�b��+w�ӈ���I~��m���O�~'��l=���
� ���X���ɻ@
��Tn�����|ǽ1���.�u�P�_m�.V���\��ec���gu��Y\�#.<�����	��F���#+��>���p<�>=��d=&�=J��=���=��=���=�   �   ���=f��=��=��=�K�=�ԃ=r�T=NW=8C�<��1<�]a��đ�����9� �j�>���ؖ�,���[��f���Ju�(WF�J����׼V��8���(�ȼc�&e{�(��� ���//�tZ�j5���~��dP��4w��k����ʓ� \��T�a���5�< �]����N��3{��*t<
�$=��y=��=��=���=Nb�=�3�=�   �   ���=\��=f�=���=���=|��=P��=rY=d5=�ӽ<�4�;�',�@漘�9��{��R��$䭽a.�������`��8���5���fY�z,��5�
��&���f�PV��%��:�!��yQ�����[�������q�� ɹ����w���7�������rQQ��@�o/ֽ �t� :����]<*=!a�=��=��=�X�=F>�=f��=�   �   <��=� �=NF�=&^�=z��=�E�=:k�=�+�=�)C=d��<��T<@'һ�ټLG?��k����������4ѽ��Խ��̽x���P(���d��B(_��@�nZ;��<Y������ǽ�7
���8��l�᠐�~訾S����mɾ*�;��ɾἾ�������Bh���.��mａ튽�X˼ �><�*=F�=q�=�S�=��=���=8�=�   �   �t�=l��=��=8�=D?�=��=`�=�j�=��W=�8=Ԝ�<@&��x�ּ�E�����M���8Ͻh(�
|�	D߽x\ͽ�3���������'_�_Z�Z�y�������ܽ���G��}������1��*�Ⱦ{L־^�ھ�O־F�Ⱦ~���6����v�-Q:�4$ ��G��Hh漨�%<�0*=니=<~�=�[�=�|�=8�=(�=�   �   
 �=�C�=>��=��=L
�=���=@�=z��=
�w="G=,C=��<p(< / ���g��żʎ�Z���M�|3��M���㼰�м��޼6��2Z�򣨽�]���\9�0M��2U���Uվ�| �_5���#��.�v�1�t.��#�`�����.Ӿ��� )r��"�P��Jj�ا<�<8=�%�=�j�=�T�=*��=( �=�   �   �S�=>�=��=��=�
�=��=6�=���=L�k=��;=�
=���<��< �f��p�("ż`=���Y�L��TT
��_��h�ӼP����ͼ~��z�O��z������ܡ4�D�z������о'���bX��� ���*��D.���*��� ��+�������ξf���Z�l���P���
�P�-<�:=�C�=��=�G�=z_�=n��=�   �   B�= 0�=L{�=�=�ܸ=gf�=�c�=>�t=6kG=JO=`k�<�gp<�cg; R�Ls���ż\��Д�HQ�x���ɼ ����P��Tԛ�~ۼC1�������Ὗ�&�H�i�j%���LľY"��		�L��aR!�Ϣ$�`!�����
	�p�쾜�¾5��y^�����٦�d��X[<�?=�[�=#�=���=��=2y�=�   �   l��=���=v��=�A�=���=B�=Ҿc=��5=x<=�X�<h�L< IC;�W��hg_��X���Aͼ伌��p�ռ ���,���(�>�P������������h�sZ���s�L�N�|���ᐰ�f&־�/����	�u����X��M�	�a�����־
m��Y<��jYG��+�l���Ԣ���ˍ<�aE=@Ò=���=2��=<��=Ds�=�   �   ���=�ͺ=,��=�e�=�,s=��>=�v
=���<�)< ��9X��X,u�`秼�;ɼ�*޼ĸ�̖޼��Ǽ����`�_��M滀��`q3;`A*;�	X�X���x� ��a���T�r�,�-�k�Z���+��am׾K�ﾹ������: ����X)پ>���_���m��J+���ݽh�h�h__�\�<4�J=h��=q|�=PU�=xE�=�i�=�   �   �í=�i�=�@�=�M=\B=,��<��;���d�,����g�L&�P�+���(�"_��e�(,�۴�(�f�p��� eH;�:*< �y<T��<��?< и9hu��l�B�?o�������<�w��n��C����Ǿk�վ��ھ�־��ɾ�赾&|�����NeE����W���@�/��O��4��<
�K=�ŋ=�0�=��=�=��=�   �   C!�=�Eh=�(=���<�6�;��~��
�5L�&���Z�����k-���Ӓ��W��l�f�f<����.��P+��}�:h�K<Pð<���<���<`��<�]�<@�;R��^[��?���<��=��lm�5����u��JA���𮾡��������'{�4M�6c��\޽; ��o��@p�:(��<�F=�v�=��=N��=��=��=�   �   >1L=�
= }_<���O��o�������ͽ����w���9��ޖ��c;��ǽ�*�������}8�Tdݼ!����;�w�<F)=�"=�3=N^/=|I=<Ͼ<�kx;����]�肹�
���+,��5P�"�m��������r���bx��K`�3A�
���d������J��⡼0��;���<R@9=xn=�ׇ=:Î=�u�=֢{=�   �   ���<К�;�|����B��M�����j��^%�f16��>�n�=�֣4�$$��\����zz�rK��S���;�j�<V�!=�dL=e=�i=�Y=�b1=�<P��;8h����B��F��8�ེf�FZ%��,6�l�>�:�=��4��$�p�_�R�	z��I��S���;�f�<��!=@aL=Ne=��i=XY=t\1=�   �   ��w;�����]��������d0,��:P�<�m�����.���t��6gx�vO`�@A�f��?h�����*�J��䡼 ��;��<~B9=:	n=�ه=.Ŏ=�w�=>�{=�7L=t
=Р_<`���C���o�Á��c�ͽ���qp���2������"6㽾�ǽ|'��󲁽�{8�DcݼP!���;�r�<&=`�"=�3=tY/=�C=���<�   �   �b���'[��E���@��=��qm�ѷ���x��D����8��������b*{��M�e�p_޽�!���q���o�:��<��F=�w�=/�=���=��=�=�#�=XLh=��(=�<���;�X~�V�
��(L�Ҷ�U��N����(���ϒ�}T���f��	<��~�h/���%+� 2�:�K<��<�{�<���<��< R�< l;�   �   ��B�pt��ۗ���<�Tw�!q���ԷǾA�վ��ھ��־<�ɾ�굾�}��� ��=gE����������/� R��x��<T�K=qƋ=�1�=��=��=��=ƭ=gl�=�C�="�M=<J=x��<�g�;@��Lݬ�����^_�&�n�+�^�(�P\�`d�,,��ݴ�H�f�Ь��`/H;�+*<h�y<,��<��?< Ե9�����   �   �e���Y�x�,���k�q�������o׾���f���ޠ�p �� �4+پ���a��̦m�L+�N�ݽ��h��`_�X�<\�J=2��=^}�=xV�=�F�=k�=���=�Ϻ=���=�h�=3s=��>=�}
=�Ͱ<8*< ��9P��u�hߧ�6ɼ�'޼ ��8�޼ȷǼ@����_��h滀��� 13;��);�XX��눼B� ��   �   $^��v�
�N��������z(־ 2��#�	����
��[��1�	������־�m�� =��EZG�v,�����Ģ���̍<�bE=�Ò=\��=��=H��=tt�=̑�=R��=G��=�C�=��=��=��c=ą5=`A=b�<��L<`~C;�C��a_�\W���Bͼ<�$�� �ռ����8���X�>����(��t��Ƙ��h��   �   ��ὃ�&���i��&��>Nľ�#�
	�-��;S!���$��`!���t	�.��$�¾����^����٦�0��[<�?=^\�=�#�=T��=܂�=z�=C�=61�=�|�=l �=l޸=�g�=fe�=p�t=DnG=R=8p�<�op<@xg;�L�<s�� �ż���\��(S����ɼH���dV���ڛ�0�ۼ@G1�����   �   +���<�4��z������оA����X�
� �(�*�YE.���*�(� ��+������ξV����l�ĳ����~
���-<":=0D�=Z�=0H�=`�=��=pT�=��=R �=Ԗ�=��=��= �=���=��k=��;=�
=о�<@�<��f�Pp�l#ż(?���Z�����U
��b��нӼ4���ͼ����O��|���   �   <_��v]9��M���U��lVվ�| ��5���#��.�u�1�a.���#�/�������ӾD��8(r�$�"��N���g���<p>8=&&�=k�=2U�=���=z �=T �= D�=n��= �=p
�=���=L�=z��=�w=�!G=�B=�<�(<�8 ��g�H�żX����\N�4�0N�P��t�м�޼����Z�����   �   7����4�b�z������о����3X�>� �N�*�|D.��*�Y� ��*�������ξh�����l��������r{
���-<� :=�D�=��=xH�=<`�=0��=�T�=�=t �=���=��=��=9 �=���=b�k=��;=�
=l��<�<�ef��p�ż�:��ZX���>S
��]���Ӽl��D�ͼ�����O�={���   �   ��2�&���i��$��Lľ�!�Y		�����Q!���$�2_!����
	������¾����^����\֦����[<�?=Z]�=n$�=���=D��=hz�=HC�=|1�=�|�=� �=�޸=Lh�=�e�=l�t=�oG=�S=t�<�xp< �g;�2��k��̍ż��񼰑�`N�4��$�ɼ���LM���ћ��{ۼ�A1�����   �   �X���r��N�����Џ��%־D.��	�	�c��Ȝ�!���	�����~�־k���:��XVG�g)�1���ܔ��׍<xfE=DŒ=Z��=���=���=�t�=0��=���=���=�C�=h��=�=��c=.�5=C=hf�<p�L<��C;�$���N_��L��7ͼ��� �漤�ռ(���y��x�>�8��������R��x�h��   �   �_���Q콳�,���k�󘗾t��Wk׾���"���/��� ����&پ�	���]���m�aG+�	�ݽ��h�8?_��)�<ޞJ=ϓ�=�~�=XW�=tG�=�k�=3��=`к=��=�h�=�3s=��>= 
=(Ѱ<�*< ?�9X��8u��է�+ɼ,޼H��T�޼$�ǼP�����_�@)� �����3;`w*; �W��و�ږ ��   �   .�B�l�����O�<��w��l������u�Ǿ��վ��ھ��־��ɾ�嵾ny�����aE�������Ҽ/�P	��� �<HL=Aȋ=43�=��=n�=]�=�ƭ=�l�=pD�=�M=TK=�Þ<�s�;ت��ج�(����[��&�J�+�^�(��U��\����̴�8�f�`f���H;@N*<�z<l��<(�?< ٺ9|l���   �   �F��T[�{;��1:�l�<��hm�㲌�=s��n>�����������
���!{�PM��^�iU޽����Y�� ��:���<��F=�y�=��=���=x�=��=�$�=RMh=��(=䯾<P��;�S~�̷
��&L�p���S�����Y&��4͒�hQ��
}f�<�Bv�����+� S�:�K<�Ͱ<$��<���<��<�f�<�+;�   �    �x;\���N�]��}��ș�(,�]1P��m�J����
���o��]x�4F`�A�Y���\�d��J�@͡���;��<\G9=�n=�ڇ=$Ǝ=�x�=f�{=�8L=^
=��_<����B���o�
���z�ͽѵ� o���0�������3��ǽ#$��>����s8�XRݼ�� �@��;0��<�.=�"=�3=�b/=N=Xپ<�   �   ��<�;�W����B��@��%�ཥb��U%��'6�<|>���=�ؚ4��$����齈경P�y��=�X�R��M�;�v�<��!=�gL=�e=��i=�Y=�c1=��< ��;|f����B�9F�����df��Y%�P,6�ƀ>�j�=��4��$��H
���z�"B�x�R��D�;w�<��!=\iL=�	e=p�i=Y=�g1=�   �   �<L=�#
=�_<H���8�<�o��z��m�ͽ\��jg���)������@-�\zǽ���䫁�o8��Lݼ� �@��;���<,-=��"= 3=�_/=�J=Ѿ<�xx;��P�]�����М��+,��5P�ņm�ƶ��V��)r��bx��J`��A�����a�i�֓J��ԡ�p�;,�<�G9=�n=�ۇ=:ǎ=z�=ڬ{=�   �   W&�=�Qh="�(=���< ρ;H.~�4�
��L�f��vM������� ��FȒ�?M���vf�N�;�(s����p +��<�: �K<�ɰ<T��< ��<��<�_�< �;�P���[��?���<��=��lm�����u��A����V��H��x��	&{�
M��a�Z޽P�� c��@7�:���<J�F=z�=�=Б�=��=*�=�   �   ȭ=�n�=�F�=��M=�Q=�Ҟ<`��;����Ŭ�D����R�\�%���+�P�(��P��Y�d�˴�H�f��p����H;0E*<��y<��<x�?< 0�9(t���B��n�������<��w��n��*����ǾD�վ��ھҫ־��ɾT赾�{�����FdE�~������J�/�'��h��<.L=)ȋ=v3�=n�=L�=��=�   �   T��=�Ѻ=Ɠ�= k�=9s=d�>=^�
=�ް<�,*<�`:pn���t�h˧��"ɼ ޼d�弤�޼X�Ǽ�����_��8��׉���3;`Q*;��W� ߈�� �}a��`T�T�,��k�K�����Mm׾3�ﾚ���~��" �b��)پ����_��F�m��I+�
�ݽ��h��O_�\$�<J�J=}��=�~�=�W�=H�=�l�=�   �   ��=���=���=jE�=2��=*�=x�c=�5= H=dp�<@
M<��C;��@C_� I���4ͼ8����漘�ռ���||����>����Ȋ����>����h�IZ���s�;�N�q���ؐ��Y&־�/���	�i����F��7�	�-�����־�l��<���XG�O+�������Xэ<�dE=�Ē=/��=���="��=ju�=�   �   �C�=2�=�}�=�!�=�߸=�i�=@g�=��t=�rG=�V=,z�< �p<��g;`#�i��H�ż\���� O�<��d�ɼl���|O��hӛ�L}ۼ�B1�v�����ὓ�&�:�i�c%���LľQ"��		�G��YR!�Ţ$�`!�w���
	�J��s�¾��^�v���ئ�����[<�?=�\�=$�=���=T��=�z�=�   �   �T�=2�=� �=X��=l�=��=� �=���=�k=N�;=4 
=xĭ<X�<@Sf�(p��ż�9��JX�B���S
��^����Ӽ���,�ͼP��T�O��z������ա4�=�z������о%���`X�� ���*��D.���*��� �{+�������ξN���*�l�������~
���-<�:=
D�=K�=,H�=`�="��=�   �   *�=���=8�=ط�=��=I��=|Ù=!��=X�m=&M=h�.=��=x	�<�G�< ;�<�<�*[<��M<��P<h�X<8�R<�#<��,;8�?����ȡ��������G�D��U�ǾDU�Bn"�G�A��]�8�s��퀿]���뀿��s�z]�FYA�^�!�X�uFþ.\����2��(Ľ��� Gz<v�R=۞=�d�=��=���=�   �   ���=���=R�=���=|�=�=���=��~=��[=��;=��=��=L��<Ğ�<0��<��g<x�M<��H<8�S<��b<��a<p8<�;�#"�z~	�5֎�`7��ڱB�)��~zþ����Z�G+>�@�Y��ao�<O}�n��O}�7Wo���Y�t�=�K���$���\���f���.��=������D1�<��T=��=��=���=$3�=�   �   ��=$�=3��=l��="Z�=(ڌ=�p=�I=��%=<K=U�<��<���<(�R<H%/<؊<8�!<�7<�Y<�j|<0L�<�/q<��
<p����ݼ�{��Q��W4�����冷���l�-�3��N���b��p���t�H!p��b�N�ՠ3�j��������}�r)"�?���Ӽ �<��Z=���=� �=Z��=`��=�   �   NM�=L߽=�ܫ=6�=��{=�7J=z=8�<l1�<�%<0p�; LN:���� �غ �7��s�:��;<8�Y<Ժ�<���<X��<`�v<`�f;���,G�	�����|8l��夾4�پ4}���#���;�?	O��b[��_�[�48O�Z<��#�me���ؾ����bc�2��A�����<�b=�P�=�e�=� �=xN�=�   �   �>�=x}�=E��=�{S=t-=�ެ<0��;��Ż���ȡ��������8��HG¼ p���\<�@!�����;��D<8ԛ<t�<���<x��<��a< w��t���Q��Rj��9G�K��}0��U��g���$���5��A���D��:A��L6�t4%��������⫌���B�&S�T}f�����`��<dRj=o�=�ɳ=*�=��=�   �   �Y�=8�n=��*=L�<�79;�t�������P��I�����4������%>��ҏ`�dx1��������������j
<���<�6�<,�=lO=�/�<�.<0�Z�JNE��F½�v��ee�%����žª�6�
�O��~6#�Ш&�A�#��/�/�����FȾ���*�h��f�3ỽ�G!� �+; =,Yo=�}�=���=�=᧤=�   �   �T=.�	=8+9<Haa��j$��e��H귽�\���(���A������W��Žͤ���i��i��҆��k�:���<���<�)=l�$=&Q=P�<`��;�)��|�}�F���+.���q�)���O���߾[(���?�Q=�����2��t⾤tþ�%��,�{���7��5��ۻ��$f��xK<$ !=�Lo=P��=�p�=tݕ=VɅ=�   �   ���<@�w;��Ѽ0�o�X���r���!��;���L�r�T���R�RPG�$�3�v$�����aۻ��~����B�HDF<T�<�[(=�sB=,�B=n�%=\��<��;,�򯎽˧�?/�(i������������|̾�Ѿ�	ξ�¾�(��b��@�w�d�?�J�	�أ��R�3�0Z����<6e,=�Vh=E�=,�=��s=��@=�   �   ���:�����팽���]���L�6u��֊�����/:������:L�� 3���,^��15�d�
�.}½8�k� Eȼ`�m; 3�<�/= kY=��h=�f\=*u2=P��<@��:����挽"��t��j�L�u��ӊ�R����6����]I���0��J(^�Z.5�̤
�{y½J�k�x?ȼ n;�2�<|/=�hY=��h="b\=fo2=���<�   �   �!�S�������C/��!i����������	��l�̾��Ѿiξ�!¾�+���	���w�\�?�t�	�Ȧ���3�Ha���<f,=�Xh=�	�=�=��s=��@=��<�*x;x�Ѽ܍o�������~!��;��L��T�V�R��KG��3�� ����!׻��~���:�(FF<tR�<�Y(=�pB=Z�B=n�%=���<@;�   �   j�}�!��(0.���q�+��������߾O,���A�M?�����5��{�3wþ�'��U�{�4�7�9��ս��dj����J<� !=^No=z��=Ir�=�ߕ=̅=��T=��	=XS9<�1a��\$�B^���᷽.�I�������=�����P�r�Žd���H
i� e��͆�@��: ��<<��<<'=8�$=�L=��<��;�:���   �   $L½|z��ie��'����ž>���
�N���8#�̪&�$�#�f1����H��HȾ:���l�h��h�+㻽�I!���+;H =RZo=�~�=��=���=��=�\�=��n=��*=<�<��9;d\��p����P��B����������Ů��9��f�`��q1� �������pv��l
<l��<x3�<��=L=�&�<�	.<��Z�WE��   �   m�l=G�&M��3��L��	�˹$���5��A���D�d<A�mN6��5%�
��؋�t���ެ���B��T�f�`�����<dSj=<�=�ʳ=~+�=��=.A�=!��=q��=0�S=�5=8�<�>�;ЈŻ����T���������\��8;¼�f�� P<�`��P��;��D<�ћ<Hp�<p��<�}�<��a<𡂻*��V���   �   "���;l��社��پ�~�3�#��;��
O�1d[���_�}�[�x9O�o<���#�f� �ؾ̑���cc��2�B��4���<�b=fQ�=�f�=��=�O�=�N�=H�=�ޫ=��=��{=T>J=�=�*�< @�<��%<P��;��O: ���4غ 7�@��: �;P<x�Y<��<짤<H��<��v<��f;Ġ��RG�����   �   Z4�۲�����γ�m�T�3�6N���b��p�˲t�G"p���b��N�_�3����
������}��)"��>����Ӽ��<زZ=R��=Z!�=2��=n��=
�=��=���=8��="\�=Y܌=��p=ԦI=\�%=�O=H]�<�	�<���<HS<�+/<��<0�!<��7<�Y<�e|<�H�<'q<ؑ
<�0����ݼ:�{��T��   �   n�B�"���{þq����[�,>��Y�@bo��O}�����O}��Wo�фY���=�T���$���\��lf���.�=������@4�<
�T=O�=���=���=�3�=���=|��=>�=���=��=;�=���=Ң~=
�[=��;=b�=��=���<h��<��<��g<��M<��H<��S<�~b<@�a< 8<���;�-"���	�.؎��9���   �   ��G��D����Ǿ�U��n"���A�H�]�j�s��퀿]��v뀿��s��y]��XA��!� ��Eþ�[����2�'Ľ��POz< �R=�۞=Je�=.�=���=l*�=���=|�=��=�=j��=�Ù=*��=P�m=�M=�.=6�=|�<�F�<�9�<8�~<([<P�M<��P<`�X<�R< �#<@t,;x�?�������2����   �   *�B�N���zþ#����Z�#+>� �Y�$ao��N}� ��\N}�rVo�ȃY���=����d#���[���e��l~.�>;��H����7�<f�T=��=��=ƅ�=4�=���=���=X�= ��=��=^�=Ԅ�=4�~=��[=B�;=�=��=���<���<���<��g<лM<�H<��S<��b<`�a<P8<`��;�$"�	��֎��7���   �   �W4�H���~���S��;l���3�EN���b��p���t� p���b��N���3�N���������}�7'"�w;����Ӽ��<`�Z=<��=�!�=���=���=Z
�=��=��=r��=`\�=�܌=L�p=��I=H�%=�P=�_�<�<d��<S<�5/<��< �!< �7<��Y<0s|<�O�<05q<�
<���,�ݼR�{�*Q��   �   ���J7l��䤾�پw|�Η#�i�;��O�a[���_�d}[��6O��<���#�d���ؾ���N_c�R/�F=��P㐼��<t�b=�R�=�g�=~�=cP�=^O�=��=2߫=6�=B�{=?J=n =�,�<�B�<��%<p��; VP:������׺ .6��,�:p5�;�"<��Y<t��<t��<,�<��v<�g;H���G�����   �   i�B8G��I���.��d��5���$��5�A��D��8A��J6��2%�(����Z�������·B�Mｪsf�������<�Wj=� �=�˳=L,�=:�=�A�=���=Ҳ�=�S=�6=��<�F�; Ż����������\�����3¼X^��p=<�����߆;X�D<(ݛ<�{�<t��<h��<0�a<�_��6���O���   �   ]C½�t��be�H#����ž�ﾤ�
�����4#���&�%�#��-�/����gCȾ�|��\�h�c��ڻ��=!� Y,;�&=_o=���=I��=j��=˪�=#]�=�n=��*=��< �9;�Z��d��d�P��A������y���E���F7��F�`�4m1����������G��0�
<ة�<0@�<6�=S=�6�<..<��Z�VIE��   �   �z}���� ).���q�ۍ�������
߾�$���=�9;����`.��z
��pþx"����{�$�7�.��m���,Q���#K<X'!=6So=6��=�s�=|��=�̅=ƐT=h�	=�V9<�.a�\$��]��U᷽~�s���/���<�g����N�X�Ž���i�z_������S�:ػ�<h��<.=|�$=U=x'�<��;����   �   ���k�����y;/��i���k�������x̾�Ѿ�ξ�¾�$������w��?���	�K���֦3��0��ŧ<�l,=�]h=^�=M�=d�s=6�@=��<�9x;ȜѼ�o�����|��~!�,;���L�d�T���R��JG�
�3��������Ի�v~�>��"� _F<<_�<|`(=xB=R�B=��%=��<��;�   �   ���:����@ጽg��X����L�ru��Њ�뵕�U3��=��E��@-��"^��(5���
�-q½B�k��'ȼ �n;xC�<�/=PoY=��h=�h\=�v2=���<�ڃ:����K挽���B��5�L��u��ӊ�#����6����I��20��Y'^�K-5���
��v½��k�@4ȼ@gn;�>�<�/=`oY=
�h=�j\=�y2=h��<�   �   ��< �x;�Ѽ�o�ы��|��y!�;��L�ȬT�'�R�tEG�$�3���G}���λ�(
~�V���kF<Xb�<�`(=vwB=؉B=N�%=��<��;�񼓯��v���>/��i�|���j������}|̾��Ѿ�	ξR¾R(�����N�w�Y�?�,�	�v���X�3��E�H��<�j,=
]h=��= ��=�s=�@=�   �   F�T=V�	=�t9<0	a��P$�)W���ٷ�-�߽�������r8����*G�z�Ž<�����h�VX�x������:࿌<���<�-=��$=bS=h"�<@�;�'��Ҁ}�����+.�n�q����:����߾=(���?�:=����J2��%�HtþT%��F�{���7��3������L]���K<�$!=,Ro=F��=t�=��=W΅=�   �   �^�=��n=��*=�(�<@�:;`E��n��^~P��:���򎽋򓽱���D1���x`�~d1�����v��`*����
<,��<�@�<��=�Q=(3�<x$.<��Z��ME�GF½�v�hee��$����ž���-�
�C��o6#���&�*�#��/���y��aFȾO��`�h�$f�w߻�8D!� ,;�#=�]o=h��=���=0��=��=�   �   �B�=[��="��=S=�==��<���;�0Ż<愼�t��t��ī�0��D$¼�Q�� )<���� �;� E<Tޛ<�{�<��<H��<(�a<�o��Ԃ��Q��:j��9G��J��r0��H��`���$���5��A���D��:A��L6�[4%�ˍ�ʉ�̗�������B��Qｄzf� ������<�Uj=d �=�˳=�,�="�=�   �   HP�=��=��=I�=2�{=�DJ=�&=�:�<LQ�<�&<��; R:�㝺 #׺ 5�@��: J�;�)<x�Y<$<��<8�<��v< g;�����G�������l8l��夾,�پ0}���#���;�8	O��b[��_� [�"8O�F<��#�Te�Ŏؾܐ��<bc��1��@���쐼X�<l�b=#R�=�g�=��=�P�=�   �   �
�=��=��=���=�]�=hތ=j�p=��I=��%=�U=Li�< �<�Ƅ<`S<�A/<�< �!<��7<xZ< t|<�O�<�4q<�
<�����ݼ��{�yQ��W4�����������l�(�3��N���b��p���t�>!p��b��N�Š3�Z��`��n��d�}�#)"�\>���Ӽ��<X�Z=���=�!�=���=���=�   �   ���=Ҕ�=��=���=^�=,	�=ƅ�=Z�~=��[=��;=��=<�=��<���<��<P�g<`�M<h�H<X�S<h�b<��a<�8<`��;x""�H~	�#֎�Q7��ֱB�&��{zþ����Z�E+>�?�Y��ao�8O}�l��O}�/Wo���Y�k�=�C���$���\���f���.��=��L����2�<z�T=$�=���=���=�3�=�   �   ��=N`�=Y��=PE�=�p�=B��=��=c=HG=´0=� =)=<�=�=��=��=� =*I(=�-=rq+=�=T�<ȜR<(�`�\�\�*A佯�B����TZ׾���}<�Zch�WQ������ɠ�� ���9��9�������ܛ���t�g���;�����ҾŅ���T0��=������T��<*&u=pͩ=��=�s�=�   �   ���=�'�=�^�=���=�r�=���=��m=�nK=��.=�M=�|=��<��<��<�;=�c=>u=�{"=�E*=ff*=�=�&�<0�f<�C�j�R��;ݽ<�=�������ҾIC��9�2>d��톿4O��q��������*����������9��������c��$8����[�ξ�p����+��s���,��@��<�Zv=�2�=��=X��=�   �   ��=�Q�=Ⱥ�=@��=�=F�U=��)=�'=���<��<��<P�l<(�x<�ď<`k�<x��<���<jQ=b�=8�&=H}=��=��<0�޻l15���Ƚ��/�T#���Nƾh���.��0X��������(^���5��fD��a=��
f��J���$����W�S?.���~�¾E���Mw�E���H�z����<ky=�/�=k��='��=�   �   ���=�b�=D�=p�a=Xb&=p��<��R< /�:���؊R��y� �l��3����;��*<���<?�<@�=�d=��!=J�=��<@Ð:�;�悔U���{t�銲�����(��SE�4-j�f���:���s��O��ل���T��5|���<j��6E�����A�S���Vk�t��ʁ��^��`�=��|=z4�=�S�=��=�   �   qٕ=�=y=F�7=��<`��;��A�$U０�2�(�]� �u�j5z�k���L�� �4�׼pK�@�:qt<��<��=K =T�=l��<��2<hR���d�����Z�N������Ծ(�M-�XdN�¿k��p��I݈�,u������䛁�^!l�/�N�5�-�x+��ԾF��H��j�t C���;
�=��~=�x�=�3�=�,�=�   �   t\=J =`�\<(�<�@���恽�v��VFؽ;@� 0 ������"�Խʰ���(5�������5��)p<�w�<�=�$=2�=�=�<��B�\6%��
���$$���z�yB��!�����.�dsH�{�\��i� <n���i�/#]��I�ɍ/����=�� ���z���!������x��H�G<-=6�|=P&�=l��=���=�   �    ��<��y;�dټ@:w�8Ľ�x�\a%�]?�^zP�b�W�&U��H��~3�p6��:�@��nc�|�ۼ�$�P��<\s=ؑ'=�(=�=�(Z<�%����v����@�K���&���l��I��ǆ#���4���?���C���?��F5��v$�7�r>�"μ�fQ����D����v��OW�4�<�;=Ut=��=�v=$�E=�   �    }6��L�����x���+��	[�ο��nÓ�����w���ɠ�YV���!���Vi�
h=����l�ǽ�xm�����К�;��<x�"=�E9=P{+=���<n�; ��9��,!�gL��Z�������۾e����l�-{�!��7�� [��� ��Z߾Ը�.��M,V�����@7);�"�<Z/C=�pd=^`=^>7=��<�   �   ����뤽����D�t���ߠ������Ҿ��Z��]k�XKվQ�����^�� �S�N����ŽXGP��Y� ��<��=`�B=XL=`�/=��< Ne9��䤽\��$�D����۠�{�����Ҿ-ᾼ���f�FGվ�}������[��S�S��`|Ž�AP��Y�ܙ�<F�=��B=L=|�/=T�< .\9�   �   �?��o%��L��]��狴��۾/���o��}�������e]��� �:^߾�ָ�<0���/V��
�$������ );("�<�0C=�sd=�`=HD7=��< �3� @�����������+�[�:�����������t���Š��R������Qi��c=����j�ǽ�qm��������;` �<��"=�C9=�w+=d��<01�;X
��   �   :�ｇ@�.���� ����뾡��U�#�g�4���?�C�C�O�?�0I5��x$� �fA�vм�#S���D���Nv�pXW�,�<�;=6Wt=j��=��v=ƤE=<��< :z;@Jټh*w��Ľ�s��[%�2?�tP��W� U�u}H�z3�>2��3�I;�� fc�d�ۼ@�纰��<ds=z�'=�(=�=8Z<L6����v��   �   ($�`�z�tE�������w�.��uH�/�\���i��>n�v�i��%]��I���/�����?꾔"����z�)�!������|��؜G<`�-=�|=�'�=v��=k��=l\=�(=Ⱥ\<��<�����ށ��m���<ؽe6�@+ �]���z�ｋ�Խ�ð�m醽� 5������o5� 3p<Py�<��=.$="�=t4�<��B��>%�����   �    �N�����֘Ծ��O-��fN�.�k��q���ވ�gv�����𜁿5#l���N�x�-�s,�\ԾL�j�H�l�C�`�;��=*�~=�y�=25�=�.�=6ܕ=�Dy=r�7=0)�<�C�;�YA��9�6�2���]���u��'z��k�T�L��� ���׼�K�@��: |t<���<�=$J =L�=��<��2<�^���h���
���   �   1t��������:*�nUE�,/j�g���;���t��P��̅��bU���|��>j�z7E�d���B�����Vk���ˁ�^��"�=��|=z5�=(U�=m�=�ó=@e�=*G�=l�a=Vj&=T��<��R< r�:�K�bR���x�(�l��`3�ສ��7;�	+<X�<<B�<��=hd=d�!=,�=��< :�:�A�������   �   �$���Pƾ��"�.�^2X���Ŏ���^���6��$E��>���f�����������W��?.�Y��ţ¾c���Tw������z� ��<Lly=�0�=n��=c��=���=dS�=м�=� �=��="�U=��)=.=���<h��<`�<اl<��x<�̏<�q�< ��<���<R=z�=��&=�{=��=�<0߻|65���Ƚ��/��   �   ����T�ҾD��9�-?d��O���d���(+��C���Y����9�������c��$8�����ξ�p��f�+��r��H)��`��<B\v=i3�=��=!��=���=�(�=�_�=솰=<t�=9��=֗m=�qK=³.=�P=d=d�<��<(��<�<=�d=�u=�{"=E*=�e*=f=h#�<��f<��C�b�R�c>ݽ��=��   �   ���� [׾��R~<��ch��Q������꠪� ���9��&�������oܛ������g�E�;����H�Ҿ���uS0�<��L������<�'u=!Ω=���=lt�=���=�`�=���=�E�=q�=p��=��=2c=LG=��0=� =�(=��=z�=�=�=, =jH(=6�-=�p+=��=��<�R<��`��\��B�ȶB��   �   ����:�Ҿ_C��9� >d�{톿
O��2�������_*��~��������8�������c��#8�����ξ�o��2�+�3q��x$��Ȓ�<j]v=�3�=��=X��=���=�(�=�_�=��=Zt�=T��=�m=6rK=�.=�P=�=��<@ �<Ј�<�==�e=�v=}"=@F*=�f*=�=�&�<0�f<0�C���R��<ݽ��=��   �   &#��vNƾ%�s�.�\0X����{����]��5���C���<��3e��s������|�W�>.������¾̂��u�����H�z����<�ny=b1�= ��=���=̂�=�S�=��=� �=��=~�U=T�)=�.=���< ��<� �<h�l<8�x<�Ϗ<�t�<��<���<PT=µ=�&=�~=��=�<��޻15�i�Ƚ��/��   �   �zt� ��������'��RE��+j�Ae���9���r��N������lS��{���:j��4E�
���>�����Rk���~Ɓ�0*����="�|=�6�=�U�=��= ĳ=�e�=vG�=��a=�j&=|��<x�R<@��:�D�0^R�H�x���l�`Y3������^;@+< �<XH�<�=�g=�!=T�=�<���::�
����   �   ��N����`�Ծ!��K-��bN�޽k��o��܈��s�����������l�ֹN��-��)��	Ծ�헾2�H�od��B��n;(�=�~=P{�=(6�=�/�=�ܕ=REy=4�7=|*�<PI�; WA��8�Z�2���]�`�u�&z�8�k��L��� ���׼��J� ��:؊t<���<�=�N =^�=���<8�2<�L���b������   �   �"$�ޘz��@�����d�G�.�FqH��\�V�i�>9n��i�c ]�I�O�/�����9꾿����z���!�X����d��(�G<f�-=2�|=@)�=��=)��=�\=�)=�\<��<���5ށ�mm��B<ؽ�5��* ����o��M�Խ=°��熽85�����.5�HDp<���<��=�$=��=4D�<�JB��1%�����   �   ����@�Y�������O��i����#�>�4�T�?���C���?�D5�t$���:�iʼ�NN���D�����v��'W����<�;=�[t=킃=�v=P�E=���<�Hz;�Hټ�)w��Ľs�\[%��?��sP���W��U��|H�dy3��1�42�{9��4bc��ۼ�)� ɗ<�x=:�'=�	(=�=�9Z<���T�v��   �   �4��>���K�0X������۾1���9j��x�v�����{X�\� �3V߾�ϸ��*���&V�`�]������`�);�2�<�6C=�wd=~"`=NF7=��< �3�&?�L���u�����+��[�!���~��������s���Š��R��2���Pi��b=������ǽ�mm����`Ӛ;T*�<<�"=(J9=|+=���< ��;l���   �   ^���ޤ�̝���D�R����ؠ�����N�Ҿ���{�b⾊Bվ;y���
���W���xS�~��sŽ�3P�@�X����<H�=ڟB=4L=�/=��< �f9����㤽2�� �D� ���۠�g���s�Ҿᾔ���f�Gվj}�����![��5~S�r��}zŽ�=P���X���<��=��B=�L=�/=� �< �k9�   �   ��1�6�\������� �+�j�Z�򸂾���������o�������N������Ji��]=�F��X�ǽ�bm�������;�1�<@�"=�J9=�~+=��<�z�;��켠8��!�CL��Z�������۾P����l�{��� ��[��� �|Z߾�Ӹ��-���+V�E�+���:��@y);�+�<�4C=�wd=�#`=:I7=�!�<�   �   ���< �z;�4ټw��Ľ�n�(V%�0?��mP�^�W�PU��vH��s3�{,��)�P2���Vc���ۼ�Z�җ<H{=��'=�	(=�=0Z<D#���v�����@�=������]��@����#���4��?�y�C���?��F5��v$��'>��ͼ�Q��ΟD�>���v��AW�@�<̛;=�Zt=X��=`�v="�E=�   �   \= 0=��\<�v<����	ׁ�Ae��D3ؽ9,��% ������｢�Խz���,ᆽ.5�����@�4��Wp<0��<��=�$=z�=�A�<`nB�`5%��
���$$���z�mB�������.�\sH�q�\��i��;n���i�#]��I���/����h=꾟 ����z���!�[���s��x�G<��-=�|=d)�=P��=���=�   �   dޕ= Jy=P8=�9�<@��;�+A�����2�,�]���u��z�B�k�$uL�n� �$�׼��J����:Оt<���<��=P =�=t��<��2<8P��)d�����H�N������Ծ%�M-�QdN���k��p��C݈�%u������ڛ��H!l��N��-�]+��Ծ𗾘�H�xi�*�B� !;�=��~=6{�=�6�=�0�=�   �    ų=8g�=�I�=p�a=vq&=���<`�R<@��:����4R�8�x�0�l��43�0h�� �;�++<l�<�O�<��=�i=,�!=ޛ=<�<��:;��>���{t�⊲�����(��SE�/-j��e���:���s��O��ӄ���T��+|���<j�p6E�����A�(����Uk���Ɂ��O����=f�|=D6�="V�=��=�   �   l��=�T�=^��=x�=��=Z�U=��)=�4=�
�<4�<��<��l<��x<<ڏ< ~�<�
�<<��<�V=��=d�&=�=h�=��<@�޻�05�x�Ƚ��/�P#���Nƾg���.��0X����􍑿%^���5��cD��]=��f��C�������W�D?.���b�¾(���w�����`�z����<�ly=�0�=���=��=�   �   ³�=2)�=y`�=���=:u�=l��=��m=uK=6�.=8T=0�=,&�<t&�<���<<@=�g=�x=�~"=�G*=�g*=�=h(�<0�f<x�C�.�R��;ݽ6�=������ҾHC��9�1>d��톿4O��o��������*���������}9��������c��$8����L�ξ�p����+��s���+�����<�[v=>3�=��=B��=�   �   Xu�=��=pD�=�ş=���=2�k=��D=��#= )
=܋�<i�<�;�<��<��=<�#=�:=H�P=.c=z5l=:|f=�J=t�=�_!<`O．G��&6+�Ub��	vվ���W(J���Uk��ݕ��[�пn[�Gvￖ���q�RI�)Yп M��L��|r����H�WI��Ѿ�l��z�<ꈽ��S=S��=��=�M�=�   �   n��=d��=|�=��=�
=4�Q=(=��=�E�<T��<�]�<���<�g�<Z�<��=�)=(~C=�Y=�ce=��b=pgI=.�=h�3<�c߼�:����&��>��e Ѿn�@yF�:b}�v���s���~Ϳp�߿Ǎ뿏��G��/�߿��̿�F���d���t|��EE�-{��̾�w��_z��σ� �^��!=��=�=�޾=�   �   m��=@֥=g`�=�p=d9=�2=p�<�=<@=�: �� �Z��욺��t;��1<�ޞ<te�<�2=�;:=�EP=�lV=H�E=z�=��g<ű�ܵ�����f#��H�ľL����;��;p����������ÿA�Կ8�9*��D�e�Կ�ÿSv��������o���:��T
�������w�����j��	":�S'=*I�=���=�e�=�   �   ��=)!�=�N=�	=�ـ<�zﺐ7��$���`#���6�x�6���$�n�����'��p�;t��<�W=��*=�5@=�H==�=�ٙ<�[X��}�����e�X���`D��+�ߠ[�����Ҏ��k���o�ÿ��ο�2ҿT�ο�Ŀ����y���Ъ��m?[��^*�6���⭾�]�֩��<�p��;��.=���=}+�=�e�=�   �   �g=4�&=hU�<��B�P��}R��Z��v���Mѽaܽȩٽ��ɽ󰮽�(�C�� ڼ@�Ļ��O<�$�<�P=*�-==�f�< �5�:�8��ٽ4�A��$��-%ܾ��XA��8n�띌�����ym��f���"K��y��S���bΟ�[ό�7mn��TA��{���ھN��Z;�Pƽ�+�x�b<��5=$~=��=��=�   �   ��=0u<8����oV������)���p��0�8
A�=�G�S�D�-�7�=#�J(�6=ӽu�����+�@m� �<��<zA=��="�<��
< 
ڼV㠽6���wx�v׶��i��}�#�ڤJ��Ip�ň��Օ��7���)���b��[�����p�d3K�l�#���������̹v�b��U����V���x�<�]9=i=`ql=-I=�   �    t�:>�ᒽc��e&�6�T��n~�3ۏ�˚���
3��ֱ���}���"`�|S4��)�����M��ۋ��<�7�<j4=:�=���<�����L��M߽ީ>��0���vɾ�o��`%�=E��a��w�!��6����9���mx�>Zb��.F��S&�FT��˾�d����?��h޽��A��L �p��<�s6=JJ=��0=\9�<�   �   ���6�����
��H����nQ��}[����վ @侉���_���׾��¾�����l���`T��J��ý*L�h�W��z_<X��<��=|K�<�w$<Ԕ������
��.YU�m�VI̾�� �����"2��zD�OP���T�ӴP��<E�<13�9��W��EϾ9�H[��a������ļ��2<&\=4�*=��=�b�< ���   �   ����6a���X�:���%�����羌4���S5���!� ��n��ڇ��뾀�¾	���?b���e����#&��
[��H�<b=(�=���< �9;���郥�F\���X�n�������q�羺1���<2���!������i�����¾D��P;b���'���&&�`�Z�J�<�=��=$��< ,9;��   �   W���^U������M̾� �m��&2�9~D��RP��T��P��?E��33�T;��Y��HϾ�󛾲[�"d������ļ(�2<�\=��*=��=�p�< �Ṕ��Ӊ����
�,H�!	��M���V��f�վ�:�K���Z��׾s�¾&����i��0\T�NG���ý�L��W���_<$��<�=DC�<�]$<����( ���   �   ��>��3��azɾ�q��c%�0@E��a���w��������X;���px�]b�#1F��U&��U��
˾�f����?��k޽d�A� c �`��<�u6=FJ=��0=�I�<���:pq�ؒ����^&�6�T�:g~�׏��ƚ�� ���.�����3z���`��N4�@�U���D�M�4Ћ��&<,:�<�3=��=8��<p7��B�L��T߽�   �   �|x��ڶ��m��߉#���J��Lp��ƈ��ו�]9��L+��4d��� ��q��V�p�M5K���#�>���B����v�޷�����Y��Py�<t_9=Ji=8vl=�3I=��=h�<�أ��_V�%~�����j���0��A���G� D�R�7� #��#��5ӽ����ܷ+�P�l��<L�<�A=��=��<��
<ڼ�蠽؇��   �   '��D(ܾ��VZA�8;n�`���%���o������L����������ϟ�\Ќ��nn�BVA��|��ھ@��H[;�]Qƽ�,�Дb<�5=�!~=��=|�=��g=��&=Hj�< �A�t���lR��Q�������Cѽ]Wܽx�ٽ3�ɽ5����芽�C�8ڼ �Ļ��O<�*�<�Q=��-=j=`�<@�5���8�&�ٽ��A��   �   ����3G���	+��[��������Ņ����ÿ�ο4ҿ��ο� Ŀ����A���p���d@[��_*��6��㭾�]����,�<����;��.=ڠ�=-�=�g�=u��=S$�=�N=�	=��<@	�h������fR#�
6���6���$����`
������pO�;X��<�Z=V�*=6@=,H==�=Lә<hoX��}����e��   �   (�ľ|��)�;��=p���������� ÿO�Կ9�,+俞E� �Կ�ÿ�v������o���:�
U
�������w�����j� T":TU'=J�=���=g�=0��=`إ=�b�=�#p=,9=F:=�%�<�_<�P�:�v� Z�  ��`8u;�1<��<�l�<(5=�=:=dFP=�lV=<�E=��=H�g<�ͱ������ ��$���   �   �!ѾP�JzF�ec}�������(Ϳ�߿[���￯��|�߿��̿�F���d���t|��EE�{���̾nw���y��΃���^���!=��=�=�߾=���=���=� �=I��=
=�Q=((=��=PN�<X�<he�<<��<�m�<�^�<��=D�)=�~C=�Y=�ce=��b=:fI=V�=��3<�j߼,=��s�&��?���   �   �vվ ���(J��󀿡k��#�����п�[�^vￖ���q�'I��Xп�L�� ��/r���H��H��ѾBl���x��舽����U="��=��=2N�=�u�=:�=�D�=�ş=6��=��k=L�D=�#=2)
=���<ph�<�:�<��<�=��#=R�:=z�P=6c=x4l={f=.~J=��=W!<�T�MI��H7+�c���   �   � Ѿ��\yF�Ab}�k���S���IͿ �߿[��
�￮�뿈�߿�̿F��d���s|��DE�Jz���̾�v���x��̃�`�^��!=	�=\�=�߾=���=Е�=!�=f��=>=<�Q=V(=�=�N�<��<f�<��<�n�<`�<>�=��)=�C=�Y=�de=�b=pgI=ġ= �3< f߼�;��K�&��>���   �   �ľ��b�;�p;p�����'���ÿ��Կ37�>)俷C�R�Կ�ÿMu��ʸ���o��:��S
�������w�e���j� \#:0X'=K�=���=�g�=���=�إ=*c�=�#p=�9=�:=L&�<ha<�_�:�m��Z��噺 Gu;P�1<t�<`o�<�6="?:=HP=�nV=��E=P�=(�g<�ı�͵�����N#���   �   ��YC��F+��[�细����v���S�ÿm�οs1ҿ�ο3ĿE���+�������U=[�]*� 3��:୾d
]�����<����;�/=3��=�-�=,h�=���=�$�= N=��	=`�< ��p��|����Q#�@~6���6�ҷ$�j��`�������^�;p��<H]=��*=�8@=XK==�=ݙ<pUX�&}����e��   �   �#���#ܾ���VA��6n�䜌�_���l���󷿆I����������̟��͌��jn��RA��y�s�ھ�
��DV;�=Jƽ�"�@�b<��5=%~=��=B�=��g=��&=�k�< �A�h��DlR��Q�������Cѽ�Vܽ�ٽ��ɽj����犽��C��
ڼ0rĻ(�O<\0�<:U=��-= "=�k�<��5��8�ԏٽ��A��   �   Xux��ն�<g���#��J�?Gp��È�<ԕ��5���'���`�����d����p��0K���#�����K�����v�q��I����C��|��<�d9=�i=�xl=b5I=ܜ=Ф<xף�_V��}������j���0�iA�j�G��~D���7���"�H#��4ӽA����+���l�(�<��<6F=��=)�<�
<�ڼ�࠽_���   �   �>��.��tɾ�m��^%��:E��|a���w�j	��i����7��5jx��Vb��+F��P&��Q��˾�a��~�?��`޽��A� �����<{6=�!J=�0=M�<@��:�p�#ؒ�����^&��T�g~��֏��ƚ�� ���.��ܭ���y��_`�N4���ꃶ�<�M��ɋ��5<�B�<9=V�=���< ����L��I߽�   �   8��fUU��#F̾�� �*��+ 2��wD��KP��T�S�P��9E��-3�6��T�]AϾ�훾J�Z�]��󔽸�ü��2<rd= +=4�=�u�< 5Ṅ��l���V�
�
H�	��
M���V��R�վ�:�+���Z���׾;�¾㻧��i���[T��F�f�ý�L�P�W�ؓ_<���<x�=�T�<(�$<(��������   �   �~���X���X�}��������9/�R��;/�n�!������~��3�Q�¾B���4b���������&��/Z�\\�<:"=�=���<��9;>��r���\�q�X�_�������d�羳1���12���!�������N��K뾽�¾����:b�W�������&���Z��S�< =ƶ=п�<�:;����   �   |�����p�
�
H����\I��cR����վ�5��龇U���׾z�¾�����e��]UT��A��{ýL�X�W�ت_<|��<��=�S�<Ђ$<,���"���ւ�YU�^�JI̾|� �����"2��zD�OP�{�T�´P��<E�#13��8�zW��EϾ�𛾬[�a�r���ļ��2<�a=h�*=��=�|�< V޹�   �   ���:�f��ђ�r���Y&�	�T�$`~� ӏ���h����*������%v���`� H4�����{����M�����@Q<L�<�;=L�=���<������L�|M߽��>��0���vɾ�o��`%�=E��a��w���/����9���mx�&Zb��.F��S&�&T�Q˾�d����?�gg޽��A�  ����<�y6=�"J=��0=|V�<�   �   |�=`�<�£��QV��u��L��e���0� �@�ʵG�xD���7���"���g+ӽ������+��l��<P�<�I=��=4*�<Ȱ
<tڼ�⠽���wx�k׶��i��z�#�֤J��Ip�ň��Օ��7���)���b��Q������p�K3K�R�#�����_���V�v�ߵ�"����P�����<�b9=�i=|zl=9I=�   �   �g=��&=h{�< A�X�� ^R�~I���︽:ѽMܽ"�ٽ�ɽ�������JsC���ټ�&ĻP<�;�<<Y=��-=�#=�l�<��5���8�{�ٽ�A��$��&%ܾ��XA��8n�Ꝍ�����vm��a���K��p��G���WΟ�Oό�"mn��TA��{�x�ھ���Y;�Oƽ\)���b<��5=�$~=u�=��=�   �   ]��=�&�=�#N=��	=p �<��캸��t���vD#��p6��6���$���� �����;��<�b=��*=�;@=nM==  =`ޙ<�UX��}�����e�R���\D��+�ݠ[�����Ў��i���k�ÿ��ο�2ҿK�ο�Ŀ����p���Ȫ��\?[��^*��5��]⭾�]�&��6�<� ��;r�.=���=.�=�h�=�   �   L��=�٥=�d�=>(p=�9=�@=�4�<��<�k�:�����Y��ט�`�u;X�1<��<0z�<,;=�B:=KP=�pV=B�E=��=P�g<4ñ��������a#��D�ľK����;��;p����������ÿ>�Կ8�1*俼D�^�Կ�ÿLv��������o�t�:��T
�p���h�w�h���j� e":�U'=rJ�=~��=�g�=�   �   ۈ�=2��=�!�=L��=�=�Q=�(=��=�V�<��<�n�<���<�v�<�g�<��=��)=L�C=�Y=�fe=��b=�hI=<�= �3<�b߼�:����&��>��e Ѿn�@yF�9b}�v���r���Ϳn�߿č뿌��D��*�߿��̿�F���d���t|��EE�&{���̾�w��@z�Oσ���^�Ȁ!=]�=��=�߾=�   �   �o�=�=T~�=���=�|X=��'=P�<\u�<�Zv<8�@<�.><�Hl<t}�<�_�<L=j�8=�*[=0�u=�H�=Z�y=��Q=� =�M$�3_�sg�Cr�z¾�����H��섿槿:`˿
H�ʺ������xj�&��<�������쿆�ʿ4���'��.%G���ڮ���Xg�_��? ���~<`T=��=RB�=�   �   �z�=|��=}��=:�p=��;=*N=,��<��A< �;@V�:��:`�;�J8<8��<�[�<��!=v�H=V�g=��x=�Gs=�O=� =���LV�~��I�l�����)��'E�h���F��;ȿ�k�؋�,d�t�b��(��\�s�y鿅�ǿ>o��8ⁿ��C�Z��ӹ�'b���齪z����<�S=���=r+�=�   �   �X�= ߊ=� d=��&=���<�<�(���x��$�μ`����9���Ox��逻��<pٸ<�$=�(==��Y=��_=�/F=�{=���:��;�eh\�>~��N�:}:���w��Ӝ�@N��J7޿Gw���u�����N�������t��x޿�����\��P�v��&9����������R��mֽ�\���<��O=I��=\��=�   �   v=�C=P�< ~<��G�Bm	���W�Ä��I����ݩ�5����7���:{��[8���׼/�؋A<P��<S$=�E==s5=�=��;��lͽ^C�f��"�H�)��}b�揿�����̿9��'���m�|��l�����m翏�̿����˨��_�a���(�Ȣ�`3��0;�)a���¼\�<��H=G�=Z�=�   �   @=���<�\���ca��:Ž����7��P"���'���$��������ٽ�����N��V�� ��:���<2	="=�#�<��<<��Ƽ�У��#����YѾ"��2zG��~�����1W����Ϳ�u��f�r��I��5��5Nο	���d�����~�7-G���7�Ͼr(���d������c��4�<;=��[=��N=�   �   ��<�����.l���ɽ0��bA;��a��������Ս�k$��XD��@9h��D�.T��s⽉f���'���Ļ0�~<���<���<�'�<��>�vl��� ��_�蚭�l�����(��	Y�Q6��{̜�����v����C̿��Ͽ��̿5@¿
��A��#����oY���(��C���Ӭ���\��l��6�S��=r�P"�<*$=8�&=��<�   �   �r���铽w���l�7��t��ۗ�zf���Ǿ�Pվqbھ"N־��ɾO��~���vq}�4�A����̽���
(�x���[<H��<���< ��9(F�[�����*�������Ǿ���`�1��h[��Ё�����)z��9l�����;����d���_��d\��L2��v	���ȾM∾�-*�ô���`g�;H��<>z= ʾ<�P;�   �   ��|�
�+(Q��������}ᾦw��������G�{h�������#H������⓾��Y���r?������,����k<$s�<`�2<��f�dMf��]���I��ؗ���ӾD�
�E-��2N���k�8U��wň��j�����lȁ�x�l�&vO��T.����<�վW�����L����i�-[�x0X<@[�<p2�<@��:\D���   �   s9��W�Vr���@ξ8%��e�H�3��JF��<R�j�V���R��,G���4�������XѾ����`]�6��[��,� ;x=�<��<�/�;h�ϼ�����4���W�[n��<ξX"�Mb���3�GF��8R��~V�:�R�)G���4�Y�����4UѾ�|���\]�V���	�����5;�:�<X��<���;�м�����   �   ^�I�Kܗ��Ӿ�
��-��6N���k�RW���ǈ��l�����Rʁ��l�yO��V.����N�վ����،L���i��4[��2X<Ta�<�=�<��:0,��͝��2|
�x!Q��܏�<����ᾔt�]�����qD�<e����8��uC�����ߓ�*�Y�3���:��T�������k<(o�<��2<��f��Xf��e��   �   ������Ǿr��X�1�Pl[�pҁ�����[|��un��5���V�����#��a���f\��N2�Sx	���Ⱦ�㈾0*��Ŵ��Ph�;���<�~=Xؾ< �;(X������������7�4xt�ח��a����Ǿ�Jվ�\ھ�H־��ɾ�J������k}��A��������(��k���[<ܼ�<4��< �9�N�������*��   �   ���u�����(��Y�8��jΜ����������E̿��Ͽ��̿B¿����B��V����qY�B�(�F��0լ���\�
o��`�S� ?r��%�<�-$=�&=��<0�<d����l���ɽ��j:;�`|a�e������э�Q ���@��d2h��D�<O��k�l`�����|Ļh�~<8��<���<d!�< �>�Dl�Ԏ ���_��   �   *\Ѿ���|G�Ȼ~�C���Y����Ϳ�w��h�n��&����࿯OοL���m�����~�|.G���x�Ͼ@)���e�������c��7�<;=z\=H�N=�=Ԗ�<���b��DX���/ŽU���"��"�T�'��$�q�����ٽ����F�N��D�� m�:���<z	=z"=� �<@�<<��Ƽ!գ�N�#�`����   �   �$��)��b�Z珿K��W�̿������xn�T��2��^����翇�̿d���e���F�a�z�(�����3���0;�wa��`¼`��<.�H=�=��=�v=JC=#�<��<8�G��^	���W�M|�������ԩ��z��+0���,{�fO8�H�׼���ФA<0��<�U$=�F==�r5=�=P��;���ͽaC�!h���   �   ���~:���w��Ԝ�iO���8޿�x��Pv�d��$O�$��X���u��޿����2]����v�+'9���������R�$mֽB[�\��<��O=���=��=�Z�=��=�&d=��&=h��<h�<�׸��c��@�μ�x��p��%���-x�@���`�<<�<X(=f+==,�Y=8�_=�.F=�y=�l�:6�;�@�Ck\�����   �   �*��(E������	ȿwl�D���d������l�"]�0s��鿑�ǿ7o��'ⁿ��C��Y�Fӹ�lb�t��lx����<�S=���=�,�=�{�=���=<��=�p=L<=�R=` �<��A<��;���: ��: ;�;8Z8<���<a�<��!=��H=�g=��x=BGs=�O=�� =@p���V���g�l�I���   �   7��7�H��섿}槿�`˿cH��� �����xj��� ��|��-��&�ʿ�3��7'���$G��󭽾aWg�6��; �p�~<FT=^�=�B�=Tp�=��=�~�=���=D}X=$�'=0�<�u�<[v<��@<X-><�Fl<0|�<,^�<8K=x�8=�)[=�u=XH�=
�y=��Q=�  =�v$�x6_��h��r�h¾�   �   �)��'E�z���K��-ȿ|k鿶���c�.�
�����\��r��鿹�ǿ�n���ၿ��C�Y�Bҹ�b�����u� ��<�S=)��=�,�=|�="��=T��=T�p=r<= S=� �<��A<P�;��:@��:�=�;�[8<���<b�<�!=R�H=��g=��x=&Hs=�O=|� = 1�� 
V�	����l�C���   �   ,��|:�P�w�Ӝ��M���6޿v��(u�*���M����2���s��3޿]����[���v�f%9�R��"����R�eiֽ2V�4��<�O=v��=���=[�=��=b'd=.�&=��<��<pո��b����μ�w��o輰$���*x����� �<P�<p)=�,==��Y=��_=1F=�|=���:��;�ih\� ~���   �   =!��)��|b�s叿��ò̿���}���l�������8����
���̿$���}���(�a��(���01���,;�J\��L¼���<\�H='�=v�=�v=C=($�<x�<��G�L^	�x�W�|��X����ԩ��z���/���+{�PN8�̥׼ ���A<���<�W$=fI==�u5=�=�;( �qͽN]C�re���   �   �WѾ/���xG�6�~������U��y�Ϳ�s��d�n��6��(��8Lο1��������~��*G����Ͼ&��a�s��� �c�lC�<�;=\=��N=�=���<������	X���/Ž������"�'�'���$�3�����s�ٽڪ����N��@�� ��:H��<f	=&= *�<�<<��Ƽ�Σ���#�.����   �   H���)���t�(��Y�5��˜�䇱������A̿��Ͽc�̿�=¿���?��]����lY�2�(��?��sЬ���\�Te����S���q�|2�<2$=Ə&=��<8�<�����l�`�ɽ���L:;�C|a�V��|��pэ�5 ��d@��2h�nD��N��j�e_�����gĻ8�~<$��<��<l/�<�r>�Lql�� ���_��   �   ˥��`�Ǿ_��L�1�Lf[��΁�䊓�2x��j��ƕ������\�A���]��~`\��I2�;t	���Ⱦ,߈�+)*�ͻ��l�����;���<$�=޾<  ;�U������C�����7�xt��֗�ra����Ǿ�Jվ�\ھ�H־��ɾyJ��y����j}���A�B��ض����'��^���[<�Ǽ<���< �9�@�����	�*��   �   `�I�Q֗�g�Ӿ;�
��-��/N�"�k�NS��gÈ��h��x��FƁ�c�l�erO�.Q.������վ����܃L��	��i�@ [�hWX<�m�<F�<�i�:�(��7����{
�Q!Q��܏�/����ᾎt�W�����fD�.e�x��#��CC�ޥ��lߓ���Y����69��2���󯻸l<4}�<��2< �f��Ef�}X��   �   X1�(~W�jk��N8ξ ��_���3��CF�15R��zV�;�R�6%G�*�4�������&PѾ�x���U]���u���켠�;0N�<T��<N�;��ϼෑ�h4�t�W�Kn��<ξR"�Hb���3�GF��8R�w~V�+�R�)G���4�A������TѾ�|���[]����.���	� �; H�<p��<_�;��ϼ�����   �   ����Dx
�VQ�^ُ�8�%��q�O��Q��A��a�/�����=����`ۓ��Y����u1����`����l<���<0�2<ȶf�PKf��\ｲ�I��ؗ���Ӿ@�
�A-��2N���k�5U��tň��j�����dȁ�d�l�vO�iT.�x���վ���(�L�D�i�0[��GX<\k�<�H�<��:l���   �   �C��Uړ�	���e�7��qt�ӗ��\����Ǿ�EվSWھ1C־B{ɾ~E�������b}��A��������\�'�:��\<4ϼ<���< ��9�C�����R�*�|�����Ǿ���^�1��h[�Ё�����'z��7l������4����Y��}_���c\��L2��v	�u�Ⱦ∾l-*�����H����;��<Ѓ=T�< l ;�   �   0�<䌮��l��ɽ���:4;�Lua����Z���(͍����C<��b*h��D��H��`�-W�����Ļ0�~<�<��<�1�<�u>�tl�6� �ƹ_�ܚ��f�����(��	Y�P6��{̜�����s����C̿��Ͽ��̿+@¿
��A������oY���(��C��zӬ��\��k��V�S���q��-�<�1$=�&=��<�   �   �=d��<��V��iP��|&Žů��L���"���'�n�$������3�ٽ졡�~�N�(�� �:dɩ<�	=�)=�.�< �<<��Ƽ�ϣ���#����YѾ��3zG��~�����2W����Ϳ�u࿽f�k��B��,��+Nο ���Y����~�%-G����ϾG(��Bd�������c��=�<,;=L\=*�N=�   �   f�v=2#C=2�<��<��G��Q	��W�$t��٠���˩��q��C'���{��?8���׼��໨�A<��<n]$=�M==�x5=�=��;����ͽ�]C��e��"�H�)��}b�揿�����̿7��$���m�x��h������d翅�̿����è��P�a���(����?3���/;�``���¼���<�H=W�=l�=�   �   \�=m�=�+d=�'=X��<�<0���O��<�μ�a�Y���0x��]���<|�<j/=�1==��Y=�_=f3F=l~=��:��;��|h\�9~��N�:}:���w��Ӝ�AN��J7޿Ew���u�����N����ހ��t��p޿�����\��E�v��&9�~��袮���R�mֽ[���<��O=N��=��=�   �   P|�=���=*��=��p=N<=�V=��<8�A<�F�; ��:�q�:@i�;Hp8<8��<�j�<��!=��H=��g=��x=VJs=�O=T� =@��V�j��=�l�����)��'E�h���E��;ȿ�k�ڋ�,d�t�`��&��\�s�u鿁�ǿ:o��4ⁿ��C��Y��ӹ�b�u���y����<�S=���=�,�=�   �   ��=�&�=j��=x�P=t=���<�4<@ӈ:�H��89�� ���U� E�;�9t<���<�#=��L=�3o=�=��r=�@=<Z�<�'�����oz9�����߁��R�8�p�~��ݦ��5ѿU�����D&�6�>�@�:RD�Β@� �5��&�����r��86п�֥�҉|���6�o���`���0�㚽�=��=��y=���=�   �   �ٖ=���=�l=Ա3=o�<H�a< �9x ,�P����﫼����Tq���Ļ01�;���<6�=0�5=�w]=�r=ʌj=<=�ӱ<���p�����4�x���Ԋ���5�z�z	��[�Ϳ�9��d��8s#�b�2�<#=�R�@�v$=�`�2��L#�,j��s����̿���J)x�>3�͵�s��<�+������4�v8=�t=�Ӓ=�   �   �\�=��]=Z#=�<��C;<<������<�doa��p�X�i��+M����¼��ۻH�1<D��<6'=<zJ=P�P=�.=�ɱ<��'W���(�h����#龯-+�x�l��Λ�4�ÿ�Q�(�	�`�x�)��Q3�ֵ6�Tc3���)�B_�ʕ	�/�뿷ÿ���	jk�X�)���P᏾������?���
=b:d=�$�=�   �   T�8=���<Ht<��4+�� ���鸽�W޽E���a �i���j�NĽ���O�<1Լ "���<��=F#=%=h�<@�6�v�����.����ҾD��T�X��玿�����ٿ����~��2�$��'��$�<4�j1�����i�ٿ�³��q���gW��i���Ͼ������ �e� �Ⱥܮ=�4G=.mU=�   �   D�<P~����� ���ݽ���
&5�P�O�i�`��eg��b�� S�d:�F��UZ�z٤�z=������ <��<��<�M�<�����MO��A��בa��^��$���t>���|���a¿��^@������p(�ޮ�4X��������]O¿��{|��=��'�#U����\��L���2���;
�<��=Xy
=�   �   ���tZ��FȽ�j��0M��؀�4`�����Q���ϻ��/���Ѭ��՚������T�&����ٽ$�~��ռ 8�8�1j< Pp< s��:(�`d���V6�$������K� ��RW����1����ÿ5�ܿnx�eD��R� ������%�rݿ�CĿj����_��>uW�� ���⾜b����2�䤶�$����y�;��<�~�<�|<�   �   �����p코M6���}������)ɾ���8��{
�[����
�r��5c�̾�ԧ�Z���֚=�!+��B'���K���O��@K�;�`�:����(��H
���k�gյ�@L��0���a�J���P����k��Fɿ�Կ ؿ߂Կ��ɿ57��⸣�-����b�[�0����ᵾ4k�ry�����,<���8�;psK<@R;h����   �   Ga���E�����.e��e^�~���(�<�9���D��	I�wE���:��^)�p�p��w¾H����;K�(��L����輀��� ��:��%�`)������,�������Ⱦ��	�o2���\����I^���e��sl��Υ���ë����_��}I��V�]�]�3��{
��Gʾn��[�-����y&���0Ԉ;@Ī�,�Ƽΐ���   �   �*B�{]��ci̾4[� �'��H�$�d��a{����������D���q|��"f��I�:)�ӱ���ξjj����E��Ko��	��@�ߺ@�������Nf�J5��$B��Y��sd̾0X���'��H���d�]{�0�������JB���m|�f���I�B7)�����ξ�g��اE�4�콞Eo������ߺ ����
��v�f��=��   �   ���j ɾh�	��r2�}�\�M����`���h��o��d���)ƫ�D��s!��NK��f�]�ז3��}
��Jʾp���-�'���|&� ���;�𩺨�Ƽ~���XW��|�E�|���`��^X����(�0�9���D��I�sE�B�:�a[)�m�(k��%s¾=���>7K� ��H������������:P�%��%)����{�,��   �   ٵ��N��0�R�a�c�������hn���Hɿ�"Կ�ؿn�Կ7�ɿS9������/��P�b�M�0���㵾�k�{�;���L<���M�;��K<@�;����ޡ��,f��F6�x�}�с��$ɾ�����(x
���c�
�`���]�I̾�Ч�#���ޕ=��#��#"���>��`6�� L�;��:h(���-��  
���k��   �   ����� ��UW����L��N�ÿ��ܿ{�G���� �5���(�tݿ~EĿޏ���`��wW�x� �����c��v�2�O���Ą��`��;(�<0��<Т<@ncZ�n<Ƚhd�)M�TԀ�j[������K��Aʻ��*���̬�uњ���cyT���0�ٽ��~�4�ռ Ԓ8p9j<�Lp< 瑺$/��i���Z6������   �   ��Aw>���|����_¿���B�������)���@Y�����r�⿞P¿���||�5�=��(�(V��ڡ\�N�
�2�`�;�<0�=Ȁ
=!�<���>��@����ݽ����5�O���`��]g���b��S��]:����Q�Ҥ��=�����
<�Ž<��<�J�<P���TO�TG����a�la���   �   ����X�鎿O��w�ٿ������ �R�$��'��$�5�$2�����X�ٿIó�_r���hW�xj���Ͼ��ƭ���e�@�Ⱥ±=�8G=�rU=��8=8�<8�<��X$+�����฽<M޽����R\ �������_EĽW똽D�O��Լ�����<��= 	#=�$=hݬ<(�6����|
�k0��7�Ҿ�   �   */+�R�l��ϛ�x�ÿGS��	��`�X�)��R3���6�d3�r�)��_�(�	����ÿ���Xjk���)����G᏾r��d��p0��0
=�=d=�&�=_�=�]=�#=��<`TD;p%���{�~�<��aa���p���i��M��H�����ۻ�1<���<V9'=.|J=�P=<�.=Xű<����YZ��(�����%��   �   �5�nz�G
��@�Ϳ�:�����s#���2��#=���@��$=���2�M#�@j��s����̿���)x��=3�P��r��|�+�0���+��:=Z�t=2Ւ=ۖ=���=l=��3=�y�<P�a< �9��+�X����⫼����>q�p_Ļ�Q�;\��<��=��5=�x]=(r=X�j=� <=�α<�%�����v�4�ǌ�������   �   �8�A�~�ަ�Q6ѿ�U�����D&�46�R�@�:RD���@���5�p&����r���5п֥��|���6�Q��������0�ᚽ@2��=��y=j��=x�=
'�=���=f�P=H =��<�4<�݈:�G���9�P� �`�U��?�;06t<���<�"=~�L=�2o=> =.�r=@=�U�<�-������{9���������   �    5�Lz��	��c�Ϳ{9��L��s#��2��"=���@��#=���2�jL#��i��r����̿���'x��<3����q��J�+������"�.<=@�t=�Ւ=Hۖ=���=Fl=��3=�y�<��a< �90�+������⫼����=q� ]Ļ`T�;��<$�=d�5=fy]=�r=(�j=�<= ұ<L!��w���>�4�勝�R����   �   �-+�+�l��Λ���ÿPQ�ȴ	��_���)�6Q3� �6�pb3���)�h^��	����uÿw��3hk�ލ)���徜ߏ�*��W���@���
=d?d=L'�=y_�=��]=<#=H�< YD;%��Z{�D�<��aa�X�p� �i�PM��������ۻP�1<|��<d:'=~}J=��P=l�.=T˱<4�3W���(�`���w#��   �   �����X�/玿����ٿ������" �.�$��'��$�3�X0�������ٿ����|p���eW�5h�A�Ͼ������,�e��Ⱥ~�=0;G=rtU=��8=��<��<����#+�~����߸�M޽P���5\ �����o��EĽ�꘽J�O�xԼ������<X�=j#=
(=��< �6����F�.���Ҿ�   �   S���s>�B�|���¿]�⿉>�����~�.'�����V��������ZM¿Z��x|���=��%�<R��Z�\��F��2�@i;��<,�=��
=�#�<����������ݽ����5���O���`��]g�c�b�jS��]:�����P�^Ѥ�p=����� <�ʽ<�"�<�T�<Pۼ�6JO��?��Y�a�~]���   �   ����� ��PW�������8�ÿ+�ܿ"v��A���� �����#�pݿ`AĿF����]��rW��� ���⾢_����2�%����n���Į;�<���<@�<x싼zbZ�<ȽHd��(M�IԀ�_[��}���K��.ʻ��*���̬�Uњ���yT��Z�ٽ��~��ռ Ԙ88Ij<(cp< 됺�#��a���T6������   �   ;ӵ��J��0�'�a�����y����i���CɿIԿa�׿$�Կ)�ɿ�4�����\+���b�E�0�(��2ݵ�hk�u����%�����;�K<`;P���/����e콾F6�[�}�Á��$ɾ�����"x
���W�
�R���]�"̾�Ч�񁂾p�=��"��� ���8�����Py�;��:$��x%��
�}�k��   �   �����Ⱦ��	��l2�u�\�A���4\���c���i��5������_������7G��J�]��3��x
�@Cʾwj����-�����l&����`)�;�V��t�Ƽ�����V��J�E�i���`��TX�	���(�-�9���D��I�sE�4�:�P[)�m��j���r¾����6K�o�PG�����ș����:x�%��)�����m�,��   �   � B��V���`̾�U���'�\H�ݺd��X{�����4����?���h|��f���I��3)�s���ξ�c����E�y��h6o��쨼�Q޺�(��@򝼎|f�o4罔$B��Y��hd̾,X���'��H���d�]{�.�������EB���m|�f���I�-7)�v����ξ�g��V�E����
Bo�������޺�=��,흼�vf�c/��   �   (P����E�R���\��kS����(�q�9���D��I��nE�%�:��W)��i��d���m¾쌑�V0K��� �B@�����P�����:��%��)�ꢿ�/�,�������Ⱦ��	�~o2���\����H^���e��rl��˥���ë����V��sI��A�]�I�3��{
��Gʾ�m����-�|���u&������;�"����Ƽ1����   �   ƛ��^콦A6���}��}��6ɾ������t
�x����
� ��UW쾇̾�˧��}��Ԏ=�i�����!���։�`��;�J�:@��1'���
�M�k�Uյ�;L��0���a�K���Q����k��Fɿ�Կ ؿۂԿ��ɿ+7��׸��u-����b�F�0�����ൾ�k��x�����h1��w�;��K<`I;,����   �   �ۋ�xVZ�4Ƚ&_��"M��Ѐ�W������F���Ļ�h%���Ǭ��̚�z탾�qT�r���ٽ��~��fռ  �8hbj<`rp< ���`$�3c��hV6�������J� ��RW����2����ÿ8�ܿnx�dD��P� ������%�rݿ�CĿ_����_��,uW�
� ����mb��r�2�d����{��@��;��<���<��<�   �    0�<@ʮ����W��=�ݽ����5���O���`��Ug���b��S�vV:�%��gE��Ǥ��=���� 9<ٽ<�,�<�Z�<�м��JO��@����a��^��"���t>���|���c¿��_@������n(�ڮ�0X��������TO¿��{|��=��'��T��E�\��K꽞�2��0;�<��=��
=�   �   ��8=4�<@�<�]��+��׸�DC޽�����V ��������3;Ľ☽��O���Ӽ`��x��<H�=�#=�+=��<X�6�s����p.����ҾC��T�X��玿�����ٿ����~��.�$��'�
�$�64�d1�����_�ٿ�³��q���gW��i���Ͼ���%����e���Ⱥ�=�;G=�vU=�   �   �`�=P�]=T#=`#�< �D;���Pp��<��Ta�ʪp���i�M�"�D���9ۻ(�1<<��<v@'=T�J=n�P=t�.=б<x탼�V��~(�\����#龰-+�z�l��Λ�5�ÿ�Q�*�	�`�x�)��Q3�Ե6�Pc3���)�<_�ƕ	�)�뿱ÿ���jk�P�)�ͺ�8᏾l��Y��p-���
= ?d=�'�=�   �   �ۖ=J��=Rl=��3=��<@�a< ��9h�+�����xի�(���`#q��*Ļp��;���<��=z�5=�|]=�r=Ώj=><=�ֱ<p��&���{�4�q���ъ���5�z�|	��\�Ϳ�9��d��8s#�b�2�<#=�P�@�t$=�^�2��L#�(j��s����̿���F)x��=3�ŵ�s���+�+����/�:=&�t=dՒ=�   �   8�=D�=�T=�=4.�< ��;D�����@�ڼ���*�T��� ~J� ��9�	t<�b�<`�0=VGZ=��l=d(^=<� =�)<"+�U���9p�S_ʾ"0���a��G����ȿO����A��11���I���^��m�t7r�m��^���I���0����Il���ǿ���3�_��*�}�ƾ^�h���彪����<eG=�Ղ=�   �   ��=��j=��8= ��<��B<�V��T��n����'��q5��.����,8̼�1�`T�;�6�<0�=E=�]]=p�S=�=@�<4g%�Ӊｬ�j��Bƾ�7���]�ß���ſͬ�����!.�8!F�"Z�Tch�TZm�&eh��oZ�<�E�<�-�6��u��hGĿ�y���[�eG�ڋ¾�hc���߽ �� |�<�tA=P�z=�   �   �kR=��'=�&�<�pw; ����W$���s�϶��㑮�����b���J���V���Dh:���˼ �o�p�<
=�-=�)4=�K=@�<̢���ݽ�s[�O[��h��U�Q��揿λ����(��$b%�ԩ;��dN��[���_�N5[�$�N�֩;��6%�44����8ݺ������P���������T��Ͻ��켤2�<6�.=\�X=�   �   
�<�IQ<�@�(G&����pϽk3���a'���,���(�(��bV�&�ٽ,���̳B�@���Z�;�<�}�<P��<`�;<��^T½r�C�姾�+�^?�H̓������DؿZd�����+��s<���G�j�K��G�R�<�6:,��-��R�g�׿�
��&��	>�������:�=��g����żpGw<,�=,&=�   �    �ܹ\%�1���@ڽd�=�E��.m��;���k���.��B*��}����Dq���J�t���Z���������R(<��{<@%�;�ͼPF��2&�s����e例�'��h� 4��n���]��"��8��R'�
[0���3�ʟ0�0p'�,_���.�î������h�� '�f⾾��4T!��w��P0��8A7<�<|q�<�   �   ��-�d����e��rJ��K��X���޴���
׾g�徜�꾺X�9�ؾ��¾N/��L%��t�P�ȥ��N��\�F�l���@��� �w�࿣�Ϋ|�Ǽ���m��[���h���E�����¥�K�ȿ�w���Z��&������	�<u�����a��ɿ��:(���E�'��Z%���j�
*��l�أ{� 4�;���;p @��   �   �jƽ@�"�ao�ؕ���Ͼ*W��TA�s� �\�*�z.��Q+���!�m�s��'aҾ�q���t�&(�d�н��^����� �-�pҌ�z�:��Rʽx9�d;����㾆&!�7�W�~\��r���Ŀ�Oݿ�4����^�S���" �Ea޿�ſ�;���䉿d:X�d!���㾱ʖ���7��ƽ��/�8	d�p�޻ ���j�K��   �   R	)�#���?A��M�ﾗZ�0�3��;N��c�pp�{@u�rq�Kd�ÚO�;n5�x����P����炾B�,��ν�LX��[̼P������,���2���Ac�=�����)��Z�s,���������|wÿ}οE�ѿ�ο�CĿ��<���������[���*��4��������c�\��,c��\����%��4��@�L�~�ǽ�   �   �}�(���\C���&���M�l)t�����X��UM��1K��k ���֋�F�u�nO�j'�� ��[��p��
!�+P���5��������2��_������
}�����v=��9&���M��$t����;V���렿���H������Yԋ�J�u��jO�Fg'�� ��X������ ��L��x�5�����&���2�g������   �   E�=��L�)��Z��.��C������{zÿ�οO�ѿ�ο<FĿR���_���� ����[��*�8��������c�D���d��̀������B�L���ǽk)�?���J<��9���V��3�L7N�c�#kp��;u���p��d���O��j5�����z򾤵��傾n�,��ν,GX��X̼����������N��hGc��   �   ���h)!�ͣW��^���t��?Ŀ�Rݿ8�����`�[����"��c޿�ſm=��i承�<X��e!�;��U̖���7��ƽږ/���c��l޻|蝼l�K�Iaƽ��"�Yo�񐢾;�ϾzP���=�� �E�*��u.��M+��!��i����R\Ҿ�m����t��!(�*�н��^�������-��،���:��Xʽ9��>���   �   k���E����ť���ȿwz�R�������0��b��v�ؤ��c�Бɿu��P)����E�N���&����j��*�
l�@�{��Z�;�=�; �?���-������_�OkJ�<G��+�������׾��;�꾏R�y�ؾ��¾�*���!��_|P����G����F�pt��@S����w�ȣ�г|�����m�_���   �   ��'���h��5��~������t������'��\0�N�3�D�0�|q'�H`��������k���fh��'�Og�y����T!��w���,���P7<$��<���< (׹�����}5ڽ� ���E�]&m�
7���f��*���%��C���;=q�X�J�����Q�������P���pb(<��{<0�;�ͼ|J��L5&�ݵ���h��   �   (`?��΃�7����Fؿfe�(�6�+�&u<�6�G�ډK�`�G�n�<� ;,�l.�@S�D�׿]���&���>���M����=�zg���ż8Tw<��=�,=�<htQ<��?�R7&�����
fϽ�-���^['�n�,�r�(�`��#Q��ٽ����n�B�������;h�<x��<���<P�;���tX½��C�X秾H-��   �   �Q��珿bϻ�����c%��;��eN�
[�ȭ_�H6[��N�r�;�$7%��4�#�鿅ݺ������P����������T��ϽT��@8�<��.= �X=�qR=��'=�7�<�x;���dJ$���s����܉����������)���郂� ]:��˼�eo���<=��-=�*4=�J=��<|��D�ݽ�v[�K]��Ú��   �   �]�����܀ſۭ�����~".��!F��Z�dh��Zm��eh��oZ�t�E�V�-�6��u��PGĿ�y����[�G�V�¾�gc��߽R��D��<�wA=d�z=��=��j=��8=��<��B<� ������ȸ���'�j5�z.�H���,̼H�1�pt�;�<�<Z�=VE=^]=
�S=��=��<dk%������j�&Dƾ�8��   �   ��a�H���ȿ�����A�D21���I�"�^��m�t7r��m��^�x�I�@�0�t���k����ǿi��c�_��)�t�ƾΌh�j��V����<gG=�ւ=�8�=�D�=��T=�= 0�<P��;�A�Ƚ����ڼ���h+缈��� �J� 
�9�t<<`�<�0=�EZ=F�l=�&^=,� =<�+������:p�c`ʾ�0��   �   ��]�埗��ſԬ�����!.�� F��~Z��bh��Ym�rdh��nZ���E���-�t5��t��}FĿ'y����[�]F�K�¾`fc�/�߽���l��<�xA=�z=��=��j=��8=(�<8�B<���x��������'��i5�P.���,̼H�1��v�;�=�<Ə=�E=�^]=��S=ܽ=��<�h%���|�j�Cƾ8��   �   $�Q��揿�ͻ�$��ԇ��a%�2�;��cN��[���_� 4[��~N�¨;��5%�\3�7���ۺ�y���P�l��������T�I�ν�z케>�<��.=D�X=�rR=z�'=�8�<�x;����:J$���s�箙����������������������\:�̴˼ [o�x�<=¬-=R,4=M=��<�����ݽ�s[�G[��V���   �   q]?��̃�����Dؿ�c�<���+��r<�j�G���K���G��<��8,��,��Q���׿*	���$����=�
�����ʸ=�~b��ثż�ew<��=j.=L�<�wQ<��?��6&������eϽ�-���L['�V�,�V�(�<���P���ٽ#�����B����P��;��<��<(��<0-�;T��bS½ʸC��䧾M+��   �   ��'���h�53��=���ݳ�6����'��Y0�$�3�,�0��n'��]�����鿳�������,h�K�&��b�4}��nP!��q�����e7<���<膎< ֹ 뼛��E5ڽ� ���E�N&m�7���f��*���%��1���=q�#�J����pQ�8�� ������0m(<�{<PE�;�ͼoD���0&�����Fd��   �   �g���E����������ȿ�u꿞���������6��s����^뿛�ɿ���d&���E�����!��Ϳj�"&�$�k�y{����;�Z�;��?�0�-�$���l_�1kJ�1G��!������z׾���,��}R�b�ؾz�¾�*��e!��|P�����F��z�F��n���͉� cv�H�����|�(����m�	Z���   �   ��㾿$!�ݝW� [��Ep��XĿ4Mݿ/2���W]������A^޿�ſ9���≿�6X�a!�:��Fǖ���7��ŽΉ/�8�c��>޻,᝼�K��`ƽ��"��Xo�␢�1�ϾsP���=�z� �@�*��u.��M+�ݦ!��i����-\Ҿum����t� !(�
�н��^�����-��ƌ�b�:��Nʽ�9��9���   �   �뮾j	����)�}Z��*������W����tÿ�ο;�ѿ�ο}@Ŀ�ﳿ��^�����[�P�*�>/��]���X�c�����[���g��x��踼ҀL���ǽ)�$���9<��/���V��3�L7N�c� kp��;u���p��d���O��j5�v���z�v����䂾��,�~�ν$CX��L̼d����5�������=c��   �   �}�?���#9��y&�K�M�� t������S���蠿�����E������ы�o�u�lfO��c'�� ��S�����l� �D��<�5��p������ 2�m^����k
}�r���k=��6&���M��$t����<V���렿}���{H������Sԋ�:�u��jO�3g'�׳ �dX�����u� ��J���5��y�������1��Z��	���   �   -�(�b����8��l��
T���3�K3N���b�`fp��6u���p��
d�*�O��f5�����t򾃰��Ⴞ�,��ν�7X�P>̼d鐼���������$Ac�!�����)��Z�t,���������}wÿ~οD�ѿ�ο�CĿ��3���������[���*��4��[���&�c�����`��hs�� ��<丼�zL���ǽ�   �   %Zƽ6�"��Ro�����Y{Ͼ�J��K:��� �N�*��q.��I+��!�f�����SVҾ�h����t��(��{н8�^�<����u-�������:��Pʽ�9�@;����㾃&!�6�W�\��r���Ŀ�Oݿ�4����^�P��� �>a޿�ſ�;���䉿T:X��c!����vʖ��7��ƽ��/�`�c��8޻T؝���K��   �   ,v-������Z�eJ�hC�����������־�~����L�4�ؾ��¾|%�����ytP���� =���tF��X���߈��=u�x���n�|���p�m��[���h���E�����¥�M�ȿ�w���\��$������	�8u����|a��ɿ
��3(���E���,%����j�B)��l���{�Ѕ�;�r�;��?��   �    �ҹ���~��$,ڽ����E��m��2��bb��R%��� �������4q�~�J����)F��
��\��@t����(<h|<pb�;�ͼ�D���1&�R����e例�'� �h�!4��q���_��$��:��R'�
[0���3�ȟ0�,p'�(_���&鿼���|���h�� '��e⾎���S!��u��d%���`7<(�<쏎<�   �   H'�<�Q<��?�6*&��𑽭\Ͻ?(���U'�ۿ,���(����!K��ٽ�y����B��蝼��;H��<���<@�<�E�;����4S½�C��䧾�+�^?�J̓������Dؿ\d�����+��s<���G�h�K��G�L�<�2:,��-��R�d�׿�
��&�� >�������һ=�kf��̴ż@^w<6�=01=�   �   FuR=��'=�D�<��x;�~���>$���s����� �������z~�����T|��$O:��˼��n��$�<2#=��-=�04=�P=��<r��גݽ�s[�D[��h��V�Q��揿λ����*��$b%�ԩ;��dN��[���_�L5[��N�ҩ;��6%�24����4ݺ������P����������T��Ͻ���:�<~�.=|�X=�   �   H�=|�j=R�8=�
�<�C<����|証���f�'�,b5�h.�:��D̼�i1����;�H�<��=�E=>b]=��S=��=h�<f%�}�ｕ�j��Bƾ�7���]�ß���ſͬ�����!.�6!F�"Z�Rch�RZm�$eh��oZ�:�E�8�-�6��u��fGĿ�y����[�bG�ы¾�hc�1�߽�����<XwA=Ъz=�   �   ^�q=P`[=^G*=�I�<�:�;`� ��Ѽ|��BZ=�~yJ� �A���$�@T�`d� �9;8�<��=d@=��U=�TD=���<`��`��Ћ��A��é�i8�(��n���������/���O��9o�]E������u�������/����n�L,O��	/�FI���濷����XR6�j��Ύ�/����d�@[2;
=��`=�   �   �2_=��B=N�
=�҃< Ec� 0��n�#��[�ND��l_�������d�@�0�,�ۼ ��H�,<@v�<"(=�C=o8= ��<�D����y�o��\+�����R�4�:Ӂ��f����z����,�\�K��sj��u�������Ҏ�����k���,j��pK�`,�B���J����Э��9�2�;P�*Ћ��h��$_��a&;�{=NT=�   �   �'=(��<��'<(%T�x���:���A���ѽ�m�1E�/��Ùս|ȳ�Ā��&Q/�t:�����;d�<z�=r�=�;�<P���F�g�����F���#߾�+�&v�����ʢٿ���>$�&A�b]��#u��܂�6څ����pHu�8]���@�F�#�dG�C�ؿ߅��7&t��J)�m�۾�/��ϔ�*O����:h��<|W.=�   �   ��<�G@�d���P���ʽ���q'�i@�ƪP���V��Q���B�Q�*�$/���ӽ�挽 ��`���6<�˧<|��< f����N��2��.q���ɾʏ�C�`�}Ǚ�Jȿ!1����6�0�,;I��^�>Cl�Fpq�ʆl�|j^� �I�v�0���I���m�ǿ�
���l_��%�Ǿ��k��_��88� Ņ�Tn�<h]�<�   �   ࣒��M��û����HB�ڹt�W���3���"���,貾EP��c8������4�x��G�|��r^ƽN2c�� ����7��*=;��f"3��gؽ%O��������c�E��$���(��!"߿���2�1�zC�Z�N���R�O�.�C��Y2��s�p��I'߿�鱿.���Z�D���0߬�2�J�Y`ϽN* �@ȓ���<`�;�   �   .���X����3�4Tz�a1��,_ƾ��澲C �ל����| 	�� �G��P�ȾҤ��S���8�01��� ���j�?�� c��p7�����D�)��$��B�㾴l'��,h�2r��V��6����<'��b0���3��0��'�Ɩ�x ��Q�����R����g�y�&����䴏�ޜ&�˛���4��/H� �C������   �   �>�֗L�煒��"ľ?���T���+���=�SI�XxM��I�n�>��-�Z�������ƾQܔ�R�P�*�a���ܪ,�(��8��f���%b��pe��������0>��|�O���^¿������b������JZ����� ��9�-Hÿ����\}�Bk>�B��R:����c�q��]��<[��ɼ�������   �   N�S��霾_�پѪ���1���S�r��儿v����O��Q⌿�y��Lxs�xeU�vP3�=���۾�Ğ�t�V�^g�\�����4��J���V��Wý �+��A���@Ҿ�#�BJH�����{��.���׋Ͽ,_�Ɋ�����7Q��п㻸�Mf��
���q3I����l�Ҿo���]+� ½huR�{�u-�9>������   �   M��˾޾[����C�ڒq�ò��,���7��G ������@l��^���򢿿���>@s�TFE���GE��d���DI����y��TE)��w(��A��'l�<�G�I��n�޾���m�C��q����4��p4�����~���-i��~����w���`<s�/CE�{���A�<b���AI���x���F)�6}(� G��Pt�"�G��   �   EҾ�&�NH����~��*����Ͽ�b�K��B�� �QT��пS���]h������6I����A�Ҿ�p���_+�½4uR��v�vl-�l7��	����S��圾��پO����1��S���q�ㄿ����M���ߌ�,w���ss�qaU�M3�}����۾���� �V�xd�*����4�ZM���V��]ý��+�<E���   �   W���3>�)�|����{a¿��[���4�������\�~�h� �<�@Jÿ����m_}�Em>����<<���c�$r��]��X��ȼ�{��x��B9���L�L���ľ���Q��+�3�=�^NI��sM���I�/�>��-���^�����ƾ�ؔ�"�P�p&������,�������{����e�1ve�ɼ���   �   [o'�00h�F𘿄t��*��Γ����&'��d0���3���0���'�4���!��S�u��������g���&�s�������&�-���X2� H��C�|�������#w���3�rKz�.,��.YƾA��"@ �%���������� �D���Ⱦq����K�f�8�)������d��8��Dd���;������)�Q'��2���   �   ��E�X&���*��|$߿J������1�jC�`�N���R��O�̜C�4[2��t�L���(߿�걿󾇿p�D����
ା �J��`Ͻl( ������<�>;����B�M�`���l��AAB�	�t�t�������Ⲿ K��z3��;�����x�yG�B��\VƽX&c�L�`�7��D=;h���'3�ulؽ�(O�r�������   �   ��`��ș��Kȿ?3��N����0��<I��	^�$El� rq�z�l��k^�D�I�V�0����E���'�ǿ/��|m_�2&��Ǿ�k��_��68� ����x�<�k�<���< �?�d����G��A�ɽ�	��j'��a@�O�P���V���Q�θB�@�*��)��ӽ~ߌ��������6<�ѧ<H��<�x����N��7���1q�f�ɾ����   �   +v�����F�ٿd��B$�VA��]�.%u�N݂��څ�?��xIu��]��@���#��G���ؿ���o&t��J)�h�۾�/��_���O�@?�:x��<�\.='=P�<@%(<`�S����2��~9���ѽ�d�<�P�꽅�ս
���Sz��XF/��(��@͏;�!�<x�=��=$:�< Ē���g���� H��&߾:+��   �   �Ӂ��g�������H�,�,�K��tj�dv�����Hӎ�_���l���,j��pK�j,�<���J㿰��������2��O龧ϋ��g��!_� �&;�~=ZQT=�6_=L�B=��
= ߃<`�b�� ���#�X�[��?��[��𒂽J�d���0�̢ۼ ����,<8{�<�(=��C=�n8=��< \��`�y�9���,����쾇�4��   �   �(��o��Y��N��/���O��9o�E������t�������/��V�n��+O��	/��H���.��&򂿒Q6�6��͎�����d���2;@=j�`=ދq=�a[=�H*=L�<�B�;� ��Ѽ��Z=��yJ�x�A�N�$��U�Xd�`�9;�5�<r�=�b@=��U=SD=��<@w��R��+���B�����xj8��   �   gӁ��f����~����,�6�K�~sj��u��W���zҎ�����jk���+j��oK��,�����I�������	�2�nN��΋��f��_���&;�=RT=@7_=��B=ڽ
=�߃<��b�\ ����#�@�[��?�� [��ߒ���d�X�0�L�ۼ0���,<,|�<$(=F�C=�o8=���<�L��z�y����+����쾨�4��   �   �v�����r�ٿB���$��A��]��"u��ۂ�{م�����Fu��]�b�@�D�#��F�΅ؿ����9$t�I)��۾.��U��|O����: ��<^.='=x�<�&(<P�S�����2��d9���ѽnd��;�3��Z�ս���� z���E/��'���ҏ;�#�<��=J�=?�<P����g�����F���#߾�+��   �   ��`��ƙ�OIȿ!0��f��T�0�:I�L^��Al�jnq��l��h^�z�I��0����3�����ǿ0	��ij_��#�jǾ��k��Y�/8� ��� �<�o�<P��<�x?�P����G���ɽ�	��j'��a@�A�P�v�V���Q���B� �*��)���ӽߌ��������6<D֧<��<@P��X�N��1��T-q�2�ɾR���   �   G�E��#���'��� ߿�����1��C���N���R�O�>�C�X2�r����$߿�籿������D���Eܬ���J��YϽ� �0x����<�c;Ԇ��H�M����N��,AB���t�n�������Ⲿ�J��k3��(���T�x�DG�
���Uƽ�$c�P콼 g7�@�=;0��z3��eؽ�#O���������   �   Vk'��*h��옿wp��`��������'�a0���3���0�"�'� ����'O�k���;����g���&����豏�m�&�۔���(�� H� �C�p���֓���v뽟�3�SKz� ,��&Yƾ;��@ �!��ۛ������ �.����ȾS����K��8�S(�������`�0��$W��2�����j�)�;#��Z���   �   M���.>�^�|�����\¿@	�����~�8�>��hX��>� �i6�XEÿ�����X}��g>����g6����c��l�eV��bN�X�ȼ�w�nw���8�d�L�8���ľx��Q�|�+�1�=�[NI��sM���I�'�>��-����?���d�ƾ�ؔ���P��%�=�����,�����������`�ne�ﶶ��   �   �=Ҿ�!��GH�����y��á���Ͽ\�u��K��!��M�Ԩпݸ���c�������/I������Ҿdk��6X+�����gR�~m�pf-��5��t��.�S�h圾��پK����1��S���q�ㄿ����M���ߌ�(w���ss�caU�M3�m����۾z���}�V��c������4��C�,�V�VSý��+��?���   �   BF����޾w��E�C�,�q�ǭ��� ���1�� ���K}���e��T񱿃좿����z7s��>E���<��]��;I��u�p���8)�6o(�-?��{jｼ�G��H��[�޾��k�C��q����6��s4�����}���+i��{����q���R<s�CE�j��sA�b���@I��}�2u���=)�p(�t=��^f�>�G��   �   ��S�4✾J�پ���k�1��S�?�q�����튌�DJ���܌�gt��tns��\U��H3������۾������V��^�^���`�4��?�@�V�~UýL�+��A���@Ҿ�#�>JH�����{��2���ًϿ1_�ˊ�����3Q��пܻ��Ef�����a3I����;�Ҿ�n���\+�z ½�mR��o�8d-�+2��|���   �   ,5�$�L��}���ľ�	���M���+��=��II��nM���I���>�e
-���z�����ƾ	Ԕ���P�w �V���ؖ,�T�����U���2a�fpe�丶�����0>��|�P���^¿������d������JZ����� ��9�'Hÿ�����\}�3k>�0��:���c��o�TZ���Q���ȼ�r��r���   �   ���kn��3�<Dz��'���Sƾ6���< ����(��0��"� �����Ⱦ����B���8���k񏽐T� ���L���/������)�W$��*�㾰l'��,h�2r��Y��8����@'��b0���3��0��'�Ɩ�t ��Q�����K����g�l�&���⾢���
�&�>����,��H�X�C������   �   �u��vM�ذ�����:B�C�t� 뢾f���>ݲ��E��'.��@���y�x���F����*Kƽc��ҽ���6� �=;����3��eؽ�$O��������c�E��$���(��%"߿�� �4�1�|C�Z�N���R�O�,�C��Y2��s�n��D'߿�鱿+���P�D���߬���J�h^Ͻ`$ �@���H�<@�;�   �   �
�<��>�����R@��)�ɽ^��d'�[@��P���V�=�Q�r�B�^�*��#��{ӽ�Ռ�ޟ�8��H7<��<lÃ<�4��l�N��1���-q���ɾƏ�E�`�Ǚ�Jȿ%1����:�0�.;I��^�>Cl�Fpq�Ȇl�zj^��I�t�0�
��E���i�ǿ�
���l_��%��ǾJ�k�`^�48� ���D��<v�<�   �   *"'=x�<XB(<��S����D,���1��U�н�[轝2���R�սd���_r��08/�d���!�;�3�<$�=l�=G�<@�����g���jF���#߾�+�)v�����΢ٿ���>$�&A�b]��#u��܂�5څ����lHu�4]���@�B�#�dG�@�ؿޅ��2&t��J)�[�۾�/��`��vO�@^�:��<|_.=�   �   8_=d�B=��
=�<��b�����#���[��;���V��^���2�d��0���ۼ���,<��<�(=@�C=s8=д�<�4��Z�y�@��O+�����R�4�;Ӂ��f����z����,�\�K��sj��u�������Ҏ�����k���,j��pK�`,�@���J����Э��7�2�2P�Ћ�`h�b#_�@�&;�~=�QT=�   �   ZxU=�_==f�=t6�<`\x��/���U$��\�(3�����T���-c�>�.�LGּ�?��(�9<H��<�(=��?=��,=`��<X�{�;p��m]9�����؜	�kP�={���ȿ���V"��F�Txl������G��}���[�������L/���H����k�z5E�vw!�d� �{Fǿ9D���[N�����r���m3������!��J�<@�B=�   �   D^A=$:"=�)�<0L�;����:����e�j���߁��� ��X[���#��~%p���%� ����jz:�ף<x�=n,=�~=��<0 }������c5��1�����,�L��瑿�Zſ�[���fwB���g������ז�����������K̖�j���=g��A���������Ŀp���)�J�=�L����/�����p�$�\��<�F5=�   �   ��=��<�o����ۼ��^��㦽�rؽz���*���p�d��X��[�ݽ�v��In�T#��pd���m<,��<p��<��<t����;����)�%H�� �����A��i������󿂾��M8�N�Z�P�|��'���W��: ��k��x<��
�|�lfZ���7��1�	������5n����?��v��Tn���$�d����1��Ӯ<��=�   �   �l�;(���?�G᩽�:��`s#�$:F�U�a��s�fz���t���c�-�H�0�&��w �jJ����P� �����:��@<�$�;H��zG��X��|�����\0� ]}�(b����߿���)��1G�܊d�@�}�J�����ڇ�HY~���d��TG�*�(�vk�}߿���@�{���.�)�u������ƴ� �T���;<�Y�<�   �   L��8������+�j�d��T�����م��z�Ⱦ�1;>ɾT���z���$�� }h�RK/�U�(.�����8�f��� �X9���rt����r���Ⱦ����w_�Y阿cPǿ�#��JY�T0��rH�v]��;k��hp�ܜk�ܲ]�>
I��0����U%���ǿl~���~^���g�ƾw"n�w���qd�X���`�y��R#��   �   �ʮ�>r���T�(����⺾�=�­��� L���:��8��^��NJ�A������N�X��^�?G��jGL�й�s��W[��3۽��H�
���#�U�=�����x��[׿��0���_+���;���F��J��-G�g<�,�j�j8�R�׿&���n����=��n�2����E�6սζN� &ԼOҼ��=��   �   �_�t#p��n����ྦe�w�)��B���V�8Pc��g��c�/_W���C���*�t��㾆q��t�s�$�!�0�ƽ�jm�`�*��N�������n�����Ѿh���V�����h���GٿA��� ��\���$���'��$������i����1ڿx����l���!W��O�KѾ�ㄾn�Ж��XDE�`7!�$�b�;���   �   ��w���o���*"��KI�no��;���c��9۝��࠿=,��c����򈿺�p���J�_#�����'���Bcz��� ���ý #w��VR�=Ɏ�i��J�J��&��sx�FR)��0b�I����p���rͿ���n���25�����|�������X�ο�W��Ρ��3c��)�e��9���}J�egｱތ��M��`q�c�����   �   L��Vy���,��\]�����U;��Ŕ���\ƿ+ѿ�	տ&�ѿ�ǿ���&��4Έ���^��-��������k�.��!��(Vk���j�3?���&��kj����[s��,�(X]�K���R8�����Yƿ�'ѿտ��ѿ�ǿ8|��#$��̈��^��	-������벾&�k����T��bWk���j��D��h+�Xrj��   �   �}�U)��4b������s��vͿ���=���*7�����~�`�����
�οZ������&c�Q�)����!;���J��i｠ތ�|�M�ZWq��w�����e�w�������3&"��FI�4o� 9���`��؝�}ݠ�=)�������B�p�ѭJ� \#��������B^z�~� �R�ý� w�<YR�͎�4���J��*���   �   �j�o�V�!���k��Kٿ������p���$�Ʒ'��$����R��+���%4ڿW��)n���#W�VQ�oѾ>儾��&����@E��/!���b�D2���Y�lp��i��6���a�)�)�*�B��}V��Jc���g��c�uZW���C���*�Q���㾚m����s��!���ƽ6em���*��#N�����w��X���ƫѾ�   �   H�=�����dz��"׿�������a+���;�<�F�l�J��/G�i<��,����9��׿����v���% =��o�<3��,�E��սR�N�lԼ�;Ҽ�=�1���l���T�F����ܺ�7���� �H�Ϛ�>�������vD�X������.�X�JZ��@���?L�Ĳ�t��\[��8۽H�!���T��   �   ez_�+똿�Rǿ &���Z�$0��tH��]�X>k�kp��k�̴]��I�T�0�����&���ǿG���^����]�ƾd#n�Kw���od������2y�H(#����铋�X���+��yd�P��jz�����f|Ⱦt+;Zɾ֝������ ���uh�|E/�L�y'�������f�P� ��<��nxt����
#r���Ⱦ!���   �   �_}��c����߿4��
)�T3G�܌d�~�}�u���4��ۇ�[~�.�d��UG���(�l�L߿����
�{�F�.��)侬�����������T���;<�i�<���;�n��n�>�>ש��.���l#��2F�H�a���s��]z���t�	�c�f�H�I�&�s �gB���P�w�����:x�@<�(�;4��kJ����z�����^0��   �   �j��x�����~���N8���Z���|��(��~X�����k��=����|�gZ�@�7��1�k������Tn���?��v��1n����$����P�1�Xܮ<.�=��=h1�<@��4�ۼ��^�Zۦ�iiؽ������k�r������ݽQo���<n�����(��P�m<���<,��<h�<D���k>���)��I������H�A��   �   p葿\ſ]��x��:xB���g�;���/ؖ�����b��7����̖�3j���=g�"�A����v����ĿA���ɣJ��<������/�J�����$����<�J5=~bA=?"=`5�<Ё�;(������R�e������|�������V��R�� p�H�%�||�� n{:�ݣ<R�=:,=`~=�ޯ<�,}�t����e5�S3�������L��   �   �{��~�ȿ���|V"��F��xl�ɀ��H������\�������#/��|H��"�k�5E�w!�� ��Eǿ�C��[N�G���q��zl3�������!�xO�<2�B=�yU=Ba==��=�8�<�Jx��-���T$�R\�3��������2.c��.�tIּpI���9<|��<��(=�?=§,=p|�< �{�br���^9�������	�\lP��   �   �瑿([ſ\��ș�XwB���g�����Qז����k��H����˖�zi���<g�B�A���k����Ŀ����֢J�<������/�����І$����<`K5=�bA=p?"=�5�<p��;ܐ�����>�e������|�������V��;���p��%�|�� �{:lޣ<��=�,=J=h�<X$}������d5�f2��C����L��   �   �i��ޟ����6��:M8���Z�V�|�'���V��V���+j���;��^�|� eZ���7��0�l��i���m��C�?�8t��wl��T�$�,���H�1� �<��=��=�2�< ����ۼx�^�;ۦ�Niؽr�������k�d������ݽ$o��~<n�����#����m<@��<��<�#�<����s;����)�,H������t�A��   �   S\}��a���߿r���)��0G�v�d���}�@��������؇�W~���d��RG���(�Jj��߿g�����{���.�
&�K���r������nT�ȼ;<�m�<��;�l����>�ש��.���l#��2F�:�a���s��]z���t���c�H�H�(�&��r �B��8�P��t��@�:(�@<�E�;P	��OF��������澏[0��   �   Gv_�}蘿=Oǿ�!��PX�0�8qH��]��9k�:fp�h�k���]�(I�D�0�2���"��q
ǿ�|���{^����.�ƾ�n��o��fd�������x�H#�\��l����齬+��yd��O��ez�����`|Ⱦl+;Qɾȝ��u��� ���uh�GE/��K��&����� �f�H� ��/���nt����Or���Ⱦ���   �   ћ=������v���׿���փ�@^+���;���F���J�,+G��d<��,����6��~׿ى�������=��l��.���E��սةN��ԼT3ҼZ�=�Y����k�}�T�7����ܺ��6���� ��G�˚�8��x�����_D�?�������X��Y��?���<L�t��f�"R[��0۽��H�������   �   ^f�~�V�T��g���Eٿ������������$�~�'���$�Δ�Ģ�����.ڿ����hj���W��L��Ѿ���������j6E�)!���b��0��`Y�,p��i��'���a�&�)�(�B��}V��Jc���g� �c�oZW���C���*�D����tm��B�s���!�j�ƽ�`m�|�*��N�T���H��Υ��B�Ѿ�   �   "u�P)��-b�k����n��pͿ�������V3�����z������ο�T��;����c���)��� 5���wJ� ^��֌�f}M��Pq��u�����w��������.&"��FI�2o� 9���`��؝�|ݠ�;)�������8�p�íJ��[#�����n����]z��� ��ý"w��NR�.Ŏ�~����J�x$���   �   � ��'o��?,��T]�)����5�������Uƿ$$ѿ�տ/�ѿHǿ�x��!��\Ɉ�h�^��-�����1精�k�������Hk�|�j�D<���%�Dkj����Hs���,�&X]�J���S8������"Yƿ�'ѿտ��ѿ�ǿ5|��$��̈��^��	-������벾��k����@���Mk�r�j�[:���#�\gj��   �   ��w�n���1���#"�8CI��o��6��$^��՝�`ڠ�&���1툿��p�#�J�X#�����l���<Vz�V� ���ý�w�~JR�?Ŏ�����J��&��Vx�AR)��0b�I����p���rͿ ��q���45�����|�������T�ο�W��ȡ��&c��)�6���8���|J��dｚڌ��M�bNq�r������   �   @U�Qp��e�����^�n�)��B��xV��Ec���g�ľc�YUW��C���*�}��{�Nh��6�s�~�!���ƽ�Tm�*�*��N� �����#���r�Ѿ�g���V�����h��HٿF���"��`���$���'��$������g����1ڿs����l���!W��O�Ѿ�ㄾT�j����9E�(!��b��+���   �   ����,g�U�T�D���غ�(1㾮�����D������z��>���=�f��������X��S�x6���.L����$[O[�#1۽܄H�Ӕ���R�=�����x��]׿��2���_+���;���F��J��-G�g<�,�j�h8�P�׿!���j����=��n��1���E�}սh�N�tԼ�+Ҽ^�=��   �   �������޹��+��rd��K��pu��vz��|vȾR%;9ɾ嗼��������"mh�>/��?�s��z���{f�، ��&���lt���Er���Ⱦ���w_�[阿gPǿ�#��LY�X0��rH�z]��;k��hp�ܜk�ڲ]�<
I��0����S%���ǿk~���~^�ډ�:�ƾ�!n��t��^kd�L��� �x��#��   �   ���;@Z��>�>��Ω��$���f#��+F���a���s�HUz�9�t���c���H�W�&��l ��7����P��Y���^�:��@<�r�;���DE�����J�����\0�"]}�+b����߿���)��1G�ފd�D�}�K�����ڇ�FY~���d��TG�(�(�vk�|߿���<�{���.��(�?������(���wT�п;<�t�<�   �   0�=�=�<@����ۼ^�^�Ԧ��`ؽ-������f�8�����}�ݽ�f��^-n������̿�`�m<��<��<`,�<����#:��;�)�H��������A��i������󿄾��M8�P�Z�R�|��'���W��9 ��k��w<���|�jfZ���7��1�������3n����?��v��5n����$�쵌� �1�`�<N�=�   �   �cA=jA"=<�< ��;H�������e�7���3x�������Q��L��pp�n�%�ll���6}:<�<��= ,=�=�<�}�*����c5��1�����-�L��瑿�Zſ�[��ę�fwB���g������ז�����������I̖�j���=g��A���������Ŀp���&�J�=�<��x�/�2�����$����<6K5=�   �   B=�(=Xb�<8<�xD�ܡ�9O��%���O���f��J��,KW����Xnu�t�;8��<��=|�0=��=�?�<�{��_���LNN��������"�a�i]���7ؿ ��F`/��hW�i��������������j0��o�����`���9g��^�V��.� �9�ֿ]L��V`��J��$��gI��㴽|U��dz�<�.=�   �   ��,=4�=�C�<`�!���μ�jC�bÊ��J��Ed���'Ƚ���b��5ӎ���M�te�p��um<8��<\{=��=T��<�4���
���
J��F��r���]�D���#�Կ�	��\,�^S�X
~�·������������2���P���d����}��R���+�(��zӿ����M\�$~�����B�D��c���Λ�@2�<��=�   �   L<�<�K<h��b��٭��i�½a����������z#�fJ�la�g���Ƚ:č�$H$�(X�(�<xZ�<t-�< �)<جż0�����=�������
��	R�:���a?ʿ~��0�#�.�G���n����.��;����ԫ��Ƨ�/�����h�n�h�G�A#��X��Iɿ9����{P��d	�����9������v���n<t�<�   �   �ٺ��μ��m���ƽ���|7���\�Wqz��ӆ��H��D>���|�� _�E0:�����Eͽ�|�DE��	����; rt9,XԼn����;+�$7������\�?�F��5���F
񿠒���6���X�4nz��Ջ�6������������z���X�:�6��U�i��J���h���P>�����F���'�Ѩ��l�����;��<�   �   j�/��?�������?���}�j����E�;��۾*���ܾ�ξZ��5���n���EC�(	�*��J=�PH��X~�,��Y���t���҅���۾�-(�Y-r�s.����ֿ 7��I"�6�>��UZ���q����J��W<��:or���Z��1?�p"�p2��ֿɤ��Eq��>'���پ���P>��ӊ��ۼX�G�\����   �   ��˽�5"�H�l�+���};+������ !�J)��,�i_)�ŭ�ys�o>����ξQ���o��T%�s�ѽ*�w�����yO��=����^�[��	��j�M��{��/���翺��ޟ#���9���K��pX�2�\���X�ąL��-:�D$�&B��#�Z���U���iM�rD�����0F\�ϴ���}�@'��`�&xl��   �   �52�)#���V��:
��;���8��zS���h�Jrv�QJ{�J�v��ui�9cT�?�9��4�����Q�~���ݴ4�5	佧򍽌�T�аz�O�ͽu92�����Cu徻(�>'i����������=� ���K�Z�(��
2�Bv5� T2��)�����*	�0��&¿<홿l<i�.�'�2�供Œ���0���ɽ�-s�@�L��ĉ�n�߽�   �   �=����ƾ�����0�D�Z������w��􉡿�����ĭ��Ԫ�� �����.-��$�[�#�1�K��VȾ�7��D#4����h��t��RF������a�&?��C_�%48��Fu�a���\l���ݿV���K����f@����:��#���Vw޿H%���?��=�u���8�"~�02���6a��)�S�����{��"���f޽��2��   �   I�þ��
�:;�Q&p��6��G*���Ŀ��տH����m��^�ֿ�Ŀ�譿�ݓ�-q���;�u��+ľvZ���*$�1�ʽ�c��<���lʽY�#��g�þz�
��5;�e!p�"4��'��k Ŀ��տy��R�������ֿk�Ŀ!歿Jۓ�^)q���;��r�](ľdX��`($�=�ʽ�d��D?���rʽ3�#����   �   b��78�YKu�����o����ݿ7�� N� ���B������w���9z޿�'���A��h�u��8���z4��u9a��*�M�����{�����^޽щ2��9��T�ƾj��ȏ0�Q�Z�ڎ���t������C���G����Ѫ������	���*���[�ׇ1�����Ⱦ&5���4��Ὗg����]J��z����a�:C���   �   � (�.+i����ߣ��GA����M���(�D2��x5�BV2��)�Z��,	����'¿��>i���'����ǒ�\�0�K�ɽN*s�P�L�����z߽N/2����"Q��g��7���8��uS��h��lv��D{���v��pi��^T�=�9�[1����컾Y���v�4��佻��T�дz��ͽ�=2������y��   �   ��M��}�����	��p��ڡ#��9�| L�psX���\�d�X��L��/:��$�VC�w%����W��(kM��E�㽶��G\�W���|�}�!��V�^il���˽�."���l�薠�8;����������)���,� [)�©��o�!8����ξ�L��f�o��O%���ѽ��w�@��8�R�����,�^��
��c���   �   p0r�c0��4�ֿl8��K"�<�>��WZ�R�q��������=��tqr���Z�23?�.q"�@3�<�ֿhʤ�>Gq��?'���پ^	��~>��Ҋ�0�ۼ�nG��虼�/�6��M�� �?�n�}���=���;��۾��ྔܾ��ξ�T���|��'j��X?C�F	����"@=��<����}��!��Q���>���ԅ���۾0(��   �   �������g���(�6���X��pz�:׋����䄙�B�������z���X��6�HV��i�K��i��!Q>���������'�����D���pP�;8 <��׺h�μ2�m� �ƽ���Iu7���\��hz�:φ�.D���9����{���^��):�b��U=ͽ�|��1�0կ� "�; u9H]Լ�á�l>+�K9��� ����?��   �   k����@ʿb��D�#���G�|�n����<��J����ի�vǧ��/��_��,�n��G�VA#��X�+Jɿ[����{P��d	�e��Z9�3����o��h�n<l�<hK�<��K<p�����˥��B�½Q������l��ru#�E�v\�r���@Ƚ�����=$���W�8�<�a�<|0�<��)<��ż=���|�=�����T�
��R��   �   +���9�Կ��	�X],�_S�|~�s���� ������!�����������d��&�}�(�R�~�+����yӿ^����\��}�!���B�D��a���Ǜ�@9�<x�=�,=t�=LP�<�z!�h�μ�aC�p����E���^���"Ƚ������+ώ�ȰM�0Z�0ʿ�(�m<8��<H|=��=��<l;������J�H����<�]��   �   �]��q8ؿ\���`/�BiW��������' ������i0��V������%����f���V���.�����ֿ�K��l`��I��#���I��ᴽ�N��`�<� .=�B=��(=e�<(<tD���68O�>%���O���f��~�q�LW���� su��i�;X��<V�=��0=��=t:�<�����þ��ON��������a��   �   z���S�Կ(�	��\,�^S�&
~�����������������������c��Ԍ}�*�R�®+�����xӿ�����\�}�'�����D�E`���Û��;�<H�=��,=Ω=�P�< x!��μ~aC�d����E���^���"Ƚ������ώ���M��Y�0ȿ���m< ��<�|=��=䤂<7������J�G����5�]��   �   ���#?ʿJ��ڻ#���G��n�E��q��Y����ӫ��ŧ�.�������n��G��?#��W�zHɿ����yP�,c	�����9�����g����n<��<�M�<H�K<���T������(�½:������b��fu#�E�d\�U���Ƚ����(=$�H�W���<(d�<4�<`�)<Ȫż����=�������
��	R��   �   �������d	�����6���X��lz��ԋ���I������S��̴z���X���6�fT��f�>I��Eg��qN>�ȟ��� ��,	'�c���@����l�;)<@y׺��μ��m�ʆƽ���8u7���\��hz�5φ�&D���9����{���^��):�@���<ͽ�|�X/��ǯ��5�; �x9�QԼ%���;+��6�����ϓ?��   �   ,r��-����ֿ06��H"���>��SZ�l�q�:������:���lr�d�Z��/?�rn"�
1���ֿ�Ǥ��Bq��<'�E�پV���:�p͊� �ۼ�]G��㙼z�/�{5��$����?�V�}���6���;��۾��ྊܾ�ξ�T��~|��j��)?C�
	�G��:>=��6��0�}�������4���х�o�۾�,(��   �   ��M�kz�����<�翌��b�#�Κ9���K�LnX���\�@�X�>�L�x+:�J$�r@�� �����S��efM�B�
����@\�����d�}���:R�~fl���˽�."���l�ז��+;���������)���,�[)�����o�8����ξ�L��$�o��O%���ѽ��w�f~���hL���
����^��������   �   �(��$i��������z;꿤���I�V�(��2��s5��Q2�J)�z���(	����B¿�ꙿx8i��'����,�Ӆ0���ɽs��L�˻���y߽�.2����Q��W��7��8��uS��h��lv��D{���v��pi��^T�4�9�O1������뻾,����4���S퍽,�T�^�z�V�ͽ�62�ȃ���r��   �   }]��18��Cu�b����i��'�ݿ��J����H>����(��=����s޿"��;=����u�ׇ8�F{��-��N0a��$�����{{�K��o\޽,�2��9��8�ƾa��0�L�Z�؎���t������B���F����Ѫ������	���*���[�ʇ1����VȾ�4��4���d��,��B��8��m�a��<���   �   }þ7�
��2;��p��1��`$��[�ÿg�տ�Έ�����=�ֿ�Ŀ�⭿hؓ�f$q���;��o�P#ľ�T���"$� �ʽo\��47���iʽj�#�����B�þp�
��5;�b!p�!4��'��l Ŀ��տ{��S�������ֿj�Ŀ歿Gۓ�T)q���;��r�+(ľX��\'$��ʽ�_���7��ogʽ�#���   �   �6��^�ƾ���w�0�B�Z�v���r���������󽭿OΪ�c�������'���[���1�8����Ǿ�0��.4����'_���|�B�����8�a��>��6_�48��Fu�`���\l���ݿW���K� ��f@����:��"���Tw޿E%���?��4�u�{�8�~��1���5a�K(����\~{����fX޽��2��   �   o*2�����L�������3��~8�qS��h�Egv�?{�?�v�Bki�{YT��|9�@-�'���h滾փ��n�4�����捽X�T���z�Ѕͽb82�9���u徴(�<'i����������=� ���K�\�(��
2�Dv5�T2��)�����*	�-��#¿9홿d<i��'� ��EŒ�։0�O�ɽ�"s��L�Ǹ���s߽�   �   ��˽�)"��l������;���������
)�6�,��V)�r���k��0��J�ξtG����o��H%���ѽ��w�Xt���,K��u����^�"�����h�M��{��2���翼��ޟ#���9���K��pX�4�\���X�ąL��-:�F$�$B��#�X���U���iM�`D�Q���QE\�����H�}�(�,N��]l��   �   Z�/�1.��9����?���}�p�������;��۾ |���۾�~ξ�N��.w��te��f7C��	�I���.=�D ����}�h
��
���j��Z҅�}�۾�-(�[-r�u.����ֿ7��I"�8�>��UZ���q����K��X<��:or���Z��1?�p"�p2��ֿɤ��Eq��>'���پ���@=�KЊ���ۼ�TG�Lי��   �    �ֺ�qμ�m�~ƽ=���n7�~�\�}`z��ʆ��?��a5����{�n�^�z":����,2ͽ��{���po���x�; �~9�IԼ����:+��6������[�?�G��8���I
񿠒���6���X�8nz��Ջ�7������������z���X�:�6��U�i��J���h���P>�ߢ�����'�i������s�;8<�   �   U�<�K<�q����(���a�½C������|��o#�u?� W�6����	Ƚm���V/$���W���<(s�<@�<��)<��ż������=�������
��	R�<���d?ʿ���2�#�0�G���n����.��;����ԫ��Ƨ�/�����f�n�h�G�A#��X��Iɿ9����{P��d	�i��`9����|m����n<�<�   �   ��,=��=�W�< 0!���μ|ZC�E����@���Y��aȽ����~��ʎ�\�M�0I� ���x�m<��<j�=��=��<00��-
���
J�|F��o���]�E���#�Կ�	��\,�^S�X
~�·������������0���P���d����}��R���+�&��zӿ����L\�!~�����
�D��b��ʛ��8�<�=�   �   2�8=hj=Y�<��; τ�f��z�e�5��Dۤ�����楽W=���k��D ��?���%;�U�<�L=�*=W=X|<(�߼J�˽QY����i_�n=k�����o�࿢3�4�6��?a��L���*��~������6i�������p��n��!��P�`�b!6�r���߿�>�i�	'�K����T��ý�q��P�<8$=�   �   ��"=y =�2u<pFһ ��� �Y�H��Qи�zνKֽ�Ͻ�ٺ�]<���_a�h��xa��E<8)�<�=|�=��]<����Ƚ�T�����-l�Bg��٣�(�ܿ����i3�"�\�7m������j��2����������/c��߀���H����\�  3�^f��ܿ�"����e��<�Ʉ��ΈP��������d��< /=�   �   ,��<��<�{b��+�|��p�ѽTH����� (��-�7�(�������ս��`06�������;���<�³<�7�;�m�M���H�D������@�Z�T���~ҿ���X[*�D�P��z�Bx��	¤�����d�����=Ȥ�Zt���z�@�P�d*����vlѿ����^�Y��������%D�޵�Ԏȼ��6<���<�   �   @߸��T���P��J�ս��QB��i�9܃��Ǎ�wL��s��ne��E�j��2D��E�f�ڽ$����o��� �4;�&6�����E񭽐�4���������G�����H��
h�������>�r�b�ϖ��X����������-��m��B��� c��>�zg���������%����F�P��m៾�X1��J��� ۼ ��9`��;�   �   �F�0o��J���<K�Ʋ�����3���׾���	��;�kؾy¾&���Ɔ�*�M��!�v���^P�<�Լ����$��Xb���|�����~��~/�'A|��ϫ�JJ߿���@�(��HG�ĵd�t~�8����և�V~���d�oG��)�4y��߿+|��Ä{�ۺ.�Gl侁���������x��p����c���   �   1{۽LY,���y�|ۨ��&׾�)��V��O&��0��24�N�0��&����X��F@ؾ����� |�̅.�=�߽S���.�.�V�/�࣏�����j�e���7:���V�IQ������񿚘�(y*���A��\U�D�b�6jg���b�@�U�B�Ʊ*����%�Wo��a%��BV���x���~th���L;��F�&��B&��t���   �   ��<��C����þ�� �P!���@�$�\���r�-s��낿�����-s�E]�^A��!��h���ľ�+����>���򽁘��^xi�򎈽��۽�^<��%'�ѐ/��s�����sɿ;��h8��� �n�/���9�*9=���9���/��� �,v�����ɿr����r��V/���ﾼ9����:�Q�ؽ>���4^c�����(���   �   {��ƆоS���8��5d����\���87�������Ǵ�x���Dy��W����t��E�d�c9����G=ѾR��P$>�s��ɂ���<��c������m�p�^p	�FY@����T5��A'ſ��.�P��n���������L����ǄſQu������s@�lj	���� Gm�����߳�����0����7)=��   �   �;�_���C��z�i��Q��A�˿��޿q����&����޿`e̿����@{�]�C����4V;8���8�-��Qٽȏ��u����)ٽ
�-��ψ��;l\���C��}z��f���M����˿�޿{����_��m�޿2b̿R�������^{�M�C�����R;�����-��Oٽi���·��/0ٽ�-��ӈ��   �   Es	�]@�y��)8���*ſ���4�x��<p���������N���M�ſdw��b��+v@�4l	�r����Im�D���߳�5����ڝ��/�x#=��v��+�оO���8��0d����,����3��.���BĴ�%���'v������7r���d��9�:��K9Ѿ���� >�X��x���3>��0g��o����m������   �   ��/��s�C���vɿ���b:�° �ڸ/�,�9��;=�&�9��/�t� ��w�f ��4�ɿ��Xs��X/�#��6;��t�:���ؽm����Uc�{��`����<�?��Øþb� ��K!���@�ط\�R�r�Ep��)肿����(s�K@]��YA���!��e�U�ľj(��j�>����m���Xwi� �����۽�b<����+��   �   ��V�^S��������d��@{*�V�A��_U� �b�mg�N�b���U��B�X�*�.���'��p���&���CV���ײ���uh�l���9����&�8&�	m���p۽ZR,��y�֨�o ׾�%�uR�}K&�Y�0�&.4���0��&������:ؾ�����{���.�#�߽軆��.�Μ/����������j������<��   �   XD|��ѫ��L߿v���(�$KG�P�d�X~��Ç�0���ׇ��X~���d�~pG� )�z� ߿}���{�û.�]m�	��ؚ�����l��4솼pL����E��d������4K���������-��q~׾��6��i4�Bؾ����Q	������M����n��jTP��Լ���Ԫ�de����������w�/��   �   �����J��Aj����@�>��c����wY��	 ������.��2n�����dc��>�h���������&��N�F�����៾�X1��I����ڼ Τ9���;����,7��fG���ս��EJB���h��׃�!Í��G���
��4a���}j�,D�l@�k�ڽ(����e�h����4; 6�����z���d�4�Q������̹G��   �   ����ҿ���z\*���P�Դz�Ly��(ä���f�����ɤ��t����z�̈P��*����lѿ����y�Y���ڢ��n%D��ܵ�h�ȼ��6<�<Ƞ�<x�<HLb���+��s����ѽC�"����'���,���(����ܾ�ڄս�옽t%6�Hχ�/�;t��<�ų<�2�;t�BP���H�>�����*�Z��   �   �ڣ�H�ܿ����j3�$�\��m��Ŗ��ek��׈���������c������H����\� 3�Lf��ܿ�"��H�e�8<�,���ƇP���������Č<3=2�"=�~ = Lu<�һ�����Y��B���ʸ��tν�Eֽ�Ͻ�Ժ�$8��XXa�x���N�h�E<x-�<�=*�=H�]<��༹Ƚ�T�@���Km��	g��   �   ������4���6�@a��L���*��<~������6i�������p��/��� ����`�� 6���l�߿��L�i�J&��I�� �T���ýk�����<B$=�8=�k=�[�<�&�;�̄�X����e��4��ۤ�����F楽�=����k��E ��A���%;�R�<\K=T�*=�T=�|<��߼��˽�Y�.���*`�e>k��   �   �٣�[�ܿ����i3��\�m������_j������n����}b��/���H����\�R�2��e��ܿ�!��:�e�y;�*���t�P�@������Xǌ<�3=ȣ"=�~ = Mu<
һ����t�Y��B���ʸ�~tν�Eֽ؀Ͻ�Ժ�8��*Xa�N���M���E<L.�<��=�=�]<H�� Ƚ¬T�;����l��g��   �   3���>ҿ��� [*���P�8�z��w��A������c�����Ǥ�Rs��&�z�ֆP�D*�ƒ��jѿL���v�Y�������"D�zٵ�0ȼ8�6<T�<ࢽ<�<`Jb�x�+��s����ѽC�����'���,���(����˾���ս�옽�$6�8·��5�;Ȕ�<hɳ<�H�;�k��L��	H�M������$�Z��   �   ����H��!g������>�,�b��� W��T��A���!,���k�����c�X�>�"f�����B���7$����F����ߟ�PU1�E���ڼ ��9 �;`x��@5��G����սi�4JB�x�h��׃�Í��G���
��,a���}j� ,D�L@�!�ڽɒ���d����5;��5�4����ﭽ��4����������G��   �   �?|��Ϋ�I߿$�� �(��GG�Գd�~�����,���ԇ�8S~�6�d��lG�)��w�K	߿-z����{�n�.��h��
�����X�������ㆼG���E�Rd������4K������-��k~׾��/��`4�7ؾ����C	����s�M����m���RP�,~Լ$����� `��p{�ڇ��@��}/��   �   �V�!P�������\���w*���A��ZU���b�^gg���b���U��
B���*�(���"��l��M#���>V����Э��oh����:4��z�&�^3&��k���o۽R,���y��ը�b ׾�%�qR�yK&�U�0�!.4���0��&������:ؾ�󩾦�{�`�.�&�߽[���<�.�>�/�����"��ڲj�����	9��   �   ��/�Is����qɿ����6��� �J�/�B�9��6=�<�9�|�/�b� �2t�]��#�ɿ�����r��S/���-6����:���ؽ�|���Nc��x����d�<��>����þ[� ��K!���@�Է\�N�r�Cp��'肿����(s�C@]��YA���!��e�7�ľ@(���>��������oi� �����۽&\<��욾�$��   �   �n	��V@�t��B3���$ſ���t�^���k���H��� ��J���激�ſ|r��`���o@�vg	�����^@m����Q׳�����}ם�g-��"=��v���оwO���8��0d����*����3��-���AĴ�"���%v������4r��	�d��9�-��&9ѾF���>����}���8���^����b�m��ﹾ�   �   9;Z�m�C��yz�)d���J��o�˿��޿�~���g�꿏�޿�^̿��������<{��C�K���M;�����-�eFٽ���}���&ٽ�-��ψ��;a\�}�C��}z��f���M����˿�޿|����^��k�޿0b̿Q�������V{�C�C�����R;������-��LٽQ������~$ٽ��-�f͈��   �   �s��}о�L�+�8��,d�<��Y����0��ۀ�����������r��P���Jo����d��9�����3Ѿ���>�����x��66���^��T��G�m�9�Pp	�@Y@����S5��A'ſ��.�P��n���������L����ńſOu������s@�Yj	�м��'Fm����e۳��֝�1)�=��   �   ��<��;��C�þ�� �\H!���@��\��r�vm��A傿'����"s��:]�UA�O�!�bb�u�ľ�#��,�>�d��`����gi�c���7�۽�]<�Q�&�ɐ/��s�����sɿ;��h8��� �n�/���9�,9=���9���/��� �,v�����ɿp����r��V/����f9����:���ؽ�~��VMc��u������   �   �h۽�L,���y�~Ѩ��׾�"��N�PG&��0��)4�:�0�n�&����H��+4ؾ~��{�ly.���߽������.���/�n���v��@�j�,���+:���V�JQ������񿚘�(y*���A��\U�F�b�8jg���b�@�U�B�ȱ*����%�Vo��_%��BV���9����sh�����6����&�/&�g���   �   ��E��\��t���-K�⩅����(��Ax׾s��[�꾎-澠ؾ�������Ľ��e~M���c���BP��fԼ~������^���{�c���V��~/�(A|��ϫ�MJ߿���@�(��HG�Ƶd�v~�9����և�V~���d�oG��)�6y��߿-|����{�Ӻ.�l�.�����P���$���ކ�h:���   �   �?��� ��@����ս���CB���h�uӃ�����C��7���\��*uj�f$D��9��ڽ�����U��|���5; |5��������4�嫡�����G�����H��h�������>�t�b�ϖ��X����������-��m��B��� c��>�zg���������%����F�@��6៾X1�.H����ڼ �9 &�;�   �   ���<��<h(b�v�+��l����ѽh>����T�'���,��}(�������3{սh䘽�6�L���Ѓ�;L��<�ճ<�n�;Td引K���H�&������?�Z�V����ҿ���Z[*�F�P��z�Bx��	¤�����d�����=Ȥ�[t���z�@�P�d*����wlѿ����[�Y���ߢ��x%D��ܵ��ȼh�6<�
�<�   �   ֤"=$� =[u<0�ѻ�u�� �Y��>��Ƹ�Hoν @ֽL{ϽlϺ��2���Na����0�hF<X9�<J�=(�=8�]<X��*Ƚ��T�����+l�Ag��٣�*�ܿ����i3�"�\�7m������j��1����������.c��߀���H����\�" 3�^f��ܿ�"����e��<�������P����,���@Č<�3=�   �   ��9=ڈ=��< ��;PO�����6�e��<���Ť�����gU���[���i��4�d� �g;s�<�=��/=4=�;�< �׼1)ʽ2�X�Rq���p��qk��ܦ�G��Zf��6� �a�;����ʠ�t@������>��S���?���ʠ�z�����a��6�*O�[��!�����j����^ ��Z�U�_GĽT-�� ,�<�9%=�   �   ��#=*v=��w<�wϻ����2	Z�Mz������d�ν�#ֽqϽ���\���v^��g �6�x�W<���<��=�=H�o<�ؼ<[ƽ�T������~��>g����eݿ����3�ށ]��߅��5���,���Y������+W��=)��y3���݅��z]��3����U�ܿ����;�f�\���3��=Q����\����[�<�L=�   �   �I�<�<��a��A,�ؔ��Tҽf���L�qA(�L&-�-�(����DW�cTԽ�d��`2�x.����;л�<��<��<�ݼõ��@{G�c���g���[��̛�`dҿz#���*��YQ� �{�����~��Rݱ��.��ر��v��!����{��KQ���*��	�d$ҿՂ��
kZ�wP��@����D��K��`:ȼh�9<���<�   �   �⵻(�������e�ֽ;��(�B��i�H9�����E����5��8m��4Wj���C�����;ٽ�ˆ��u��/����w;@��(��v���L4�❡������G��Ꮏ����C���j��6B?�f�c�(&��#��`֞�⨢��Ξ�q������̽c��,?������3c�����#fG��"��e����1�Ü��p�ڼ '�9p��;�   �   �[F����4��K�(2��]���\����1ؾ0��U�뾈��tXؾ¾� ����� M�
l��Ϸ�&�L��3ͼ@p���e	�G����!���P)���/�־|��/����߿>��J�)��H�(�e��9�jY��s��dQ��z�D�e���G�n)�*��<�߿�����A|��B/���mr��X��
��q�xF������   �   0ܽv�,�v�z�����-�׾ާ������&��1���4��"1�Y�&��������?ؾ�ة�Ύ{���-�Od޽?����+��,�w{��&���j��	����B8W�@���E��:����+���B�R?V�z�c�;h�b{c��'V��tB��+�B������������l�V�+�U.��k�h����I����&�2&�詂��   �   Ђ=�GČ�9^ľ�^���!��A�q�]���s�7ր��A���ր���s��]�R�A���!�rq�5�ľ���(>����n���4g�񙇽�E۽�[<�y%�����0���s������ ʿ˃��|���M!�ta0��S:�$�=�bI:��O0��8!�v���[����ɿfg���{s�Y�/���򃚾�#;���ؽ�n���9c�����o4��   �   R�-EѾ����?9�!e�(���Y9��%ɨ� ���?��!��Ĩ��3������,e��99����wJѾ=����=��;�y���H���鴽|��'?n��d����	���@�&Q��Lʢ�Q�ſYh�h��,O����������C�`}�]K��ſ�����5��(�@��	�����(~m�0��害�1s���ԝ�\��O�=��   �   ��;��� DD��t{�����b ���̿$[߿R>뿿R��6��M߿�̿�﴿@U{�\&D�W���;���"�-�g�ؽ����+���$ٽ��-��(��~�;V���?D�so{��������I�̿EW߿Y:��N�3�qJ߿��̿�촿�왿2Q{�K#D���k|;�����-�M�ؽr��/��+ٽ��-��,���   �   ��	���@��S�� ͢���ſ
l�n��VQ����֊�(��vE��]N翈�ſ����Z7����@���	������m����򮳽�p���ϝ�
��2�=�퐾�?Ѿ7��H;9��e�=���&6���Ũ����g<���
�������0��8����e�#69����tFѾi���6�=��7�!�������.�>��En��h���   �   B
0���s�/����#ʿE���x���O!��c0�`V:���=��K:��Q0��:!���^����ɿi��~s�'�/��p���%;�w�ؽ�l���1c�����*�|=�Ŀ��rXľ7[�k�!�C�A��]�ڐs�LӀ�?���Ӏ�_�s�U�]�(�A��!��n�ɌľV��x#>����k���3g������J۽`<��(��J���   �   �;W�V������C��l� +���B�
BV�Z�c��=h�~c� *V��vB�x+�� ���|������V�K��/����h�D���G��.�&��'&�8����ܽ~�,���z�$~����׾�����S�&�`1��4�%1�-�&������:ؾ&ԩ��{���-�-]޽�:����+�h�,�~����v�j�7��y���   �   �|��1�� �߿����)��
H���e��<��Z���t���R���!�8�e��G�8o)�����߿���� C|�kC/����r��������l�@6�������KF���~-�	�K�Z-��Ԫ��7���3+ؾX��{����FRؾ¾�������m�L��f�Hȷ���L� 'ͼ�k��~g	�J��`�t����,�1�/��   �   ㎿{���y�������C?�|�c�e'������מ�I���>О���������c��-?���������c�������fG�#��e����1�������ڼ H�9P��;�����c��~���*�ֽ�����B���i��4���������/1���h���Oj�I�C�h���2ٽ�Ć��k�����@x;���4���y���O4����"����G��   �   �͛��eҿf$��*�j[Q�ƕ{�������qޱ��/��ٱ��w�������{�LQ��*��	��$ҿ����'kZ�tP��@��z�D��J��3ȼ`�9< ��<@Y�<�<��a��3,��ϔ�)Kҽ)��G��;(�� -��z(�j���R�JLԽ�]��ht2��� ��;�ì<�<��< �ݼݸ���}G�[�������[��   �   �	���ݿ����3��]�1���p6��F-���Z��<����W���)���3���݅��z]��3����$�ܿ_���іf����^3��<Q����p����b�<�P=�#=�{=�x<0<ϻ�z����Y�$u�����ՃνHֽ@Ͻ��� ��^o^��a �`#���W<L��<��=��=��o<��ؼ^ƽT������i@g��   �   �ݦ���࿼f���6�~�a�~���*ˠ��@������>��9����>���ʠ�6���^�a���6��N���࿍�����j�Ѽ�?�����U�EĽ�&��1�<z;%=2 :=^�=��<@��;M�����`�e�^<��sŤ������U���[���i��5��􏼀�g;,p�<�=��/=�1=\6�<��׼�+ʽԃX�sr���q��rk��   �   ����ݿ����3�Ё]�y߅��5��?,��rY��!����V���(���2��&݅��y]�<�3�>��8�ܿ����f�>��]2���:Q�`���D����e�<�Q=��#=�{=px<p:ϻtz����Y�u�����΃ν:ֽ/Ͻ�����2o^��a ��"��W<��<B�=��=��o<@�ؼM\ƽ�T����1�Z?g��   �   �̛�!dҿD#���*�rYQ�,�{�����}��cܱ��-���ֱ��u������{�JQ���*����"ҿ����!iZ�O��>����D�SG���*ȼ �9< ��<<[�<�	<��a�H3,��ϔ�Kҽ��G��;(�} -��z(�]���R�1LԽ�]���s2��
� ��;�Ŭ<��<h�<��ݼ����J{G�l���b���[��   �   -Ꮏ���\������NA?� �c�K%����՞�{����͞���������c��*?����ݱ��ea�������cG�
!�Cc��j�1�3�����ڼ �9���; {���a��1����ֽ���x�B�r�i��4���������(1���h��~Oj�2�C�N���2ٽ�Ć��j�`��� 2x;@뺨��Tu��BL4�o���(��)�G��   �   {�|��.��h�߿d��*�)�.H�4�e�B7�X���q���O������e�X�G�Pl)����˜߿�󫿓>|�@/�3��o��m���엽f��-��$��IF�"�U-���K�L-��ʪ��/���,+ؾR��t�����=Rؾu¾����񕆾J�L��f��Ƿ��L�|!ͼ�b���`	��
��7�H��(���/��   �   �6W�����	��D��d�b+���B��<V�Άc�@8h��xc�%V�JrB��+�x����j����}��#�V����*���h����
B��̪&��"&�̠���ܽ8�,�^�z�~����׾�����N�&�[1���4� 1�(�&������	:ؾԩ���{�@�-�5\޽9����+���,�Kx��f����j�'��ڀ��   �   @0�R�s�����ʿ9������K!�N_0�nQ:���=��F:�8M0��6!�z��X����ɿ�d��yws�%�/���d���:;���ؽ g��"*c�����7)�{=�����]Xľ/[�e�!�=�A��]�֐s�JӀ�?���Ӏ�X�s�N�]� �A��!��n���ľ/���">�6��i��X,g�����A۽DY<��#�����   �   ��	�@�@�~O��7Ȣ���ſWe翬��6M����`�����XA�X{��G翸�ſ̫��V3��U�@��	�����wm���k���3k��̝�؄�=��쐾r?Ѿ/��A;9��e�:���$6���Ũ����e<���
�������0��5����e�69����SFѾ0�����=�\5ｎ��� ~���䴽�~�s;n�b���   �   
�;����<D��k{�G���;����̿�S߿�6��J�	/뿑F߿�̿~鴿�陿L{�D����1w;������-���ؽ#���&���!ٽ��-��(��X�;K���?D�no{��������H�̿EW߿X:��N�3�oJ߿��̿�촿�왿+Q{�B#D����>|;6����-��ؽe��5'��nٽ3�-�_&���   �   ꐾj;Ѿ~���79��e�����Q3���¨�O
���8��Q�������-��J����e��19�D���@Ѿ����r�=�-�y����{���䴽$��\>n�od����	���@�#Q��Jʢ�P�ſVh�h��*O����������C�^}�[K� �ſ�����5���@�Ӡ	�R���V}m��������ml���ʝ����Қ=��   �   �v=�V����SľVX���!�}A�V�]���s�zЀ�<���Ѐ���s���]�L�A���!�k��ľ����:>�v��b��R$g�]���B۽�Z<�(%��v��0���s������ ʿ˃��|���M!�va0��S:�$�=�bI:��O0��8!�v���[����ɿdg���{s�N�/�o𾟃��i";�]�ؽ�h���(c�����<#��   �   �ܽ�,�r�z��y���׾̠����!�&��1�_�4��1���&����ڹ�~3ؾ�Ω��~{�H�-��Q޽z1��z�+���,�w������j��	�����?8W�A���F��;����+���B�R?V�z�c�;h�d{c��'V��tB��+�B������������f�V��.����h�����D���&��&�@����   �   \?F��崽2(�Q�K�:)��便������$ؾ�澛y�	�澣KؾP¾R���%���8�L�+`�O����L�L
ͼ�R���[	��	��n����*)���/�ؾ|��/����߿>��J�)��H�(�e��9�jY��s��cQ��z�D�e���G�n)�,��=�߿�����A|�{B/���r��D����g��(��h侼�   �   �B���L��!���܄ֽ����B�Щi�}0��a��܃��v,��ld��Gj���C����Y'ٽJ����[����@�x;�S�|��;t��/L4�����x����G��Ꮏ����E���l��6B?�f�c�(&��"��`֞�㨢��Ξ�p������ʽc��,?������5c�����fG��"�ve��6�1�R���|�ڼ ��90�;�   �   8c�<�"<�ga�2(,��Ȕ��Bҽp���A�
6(��-��t(����JM��BԽ<U���e2���~�`�;Tլ<���<H<T�ݼ5����zG�C���a���[��̛�adҿ|#���*��YQ��{�����~��Rݱ��.��ر��v��!����{��KQ���*��	�e$ҿւ��kZ�oP��@����D�\J���0ȼ �9<���<�   �   ��#=4~=`%x<�ϻ�n��6�Y��p��A󸽐~ν�ֽ�	Ͻs������e^�Y �����W<��<�=��=��o<\|ؼyZƽ�T�u����~��>g����fݿ����3���]��߅��5���,���Y������,W��=)��y3���݅��z]��3����U�ܿ����:�f�[���3���<Q���������b�<bQ=�   �   ��E=ܭ+=��<��< vB�4����O�_e���<������?=���v���OP����YJ���<ȼ�<j&=�a?=�*=l��<���!Թ�\�L�-���~ �Ɯb���ٿ�i��W0��Y�������V)��E ��ѝ��� ��{2��^������t]Y��0����`ٿ�����b���:��@HK�����@���<�d1=�   �   ��/=[=���< ���\ϼ8jD��z������߽����ǽ۲��3�������>E�D�Ҽ @��I�<�f	=�)=�8=d��<�/��J1���sH�?��XJ�N�^�5���տ�"
�HZ-��T��E��/G���D������]��C��OE���U��Uc���DU�r�-�rZ
��տsX��ٛ^�)����AG�9���$`��L��<��"=�   �   8��<��Q<�U�~���؈���Ľ��������[��#�3E��������x�Ľy6���d���&�x�A<���<�e�<0:]<������P<�Lr��6�n�R��B��&5˿���x�$���I�mq�Ì��-��������������������uq���I�r�$�4���_˿�T��(�R�t�
�B驾B�:�z����񡼈ev<��<�   �   ����<�ϼ�p�7�Ƚ�Z�i9���^���|�0Շ����B���	L|���^��9�)�/�Ƚ>tq�̼Լ ����< �M;��	w��d�)�������	h@��ɉ�-	��N�򿚬��}8�|)[�L�}��������v���Ǘ�׉���=}��Z� j8����6����ĉ��E@��:��`���h�(���������;xR<�   �   �0�ꧽ�,�<,B��O���ў�	����Ͼ�tݾz'⾬Eݾ�PϾ"���\f�����,�A�.��E��B�2�X�����S����֍�މ�ƅ�2�ܾ�)�ܬs��O��vrؿU���#���@��]�.u�$���?�������z�t���\� �@���#�p1�Gؿ�0���ts���(�"ܾ69���b����Jۼ�hD�H���   �   ��ͽ* $��zo�����I�Ͼ�z��mO��� ��*�V�-�x*�G{ ���������ξ������n���#���ͽ�1o�h��@��> ���
����^�J¸�O��CfO����������Ba�r%��;�JtN���Z�>A_�ҭZ��N��Z;��	%�~�p�鿑]��8d��NO��m�6����]�{��w~�\���v���m��   �   �4�Z�������b�����:���U�-)k��x�NQ}��x�Ѿj�yOU��!:�ю����Wڻ��)���|3�_�ན����.N��Lu�K�˽�H2�^4��9��)��Bk�l0��٘ÿQ���5
�.�Tw*�<�3��7��3��*������	��쿩ÿ�Қ��j��)��e澊����f1��sʽ(s�R�L��V���M��   �   ڟ����Ⱦ[�	��2��;]��������4���&���)�������梿���W���q|\��	2��	�@=Ⱦ����p3�W߽�,��Ҋ{�)
��)����b�����:��:�a�w��m������;�������	���v�n���s	�� ��"i߿��K����w��{9�z'�����j�a�,K��*��&�z�Z.��Α߽J4��   �   �jžm��P=���r��딿�&���/ƿ0ؿ��㿢w翆a�]�׿�ſ;����n���r�ҫ<�d��m�ľ�����#���ɽ�+���d��7�ʽ��$�w ���ež�i��L=���r��蔿y#���+ƿC,ؿ����s��]��׿ҥſ����rl���r�ب<�&��=�ľ�%�#���ɽi,���g��[�ʽb�$����   �   
���:���w��p��΍����������	�"�Bx�z���u	�+$��l߿K���O����!w�2~9�7)�� ��5�a�zL��*��`�z�Y)����߽b4�����>�Ⱦ�	�Ũ2��6]�������O1���#��G&��R����㢿W���𪂿]x\�P2�1	�^9Ⱦ���Pm3�G ߽�+��H�{�1�����B�b������   �   �)��Fk��2����ÿ����7
�R��y*���3�&7�Z�3��*�P��t�	�5쿮ÿ6Ԛ�Y�j�m)�Ah�����-h1�tʽ�s�f�L�yP��UD�i�3��������{�����5�:���U��#k�?�x��K}��{x���j��JU��:�j��"��ֻ��&��x3���ཅ����-N��Pu��˽�L2��7�����   �   miO�����������b�t%�V�;��vN���Z��C_�X�Z�N��\;�^%���W��_��Xe���O��n�d7���]����t~�*���l���m���ͽj�#�;ro�I�����Ͼ�s��bK��� �s�*���-�,t*�=w ���������ξ�����n���#���ͽL)o�F����������<�^��Ÿ�����   �   ��s��Q���tؿrV�4�#���@�^]��u���������N�����t���\���@���#�D2�`Hؿ�1��#vs���(�3ܾ�9���b����,@ۼ�HD�lh����0�৽6&�f$B��J��i̞���O�ϾPnݾ� �C?ݾ�JϾ�����a�����ήA�< ��>���2� �����S����ٍ����Uȅ���ܾT)��   �   -ˉ��
��p����8�p+[���}����u���w���ȗ�ފ��>?}�R�Z��j8�D����_���ĉ�%F@�);������T�(�����t�����;t<@G���nϼ�p�R�Ƚ(T��a9�h�^�2�|��Ї����޶���C|��^�|9��#�t�Ƚ�fq���Լ@n���< �M;���z���)����$���2j@��   �   D���6˿n����$�R�I��nq�Č��.������������i��'����vq�|�I���$�j���_˿�T��C�R�s�
�驾��:� ����꡼0xv<��<���<��Q<P'�����Ј�P�Ľ����Z��WV���#��?����{�����Ľ�/��8Z���&�8�A<���<i�<88]<칮�����R<�3t����H�R��   �   �5���տ�#
�[-���T�*F���G��xE��d����]������E��1V��oc���DU�l�-�`Z
���տ?X��s�^��(�����@G�����Y��4��<^�"=@�/=X`=x�<�U�@Lϼ�`D��u��g����\�ǽϭ���﫽~���7E���Ҽ��?�hP�<i	=*�)=b8=`��<6���3���uH����jK���^��   �   5�Uٿj�.X0�Y�"���Y����)��] ��ѝ��� ��L2��!�������\Y�~�0����8`ٿ.����b��9���FK������꙼��<�f1="�E=N�+=��<��<�qB�4����O�e���<������h=���v���PP�&��x^J���< ��<~h&=:`?="�*=|��<�"��Yֹ��L�E���8!���b��   �   85��:�տ�"
�PZ-���T�~E���F��}D��W����\������D��UU���b���CU���-��Y
���տ�W��k�^��'������G���`U��䖫<2�"=��/=�`=��<�R�Lϼ�`D�zu��`�t���T�ǽ­���﫽s����6E�h�Ҽ �?��P�<Ri	=��)=B9=��<�1��O2��TtH�����J���^��   �   �B���4˿X��&�$�x�I�Plq����,������������������6tq���I�\�$�P��E^˿_S��L�R��
�@穾T�:������⡼@�v<�"�<���<h�Q<�%�F��`Ј�:�Ľ����T��QV�y�#��?����h�����Ľ�/���Y���&� �A<���<8l�<xB]<䱮����&P<�Ur��2�U�R��   �   Yɉ����q�� ���|8�J([���}��������Du��hƗ�����D;}�"�Z��h8�Z���������kC@�V7��
�����(�?���l볼��;�|<@���lϼ4p��ȽT��a9�X�^�%�|��Ї����ض���C|��^�f9��#�:�Ƚfq���Լ W���<`�M;����u����)�J��T���}g@��   �   ��s��N��<qؿ8T�n�#�`�@�]��u�Ӵ��ґ��������t�D�\��@��#�0��Dؿ�.���qs�f�(��ܾ�6���^�​��2ۼ08D�0c���0��ߧ�&�I$B��J��`̞���I�ϾInݾ� �=?ݾ�JϾ�����a�������A� �>��h�2�������S�l伣ԍ����FŅ���ܾ)��   �   �dO�����"����`��p%�,�;�rN�P�Z��>_��Z�NN��X;��%������[��3b��
O�Uk��2���]�q��^i~���(h��m���ͽ'�#�ro�9����Ͼ�s��]K��� �p�*���-�'t*�8w ����~�����ξ{���ܵn�k�#���ͽd&o����V��%���^����^�����+���   �   F~)�'@k��.��Ӗÿս�f4
�f�Du*���3�T7���3�`*�f��
�	�Y��ÿ+К��j��)�8a�����a1�kkʽx�r�,�L�0N���B� �3�ܝ��텼�k���|�0�:���U��#k�:�x��K}��{x���j��JU��:�c�����ջ�c&���w3�0��9���r&N��Eu�R�˽*F2��2���	��   �   p���:�.�w��k��*���O�|�����	�����s�F���q	�����e߿�𾿊��w�x9��$�;�����a�BF�b"����z��%����߽�4�����%�Ⱦً	���2��6]�������L1��#��C&��N����㢿S�����Vx\�I2�'	�@9Ⱦ����l3� �޽&(����{��������b�	����   �   ^bž�g��I=��r�b政� ���(ƿ�(ؿ����o� Z�0�׿G�ſG����i���r���<����.�ľ���\�#���ɽ]$���_��(�ʽ��$�2 ���ež�i��L=���r��蔿w#���+ƿA,ؿ����s��]��׿ѥſ����pl���r�Ш<����ľ����2�#���ɽ�'��X`���ʽ�$�����   �   Ϙ��@�Ⱦ=�	�i�2��2]�������D.��B ���"�������ࢿ;������[s\�2��	��3Ⱦ����f3�!�޽1#���}{���������b�\���,��:�_�w��m������8�������	���v�n���s	�� ��i߿��I����w��{9�k'�O�����a��I�[&��
�z��$����߽$4��   �   ��3��������������%�:��U��k�Űx� F}��ux�6�j��EU��:�N��0��cл�"��q3����Ғ���N�"Bu���˽�G2�4����)��Bk�l0��טÿQ���5
�.�Rw*�:�3��7��3��*������	��쿧ÿ�Қ��j��)��e�<����e1�#pʽ6�r���L�K��'=��   �   ��ͽ&�#�Uko�恢���ϾCm���G��� ��*�^�-��o*��r ����7���7�ξ+���C�n���#���ͽ�o����B������ ���^�¸�C��AfO����������Ba�r%��;�LtN���Z�>A_�ҭZ��N��Z;��	%�~�p�鿒]��8d��JO��m��5����]����Ln~�B���c�B�m��   �   ��0�ا�!��B��F���Ǟ��	��I�Ͼ�gݾ2⾟8ݾtDϾğ��H\�����ަA����4���2�$u����S���㼛Ӎ�׈��Ņ��ܾ�)�߬s��O��xrؿU���#���@��]�.u�$���?�������z�t���\� �@���#�p1�!Gؿ�0���ts���(��
ܾ�8���a������5ۼ�.D��V���   �   �>��`Xϼl�o�I�Ƚ�N�&[9���^��|�:̇�d
��L���;|��}^�
9�$�^�Ƚ(Tq�$�Լ���8< BN;�����t����)�������h@��ɉ�/	��Q�򿜬��}8�~)[�L�}��������v���Ǘ�׉���=}��Z� j8����9����ĉ��E@�u:��+�����(�E���𳼐�;H�<�   �   D��<�R< �~���Ɉ�R�Ľ����H���P���#�,:�Z��?���F�Ľ�'���K�P�&��A<���<x�<�T]<䪮�r���O<�.r��1�n�R��B��)5˿���z�$���I�mq�Ì��-��������������������uq���I�r�$�4���_˿�T��'�R�n�
�#驾��:�����`衼��v<X&�<�   �   ��/=�b=��<��T@ϼ�YD�Uq���a�����ǽd���9꫽m����-E�̒Ҽ�E?�\]�<�n	=(*=== ��<(+���0��TsH�2��VJ�M�^�5��
�տ�"
�JZ-��T��E��/G���D������]��B��OE���U��Uc���DU�r�-�rZ
��տuX��ڛ^�)����G�w����[�����<�"=�   �   �dZ=ҰA=��
=�N�<��w������&��]�恀�Hd�����F�[���#�X���@9X�t��<�=|�@=,�X=<�D=���<2,����.�6��l���&
�"�Q�銕��8ʿ�����#�
wH�F$p�$��-v��7B��+h���C��M���7����p��I�6}$�`���ʿO���nR���
�<Ϩ��7������&#��1�<�bG=�   �   ��E=��%=H��< �;�������h�����~�������䥽M���?f��C�X���о�;|��<2X%=�ED=2P7=܉�<��.�p=��p3�v����.�M�H�����ƿ4� ��2!���D��rk���������q��Oz��Nl��e����1����k�*fE��!�-8��ǿ>~��=�N�����Z��^3�}���(&�dy�<��9=�   �   d�=��<@���0i�bcc�K����ܽ���@��m������ �E.ڽ[����_���ڼ �v���<�2=��=���<�~:��㏽��'��)��
�����B�Ց��(N���[��k�h�:��4^��������z����J��y������m���.K^�< ;������$ͽ� ����wC�G* ��f���'�dE���3�y�<�=�   �   `�;U��~=C�!���Co����&��I��e��Fw��+}��v��d�|H�0%����i �� �?� �����;|%�<0R=<x`[�������H������1����0��cK��l�
v+��J�0�h�����]���B����i���b��&�h��UJ�Rd+�`z�ӂ⿓k��5��@2��X辆�����`�U���A<��<�   �   {�����4��a�.�nXi��8��岪�GϾ�B�˾��Ͼ�6˾F
����������/g���,�����x������� ��-s�h֑���h����>r��3ʾ��� b�Dʚ�<�ɿ?���z���33�*PL��a�~�o�z�t�܅o�r�`��K�H�2�\c�+T��w�ɿU�<b����3ʾ(r������g�<m�� �r���$��   �   �@��:v�W;Y�i����־���美:�l������� ���I�ڂ�O�L��"T����V��������q>���Ѽ�Լ>@Q�^ؽs�H��訾j��?@�ꕄ����u�ڿ��@��.�bW?��gJ�&)N�J�~�>���-����Ԏ���ٿ����sY����?��X�����gH���׽N�P��,ռ|JԼ #A��   �   \m!��u�(������Y��-� kF�[Z��g�54k���f���Y�HkE�v�+�N�#��`y���r�y���X½H?c��!��&F�Zr���B��ᆾVԾخ��[Z��|��ԃ��+-ݿ��Ң�����X'��1*��'�A�����~ �#'ܿ�������Y�v2��Ӿ�t��o���ٮ���E��!���e�>~Ľ�   �   �k|�Z��������~%�ngM���s��Ҋ�����b���%���������%��_r�"L�R$�O��}���Uz�������ֹp���L� >��Ձ��L��o��;_���D,��Jf�`�������Tѿ45�p� �8V���	��� , ���	9п�ɱ��ᑿ�!e�Ao+�J5�������K��L����� M��or���½:h!��   �   �$��$���l/�-�a������W��}�����ɿ�zԿ��׿�Կ=ɿ���m���׉�R`��R.��� �����Hql����ϭ�0Oh�Hi�ꮽ���n� ����i/���a������T��'��� �ɿ�vԿ��׿�Կ	ɿ����j��dՉ��N`�P.�y� �����Mml�8��ͭ�,Ph�8	i��﮽F���n��   �   �d��[H,�2Of�����Ĳ��Wѿ�8�c� �6X��	����- ����;п�˱�u㑿�$e��q+��8�%���0�K�5O�#�����L�fr�<�½�b!�Dd|�D���y��� {%��bM���s�Њ�����_��v"�����}��
#���Zr�RL��N$�s
������Pz�t�����H�p���L��A�������L��s���   �   ���X_Z��~������R0ݿ��̤����*['��3*��'��B����� �x)ܿ����U�2�Y�4�M�ӾLv��Ǹ�Dڮ�x�E���!���e�RuĽ2g!��u��������&V�^�,�)fF��UZ�0�f��.k�i�f�֏Y��fE���+��J����`u���r�H��S½|9c��!�`*F��v���F��䆾CZԾ�   �   6@�Η��=
��4�ڿ,��A�0�.��Y?��iJ��+N�JJ�z�>���-�������ٿ`����Z��^�?��Y�ĩ��`hH�C�׽�P�� ռ@7Լ A�@7���o�B3Y�n����о�����6�`������� ��~���q�/I�$G��P��Y�V�:���𯽢i>���Ѽ��Լ�DQ�
cؽ��H��먾����   �   �b�̚�s�ɿ���
���53�NRL���a��o���t�,�o�t�`���K���2�\d��U����ɿ6Ú�|b����4ʾ'r�0����g�d���Ar���$�ll����8��	�.��Oi��3��R���Nɾ��˾��Ͼ�0˾�������W��Z(g���,����r����h� ��	s�,ّ�څh� ��BBr�7ʾ���   �   ���d2��`M�n�zw+���J�<�h���������n����j��ic����h�WJ�e+��z����-l������2�CY���������U���A<p��<c�; :���,C�����-c����&�h�I���e�T>w�z#}���v�r�d�0uH�*%�����3��,�?���P,�;�,�<PU=<Hi[�Ɗ��u��E��k��1��   �   򒋿�O��u]��l���:�6^��������p����K��H���i����K^�� ;�@��w���cͽ�B����wC�G* ��f����'�!D���2� ��<v=��=�̡<�U���N�
Tc�����ܽ��r;��h������ ��%ڽ�����_���ڼ��t�H��<`6=J�=���<`�:�N揽�'��+��������B��   �    �����ƿ�� �`3!���D��sk�M��:���Nr���z���l�������1����k�8fE��!�8��ǿ~��ܘN�B��cZ��n3�ٛ���&���<>�9= �E=��%=��<�F�;4������h�����y����ॽ����f7f��<�l0�;���<:Z%=�FD=P7= ��<��.��?��`3��������M��   �   q���j9ʿ���#�vwH��$p�Y��Xv��NB��+h���C��#����6���p�"I��|$��_���ʿ����mR��
�8Ψ�"7�~�`#�H6�<�dG=@fZ=(�A=��
=Q�<�w�����&�d�]�����Kd��F����[���#�H����JX�4��<�=�@=��X=n�D=X��<0>,������6��m��^'
��Q��   �   |�����ƿH� ��2!���D��rk����[���Yq���y���k�������0����k�NeE�8�!��7��ǿf}���N����vY��:3�H�����%�t��<�9=|�E=
�%=|��<�G�;��������h�����y����ॽ����L7f��<�8��;4��<�Z%= GD=�P7=���<��.�_>��.3����?����M��   �   �����M��t[���j���:��3^�(����������I��������������I^��:���h����˽��uC��( �e��M�'�0A����2����<�=��=Ρ<@J��pN��Sc�����ܽ��k;��h������ ��%ڽ����l�_� �ڼ��t����<l7=Ȋ=���<hz:�e㏽��'�*�������B��   �   @��-0���J�Nl�Hu+��J���h�����M������\h��Ya���h�,TJ��b+�.y�Ҁ��i�����62��U�V��ی���U� �A<���<0m�;d8��",C�����c����&�Z�I���e�J>w�p#}���v�h�d�&uH�*%�ӆ�� ����?�p���6�;�0�<�b=<�T[�����P�������辄�1��   �   l�a�kɚ��ɿ��������23��NL��a�.�o���t�R�o�
�`���K�n�2��a��Q��<�ɿ����Tb����0ʾlr�n���|g��W��`r��$��j����������.��Oi��3��L���Hɾ��˾��Ͼ�0˾�������N��B(g�y�,�E�뽇q��|��hx � �r��̑�*|h�`���<r��2ʾ���   �   �@�ߔ�������ڿz��>�n�.�fU?�FeJ��&N��J�2�>���-���8���ٿ�����W����?�YV�/���6bH� �׽d�P�hռ�.ԼvA�u6���o�3Y�b����о�����6�\������� ��~��l�#I�G��P��.�V�����ﯽ�f>�@�Ѽ�Լf:Q��Zؽh�H�稾Z���   �   1��\YZ�/{��񁶿�*ݿT�.������V'�f/*�T'��>� ���| ��#ܿ��������-�Y��/���Ӿ�q�����Ү���E���!�<�e�
tĽ�f!�_u��������!V�Z�,�$fF��UZ�,�f��.k�e�f�яY��fE���+��J���Ju��̳r�����Q½>5c��� ��F��n���@�K����SԾ�   �   �[���B,��Gf�{��������Qѿ2쿰� �PT���	���0* �뿮5п�Ʊ��ޑ�oe��k+��/�𡢾��K��C�X���`�L��_r�?�½b!��c|�.���k����z%��bM�{�s�
Њ�����_��t"�����}��#���Zr�LL��N$�b
�����nPz�������ڰp��L��9���|�6�L�Tm���   �   ������Gf/���a�Ϩ��R��=���ɿ�sԿ_�׿�Կ�ɿ[���g���҉��I`�?L.�i� ��ﳾ-fl�����ĭ�Ah��h�$箽����n������i/���a������T��&�����ɿ�vԿ��׿�Կɿ����j��bՉ��N`�P.�p� ������ll�U��5ʭ��Fh�
�h�3宽���� n��   �   �^|����������w%��^M���s�u͊�����\��N������y��  ��7Ur��L��J$��������Hz�X��?	����p�n�L�:��\���L��o��%_���D,��Jf�_�������Tѿ45�p� �6V���	��� , ���9п�ɱ��ᑿ�!e�:o+�.5�¥����K�?J������L�]r�h�½�^!��   �   �b!�`�t�����m���R���,��aF�$QZ��f��)k��f���Y�bE�M�+�G����p����r�����H½()c�l� ��F�o���A��ᆾ�UԾҮ��[Z��|��Ճ��+-ݿ��Ң�����X'��1*��'�A�����~ �"'ܿ�������Y�m2��Ӿ�t��f���֮�b�E���!�r�e��nĽ�   �   �/���j��,Y�T����˾����T3�������b� ��z�u��{�YB�1A��K��%�V����,毽Y>�L�Ѽ��Լ
8Q��[ؽ��H�N訾_��=@�아����w�ڿ��@��.�bW?��gJ�&)N�J�|�>���-����Ҏ���ٿ����tY����?��X�J���NfH��׽�P��ռ�&Լ,
A��   �   >a����������.�@Hi�u/��=����þ��˾g�Ͼ�*˾��������Q���g�.�,�W�� h�� ���M � Ur��Ñ�6zh�����=r��3ʾ��� b�Gʚ�?�ɿC���~���33�*PL��a���o�|�t�܅o�r�`��K�H�2�\c�+T��x�ɿW�<b����3ʾ�r� ��2�g�4Z����q�X�$��   �   ���; %��*C�h{���X����&�k�I���e�6w��}�1�v�6zd��mH�(#%��z�����ڌ?��瀼0��;�@�<@y=<XE[�����@�����l��1�
���0��fK��l�v+��J�2�h�����^���C����i���b��$�h��UJ�Rd+�bz�ւ⿕k��6��=2��X�R��d������U�`�A<��<�   �   >�=�١<@M��:�bGc����۽1��^6�Lc�@���� �8ڽG.�_��ڼ �q�pǢ<p>=`�=`��<@m:�⏽R�'��)�� �����B�֑��+N���[��
k�j�:��4^��������z����J��z������n���.K^�< ;������%ͽ�!����wC�@* ��f����'��C��p�2���<�=�   �   ��E=.�%= ��< k�;���6 ���h�=��u���ۥ����-f�$4��ށ��;���<�_%=VKD=xT7=��< �.��<��>3�i����.�M�J�����ƿ6� ��2!���D��rk���������q��Pz��Nl��f����1����k�*fE��!�-8��ǿ?~��<�N�����Z��(3�Ü���&���<��9=�   �   t�v=\�_=��,=b�<`��;0�,� �ؼ�F��j?�<�I�"g=�.��`�μ�G�(�<Ht�<�1=��b=��x=R�f=�=�V5;N�j�,w�l3��2|��o:�Ʌ�v���F��Z9���2��T��u��߈������<��R������z[u�Z�T��~3�����쿌¶�Ǖ��;�;�/'���S��D��.,n��!;{=�@e=�   �   j�c=�F= F=�l�< ����_ü�))��a��4���燽6��]���#�`K�� p0�u�<��=��I=P.f=�ZZ=�d=@�);\�d����j$����	
7��z������5��H����/��4P��,p�+���n����������M���ap��P��]0��v���N���n7��}#8�\R�P4��"U�"%h��@;�=�tX=�   �   ʡ)=l��<�!<�&f��#�X������ނֽ�)�<���w��$ԽAb���E��t���[J��$9<�<-=R�3=�u=@�:fT�H��RS�����)-���y�v����ܿ�
�*'��8E�~~b�T�{�K���Q����o��X�{�veb�SE�Dq'�$e
��ݿ���]�z��	.�W�6����2IW���:tT =�71=�   �   ���< fu�z�>ه��ѽ{����,�ҚE���U���Z���T���C��W*��(
�z�̽�4��H���"�l�<L�<�׹< `�΀<��;��L|q��˾G��Knd�ST���˿���������4��DN���c�f�r�̾w��Rr��xc�|�M��|4���������̿(����e��H���̾w�r�����F?��GB�t]�<���<�   �   ����L�V��&ý��l�H���|�MI���g�� 鲾ʪ��O���J���Γ�;y���E�X���Ƚ�=N�O��@ K;P�<P���(h#��6ԽO�O�� ���
�wI�@���M���9����	�J� ��E6��H�\�S�rX���S��vG�4�5�R3 ��$	�=]�E���������I�'X
�k��_P��qս��%�� ����; Z�:�   �   �勽��� ::��c��!w��<�̾Ն�U��t����0�������(Mʾ�=���~�P�6�Z{�R������8�=�0<E��9�o6���w*�����辙�*�8+m��T��o�Ŀ����
����&8+�d�4�ν7��04�"�*���n4
�� �|Ŀ�⛿.�l��*����_��l�*��߭�r4���P�$O����   �   ����SS�{L��!nʾ��������0���B��;N���Q�w�M���A��z/��^�������Ǿ���p�O�����̘�2����Ǽ>������)�<i��u����
���B�sy��3!��.Uǿz�连A����"d�x����H�H}��k翃ƿ�4���Ӏ���A��V
�hչ�Wjh�������������ͼV�$������   �   ��Y�'����f�	�-7�mZ���x��X��揿1\��9��������v�J$X��c5�vv���ݾ;�����V�z�K��N-�l��`�S��Ľ��.�q���׾��M�W~��S���Γ����Կ�翬�����1P�@��4�ӿy:��򋟿ه��c9L����־셍��-���ýpS��%�dI0�������   �   �O�l��$�I���x�$���?a�������N���n¿о��˴��E��F����av�I�G�������Z���T�J����a���t&��`'�mԈ�������L�Ƀ��������I��}x�Z���4^�������K���k¿�̾��ȴ�SC�������]v��G�����⾦�����J�����_���u&��e'��و�ڈ����L��   �   Č׾�ΰM��������ݖ����Կ���B��4����S�e��	�ӿ�<���������<L���� ־凍�r�-���ý(pS��!��@0��������Y�����
a�m��(7���Y�>�x��U���㏿SY��v���o�����v�3 X��`5��s�&�ݾ𰟾$�V�w��G���-�n���S� ŽY�.��t���   �   ��
��B��{���#��Xǿ���bC�r��f�`�����I��~�3n翢ƿE6��TՀ���A�+X
�m׹��lh����"������\�ͼ<�$���� ��DLS��G��Lhʾ��������0�8�B��6N�'�Q�֧M�0�A��v/�u[�����I�Ǿ]���O����ǘ�ޅ���Ǽt�����1-�}i�Yy���   �   I�*��.m��V����Ŀ��l�
����:+�n�4�Կ7��24�ԅ*�f��5
���!Ŀ 䛿�l���*���羅����*�0୽D2���P�O���܋�R���2:�_���q���̾�������T��������|���Gʾ9��ȩ~���6��r�`���������=��<E��=��:��c{*�c�����   �   �yI�車�P������\�	��� ��G6��H�vT��X���S�NxG���5�p4 ��%	��^�Y�����ըI��X
�gl���_P�rս$�%�P��� U�; ��:�n���V��ýh����H���|�ED��sb��l㲾5����I���E��[ʓ�63y��E���l���f0N��=��@vK;��<ൎ��l#�q;Խ�O�t��� 
��   �   �pd��U����˿���������4��FN���c�^�r���w��Tr�lzc���M��}4�H������m̿�����e�CI�1�̾��r�����D?� gA��g�<��<,ъ<��t����χ�"yѽ:���,�j�E�LyU��Z�Y�T���C��Q*��#
�Ry̽-������@��x�<�<dٹ< R�؅<�@���q���˾���   �   ��y��	���ܿ�
�+'��9E��b���{�������Fp��p�{�Lfb��SE��q'�je
�v�ݿG�����z��	.�W��5��d��FW���:tX =�<1=d�)=���<8�!<��e��#�s���󧲽�yֽp ��w��S�뽤�ӽ�Z��?��2y�`7J�8A9<P�<z-=��3=�u=���:d$T�X���T��+�P+-��   �   E{������G�����p�/�f5P�z-p�����爏�>��N������bp��P��]0��v�q�'���B7��&#8��Q��3��LT�"h��n;�=�wX=N�c= F=hK= y�<�|��Pü6!)��a�60��nㇽ���@]���#�T?��  0��|�<��=��I=H/f=�ZZ=^c=`�);ضd�n���%�����>7��   �   }Ʌ�����뿮9�:�2�@T��u���������<��?������"[u���T�2~3�>��z������M���r�;��%���R�����h(n��N;:}=tBe=�v=��_=�,=d�<0��;��,�̘ؼF��j?�H�I�dg=����ȴμ�K��<r�<�1=L�b=X�x=��f=�=�*5;�j�zx�S4��j}�p:��   �   �z��ʽ��V��P����/�p4P�D,p��������j������ ���`p��P�.]0�"v�w �`����6��D"8��P��2��3S�@h���;�=�xX=ƥc=hF=�K=dy�< |���Oü2!)��a�10��kㇽ���4]���#�@?�� 0�$}�<��=ޚI=�/f=`[Z=�d=��);�d�[���$�����b
7��   �   Åy�E��O�ܿ�
��)'�,8E��}b�D�{����������n��Ɗ{�db��QE�8p'�@d
���ݿ̸��U�z�.��T�X4��O��AW���:�Z =J>1=8�)=���<p�!<��e��#�e���槲��yֽi �w��K�뽙�ӽ�Z���>���x�X6J��B9<x�<T-=B�3=�w=@-�:T�L��XS���ᾭ)-��   �   �md��S��)�˿���������4��CN�d�c���r��w��Pr�wc���M�H{4�R��Y����̿�����e��F��̾��r�
��t=?� 5@� n�<p	�<tӊ<��t�����χ�yѽ0���,�b�E�HyU��Z�T�T���C��Q*��#
�5y̽�,���������Tz�<�"�<d߹< ���~<�i:���{q���˾Ҹ��   �   �uI�|���E����� �	�4� ��D6�BH�v�S�`	X���S��tG�b�5��1 ��#	��Z�?���H����I�&V
��h���ZP�5kսD�%��ѣ�Pr�;���:Xl��:�V��ýR��z�H�|�|�DD��qb��j㲾2����I���E��Vʓ�*3y���E�ܽ�&����/N��:�� �K; �<����0d#��4Խ�O�����9
��   �   >�*�W)m��S����Ŀ��
�h��v6+�~�4�Ȼ7��.4�*�*� ��2
�����Ŀ������l�i�*����a����*��ح��(���P�8�N����'܋�����2:�
_���q���̾�������Q��������t���Gʾ�8����~���6�|r��������=�h$E�D4��3���u*�N����   �   }�
���B�x��}��Sǿ���*@����Rb����� �6F��{�zh翦ƿ2���р�;�A�T
�yѹ��dh�@������Χ���ͼL�$�m~�����LS��G��Chʾ����
����0�5�B��6N�$�Q�ҧM�-�A��v/�p[�����;�ǾK����O�����Ƙ����(�Ǽ��;����'�Li�ts���   �   �׾��/�M��|��9���T�����Կ���D������L�����ӿm7��9������y5L���־J�����-�P�ý�aS����:0�����]����Y�~���a�j��(7���Y�<�x��U���㏿RY��u���n�����v�0 X�|`5��s��ݾڰ����V�}v��E��
-�4����S���Ľ��.��n���   �   ���� 
�i����I��yx�����[�������H��uh¿�ɾ��Ŵ�L@��.����Xv���G������d���I�J�����W���g&�X'��ш� ����L�����������I��}x�Z���5^�������K���k¿�̾��ȴ�RC��􉑿�]v��G�����⾄���C�J����]��Vm&��X'��ψ��z����L��   �   �Y�2����\྘�W%7�y�Y���x�)S������sV������������v�aX�@\5�p�A�ݾG�����V��q��>���-����S���Ľ�.��p���׾���M�X~��S���ϓ����Կ�翫�����0P�?��2�ӿw:������؇��a9L����־����`�-�l�ý�hS����80�X���J���   �   ؎��FS�D���cʾ#��������0���B�<2N�U�Q��M���A��r/�~W����r�Ǿ���{�O��������v���Ǽ�������(��i�qu����
���B�vy��5!��0Uǿ}�迠A����$d�x����H�H}��k翁ƿ�4���Ӏ���A��V
�Gչ��ih������������ͼ�$�vy���   �   2֋�_���,:�`[��8m���{̾�y�?�� �����������z뾩Aʾ�3�� ~�C�6�g���������8�=� E�2�4���v*�l���辚�*�=+m��T��s�Ŀ����
����*8+�f�4�н7��04� �*���n4
�� �}Ŀ�⛿.�l��*����,����*�@ݭ��,�p�P���N����   �   �Z����V�@ý�����H��~|��?��a]��޲�����D�� @��Wœ�$*y�"}E�F��\���zN�� ���5L; �<pg��bb#�5ԽʧO�� ���
�wI�D���R���?����	�N� ��E6��H�`�S�tX���S��vG�6�5�R3 ��$	�?]�G���������I� X
�\k��~^P��oս�%��ڣ�p��;���:�   �   pߊ<�t����<ȇ��oѽ����y,�o�E��qU�c�Z���T�z�C��J*�H
�Mn̽�#��h������h��<L1�<��< *��|<�J:���{q��˾F��Pnd�UT���˿���������4��DN���c�h�r�оw��Rr��xc�~�M��|4���������̿+����e��H���̾�r�����B?���@��o�<<�<�   �   ��)=���<��!<��e�\�"���$���	qֽ@�An�����b�ӽ�Q��7��k��J��j9<�*�<�-=\�3=�{=���:�T����8S�����)-���y�y����ܿ�
�
*'��8E��~b�X�{�M���S����o��X�{�xeb�SE�Fq'�$e
��ݿ���^�z��	.�W��5��h�xFW� ��:bZ =�?1=�   �   Ȧc=pF=�N=h��< T���Cü)��
a��+���އ�J��$]���#�d/����/����<D�=r�I=�3f=�^Z=vg=@�);�d����_$����	
7��z������7��H����/��4P��,p�,���o����������M���ap��P��]0��v���O���n7��|#8�WR�C4���T��#h�@a;֨=�xX=�   �   ��=���=�CU=RY=�D�< �; s�86�� .⼘���ܼ�ɞ�p( ����;��<�� =��\=�=��=O��=`M=�;�<���:��Rp�A�̾|���&f�W^����̿ ������5�n�O���e��t��Uz�\�t��e�B�O�h,6�M�h� �T*ο�z��h�g�-c �c#Ͼp�s�x��(m��<��G=�D�=�   �   �n�=-l=�)8=���<�',<P|軈���t����-���7���*�D	����𜢻�P<�X�<`R@=�[s=L��=�R�=f�F=8��<��	�M���k�8�Ⱦ���8b�彚���ɿ����`/���2�:�K�>Va�p��7u�.�o��Za���K� �2�ִ��#��`�ʿG��c�7W���ʾE7n�̳��*�$��<TqA=�}=�   �   X�R=*O&=�R�<���:�~��
�1�_[��?���Zഽ���� �����<�y�Ns'�����	�;�N�<��.=
�Y=��_=��3=�_�<(��a|ֽ �[�(����d�YV��������3�@����)��$A���T�l*b��f��b���T�2A���)��?����T����ؓ�ϮW���D���̅^�6�ڽ0t�|v�<�2.=��Y=�   �   ���<h_7<�(k�^�5�����E;۽��	�0���y-���1��^,�F��&��+�Խ�K��N�(�ؠ<�hz_<P�=Z�#=�=�x{<l�μ ���HD�a��������C�U���谿�ݿ ���Y��1�>PB���M�ܶQ��}M��A���0���,����ݿA���r��6�D����ҫ�/bF�Q���Lۼ0Jd<��= �=�   �   �� �6����.��LW"�)�O�A�w�����磕�-Ԙ��ꔾVP���#t��nK����߽�ˇ�T��  j���<��<p�:<<v������&��W����龷T,��o�<x��ƿn������8.,�`�5��8��R5�"�+��������ſ0^���>o�4�,�b��P���](�N����ͮ��$<��<�ʄ<�   �   <_<�����:[�Y�T�����<��b�Ⱦkc߾P���E�?��.�ݾzpƾ�`������O���Н����0���?��t�;@��;T߂���t����I�r�u�þ����K��$��C��BϿ���L��r�Z;����������Ċ�u��V+ο�0��v���kJK��i��þU@s��f�hx�(G�� �I;�_Q;�d��   �   T�ѽ�B+��{��(����ؾe��6�)�&���0�%�3�20�J�%�%���O��jվQ��r�u�D�&�˽*�O������ݻX:i��85�ѫ̽��=��᛾���٠&�R_���c*��`�ʿǜ��������2��\m��������:ɿ)櫿�����]��%�4i꾆I��4E=��̽F�6�h v�X������l�Y��   �   >�0������F��������&;�=V�G k��\x�ƞ|�[�w�ģi�Y-T�9�E��Z{��>F���1���e-��̽�QP�.���)��� ��7��6�
��6k�V\��8��G0��b�&��V���*����ɿ�PԿ�׿Z�ӿȸȿfȷ�HD��։�\�`�E�.����̳��8i�4�	�2>���6 ����<�¼FYW��ѽ�   �   b����G��<����,���U�#r}���2���!���q����z��s����⎿x�z��S�]�*�7�nӾ�
�����"�|!��J�3�`���4���&7��8���g%�Ʒ���B��3��Ѻ,�/�U�:m}�n��^���=������� x������A���d�z���S���*��4�о���s�"���� �3�،������B/7��?���l%��   �   w`���:�gK0�>�b����	���l-����ɿ�SԿ��׿T�ӿ��ȿ�ʷ�xF���׉�f�`���.���ϳ�><i�M�	�/@���6 �����,�¼*MW�Q�ѽ0�0������A��o��(���";��V�Uk��Wx���|�}�w�:�i�?)T�m9�>��qv��hB���.��za-�~~̽�KP��)���,��� �=��Z�
��<k��   �   ~��ɣ&��_�6���,��1�ʿן�.���L������n�r�����*=ɿ	諿S���]�ܺ%��k�HK��^G=�@�̽��6� v�Pn�$뭼$�Y���ѽ`<+�}{��#��ѽؾ���b��&�u�0���3�$0���%�����L��eվD�� �u���&�J˽`�O�p����ݻHEi��?5�̱̽/�=�3图�   �   5����K�u&��u�~EϿq��N�<t�
=�������>�������-ο2������LK�/k���þXBs��g�Px�4C����I;��Q;h�c��O<����T�|�T�O������l�Ⱦ]߾���@?���@�ݾ!kƾA\��������O�"��f���2�0��k?�`��;���;�悼��t�"���r��þ�   �   W,��"o�z��!ƿep�:��$���/,��5���8�T5�z�+���������ſ$_��N@o�7�,������o^(�����lʮ��$<��<0܄<@�� �6������dP"�?�O�|�w�����QϘ�'放�K���t��gK���zz߽xć���� ��6<��<��<`�:<�~����'�BZ�����   �   �C��	��]갿��ݿ���Z��1��QB�X�M�Z�Q�M�<�A���0�L������ݿ�A��as���D����ҫ��bF�3����ۼ�Vd<V�=��=��<��7<��j��5�*�L0۽��	����0s-�B�1�`X,�>�������Խ�C��.�(��w<�8�_<��=V�#=�=r{<0�μ���KD�����$���   �   �ZV�������W5�����)�&A���T��+b�B�f��b���T��A���)��?�U�����
ٓ��W���E�����^���ڽ r� |�<H6.=:�Y=B�R=zV&=�d�<�+�:4f���1��S��$���ش�������������y��g'� 薼 J�;4[�<"�.=�Y=��_=��3=`[�<�0���ֽ��[� ���If��   �   �b�������ɿ�����/�\�2���K� Wa��p�H8u���o��Za���K� �2����#��H�ʿ%���c��V�h�ʾf6n�T��6(�$��<tA=�}=�p�=01l=~.8=���<(A,<D�h��������-��7��*�Z	�����pr����P<�_�<�T@=�]s=���=�R�=Z�F=���<��	�P��
k���Ⱦ����   �   x'f��^��C�̿f �����5���O���e�$�t��Uz�@�t���e� �O�,6��L� � ��)ο8z����g�}b �S"Ͼܨs�)���i��
�<��G=rE�=��=P��=�DU=@Z=�F�<@�;�p�d5���-⼬��t�ܼ�ʞ��* �@��;8��<�� =��\={�=�=���=�	M=�6�<���~��Sp�Q�̾,���   �   �b����ǚɿ����\/���2��K��Ua��p�7u�t�o��Ya���K�T�2�:���"��l�ʿu�����c�'V�S�ʾ�4n�c�콲%�`��<uA=f	}=�p�=b1l=�.8=,��<�A,<�C�X��������-��7��*�X	�����Pr����P<�_�<U@=�]s=���=S�=T�F=���<�	�p�罖k���Ⱦ&���   �   �XV�o��]��i3����h�)�J$A���T�l)b���f�bb�v�T�A���)��>�Q������ד��W�3~�8���Ԃ^�ؽڽ^m���<@8.=r�Y=��R=�V&=�d�< 1�:�e��
�1��S��&��� ش�������������y�~g'��疼PL�;�[�<��.=��Y=8�_=t�3=Xa�<x'��f|ֽ+�[�!����d��   �   Q�C����(谿I�ݿr���X��1�OB�z�M�`�Q�.|M���A�4�0�N�����ݿt?���q���D����ϫ��^F�!����ۼ�gd<�=X�=��<Ѝ7<��j���5��B0۽��	����0s-�A�1�\X,�:�������Խ�C����(� v<���_<��=�#=J=��{<h�μ��8HD�〉�*���   �   �S,�Uo�Vw���ƿ�l��������,,�ޮ5�|�8��P5���+�:�������f�ſe\���;o��,��꾾���Y(���������X�$<��<��<���R����d��ZP"�<�O�}�w�����RϘ�'放�K���t��gK���[z߽Eć���� �7$��<��<`	;<o������&��V��S���   �   ���J�K��#���謹CAϿ���ZK�0q��9�:��B��,��8������(οr.������bGK��g�T~þ;s��b�8x�2�� %J;�R;�c��N<�B򹽻T�l�T�L������m�Ⱦ]߾���??���>�ݾkƾ<\��������O�������0�Pc?�p��;@��;�Ղ�Ьt�Q���r�σþ�   �   g���&��_�����(��0�ʿ@�����������k�`�����"8ɿ�㫿����]��%��d�F��@=�Z�̽��6�X�u��W�8䭼�Y��ѽ;<+�l{��#��нؾ���b��&�w�0���3�$0���%�����L��eվ<���u�^�&��˽L�O�����0�ܻH#i��25��̽�=�����   �   �Y��J6��E0��b�N��+���(����ɿ�MԿȪ׿9�ӿ��ȿ}ŷ��A���Ӊ�9�`�׬.���ȳ�p2i�n�	��6��$* �P�����¼�IW�`�ѽ��0������A��p��*���";��V�Xk��Wx���|�}�w�:�i�<)T�k9�;��jv��^B���.��2a-��}̽hHP�8����������3����
��2k��   �   V���m?�� ���,���U�&i}���˄��z�������u������ݎ���z�?�S�ٵ*��1�K˾����"���4�3�4t��$���V!7�E7��"g%������B��4��Ժ,�4�U�@m}�q��a���?������� x��ᘜ�A���d�z���S���*��4�о����"�J��`�3��}������D7��3��d%��   �   ��0������=���	����;�vV��k��Rx���|�l�w�K�i��$T�4
9����*p��H=���*��.[-��t̽N<P�$��T�������5����
�`6k�H\��8��G0�!�b�)��[����*����ɿ�PԿ�׿[�ӿȸȿgȷ�ID��։�Z�`�C�.����̳�t8i���	�"<��&0 �脆�l�¼�CW� �ѽ�   �   :�ѽ|7+�{����ȸؾ�����D�&�e�0���3��0�n�%���II��_վ2��׼u���&��˽�O��v��P�ܻpi��35�$�̽$�=��᛾���ܠ&�X_�
��i*��e�ʿΜ��������4��\m��������:ɿ)櫿�����]��%�&i�fI���D=�g�̽��6���u�0T��ڭ�T�Y��   �   D<��깽�O��T�Z���+���	�ȾW߾T��8�J���ݾ0eƾ�V�������O���������~0�86?�@�; �;�т���t�L����r�f�þ����K��$��I�CϿ���L��r�^;����������Ċ�u��X+ο�0��v���lJK��i�΁þ�?s�5f�
x�l9���#J; HR;(�c��   �   `9�����؅�~J"�H�O���w�����V���vʘ�LᔾFG��>t�`K�
��n߽Ⱥ��hl� �7l�<�(�<x;<�k��^��O�&��W����龼T,��o�Ax��ƿ	n������>.,�d�5�$�8��R5�"�+��������ſ1^���>o�6�,�U��0��(](�����î�X�$<h	�<��<�   �   ���<p�7<��j�^�5��꛽�&۽ �	�����l-���1��Q,�Ł������ԽG:����(�@<�@�_<0�=x�#=�=؎{<�μ���HD�P��������C�Y���谿%�ݿ���Y��1�DPB���M��Q��}M��A���0���,����ݿA���r��7�D����ҫ��aF�%����ۼad<��=b�=�   �   
�R=�[&=�q�<�9�:�Q��,�1��L����ϴ�D�����������y��Y'�xϖ����;dm�<�.=�Z=��_=�3=�f�<P#���{ֽ��[�����d�YV��������3�D����)��$A���T�r*b��f��b���T�4A���)��?����U����ؓ�ϮW���8�����^�|�ڽ�q��}�<�7.=��Y=�   �   >q�=43l=@18=X��<HS,<��ĥ������-��7���*�\	�����0:���P<�j�<�Y@=�as=���=�T�=��F=ԭ�<��	���罴k�4�Ⱦ���:b�罚���ɿ����d/���2�>�K�@Va�"p��7u�0�o��Za���K��2�ش��#��`�ʿI��c�8W���ʾ27n�q�콜)����<�sA=`	}=�   �   �=\��=ȋ�=�K=^�=�n�<x$<�aR��߻���WĻ zB:��3<�<��=F�V=~�=���=��=n��=��~=�=�3�҈����8��壾p����=�H���ȫ�oX׿�����n�+� X<�||G�ZkK�&}G��i<�l�+�
�6o��~ؿ�﬿8��h�?�z��k��h=���� �^���=�Iv=�R�=�   �   hz�=���=��g=
�,=|��<��6<�!��$T�$ş��ׯ�d����9� j<�@�a<�;�<�}8=�r=ݏ=2�=���=�y=�L= �"� p���4�w{���*��r~:��Ѐ������ӿ�����?���(�b9���C�r�G�&�C��9���(����N �~�Կ\���ʁ��6<��� ��ߢ��o8�H�����L��=t�p=�F�=�   �   p�=4�X=��=��< �7�����*���<N��+p�vz��l��F�\]��H�� Y%;�m�<'=��c=-�=y�=��h=�/
=�t��ܐ���'�͔��3�ﾏ�0�ړt��Ǡ�9�ɿ��9�z� ��/�R�9��#=�ʏ9�*�/�� ��H�'I����ʿ��v�R�1�>%�'���2+�ω������8=D�_=`ׂ=�   �   R�1=�]�< �;\ڨ��HD�Q��!4Ƚ7��Z�_��A���� ���zܐ��~4�(����i<�?�<��<=nAZ=R�J=��=@F���u�(��-��P;پ�� ��`��ݓ��F��o>ῄS����!�8]*��Y-��#*�.9!���@��Όi��	/���`�q�!���ھ���L�����Ǩ����<X�A=�XP=�   �   ��<�[!��l-�Zx��*��D@�xEA���[��l���q�k��X�H=����!���H�P�ʻH^�<��=�4=�*�<@s�:@� ?����g�������#�E��?��-���^ɿ�뿶a��&����6�Xg�$������꿮�ȿ����&��N�E��j�)����Si�5���P@G��� �P;�<�'=N�=�   �   ����Șv��`۽f�#�^�[��6��bq���q���k��3ľk��P���|�X��!�U����mLѽhe������
<<@�<x��< 6�;v{�E���<�����(�o�'��f`�"ӎ�a𭿙~˿�f� ����8�dN����%�����@ʿ.﬿���_�NV'�E��z�����<��ýBh� E;8�<@ �< z�;�   �   Q����6 �&�C�	����ܮ���Ծu�����H�M���]��w����rѾN���B���>����D函�Wμ 8�:P�H<�]�;q��4����n��tv��U��Ij��68��Ml��������1+��$Tѿ�ܿ>�߿�tۿ%2п�˾�������[lj���6�����?��4Xu����ک����;8'/<��5�����   �   ��`�R�������ʾ[ �����0���B�h�M��OQ���L��A���.����<��hǾ�q����M�j�5���,�Ѽ�]غ@e�;�����.�**ɽ�6��А��xӾߣ��Y;�Fg�������5G���5��f������%>������"J��%�d��H9���X Ѿl5���4�6�ƽ-����w^; �@�����y���   �   �N�9󚾖�׾
���0�}*R��o��Y��g���'܌�����u�� nm� �O�A.�����Ծ�^��GKJ�_�2&p�����.i� ۚ�������v�G���N�6w�׾��m�0�N&R�{�o�WW��팊��ٌ����Qs��jm���O�>.� ��*�Ծ\��HGJ���p�t�� Ti�@\������4�v��O���   �   _Ԑ�}Ӿæ�)];�'Jg�a������I��D8��������@������L��Q�d�.K9��
�e#Ѿ�7���	4���ƽx-������^;�~@����jr�������R�5���b�ʾ8 ������0�}�B��M�MKQ�p�L��
A�j�.���� ��BǾ�n���M�������t�Ѽ� غ�Y�;�����.�.1ɽ�6��   �   QY���l�:8��Ql������-���Vѿzܿ��߿wۿ�4п�;�ӱ��5����nj���6�O���A��0[u���x�<۩��Ǘ; </< �3���򁏽1 �0�C������׮���Ծ��������������Z��t�ڢ�mѾ�I���?��r�=�����߇�xHμ���: �H<�K�;�|��E���tr�(zv��   �   �,���'��i`�Վ�����˿i�إ��:��O�F���������Aʿ��U����_��W'�V��ޕ����<�Fý�h��6E;h#�<�-�<@Ⱥ;ڲ���v��U۽��#�z�[�w2��`l���l��(f��y-ľ�e��R����鞾�T����U�(��DѽV[e�h���P�
<F�<���<��;�������<�~����   �   ����E�1A������`ɿ���b�4(�H��L7��h�:�����}���ȿ+����'����E�[k�H���$Ui������@G� E ��A�<�,=�=X�<�&!��\-�in��t��9�>A��[�ԟl���q�(k���X�hA=����-��� <���ʻ�k�<�=�6=$)�<��:�	@��D����g������   �   �� ��`��ޓ�DH��8@ῂT�.���!�b^*�[-��$*�:!��������j���/����`��!���ھ~�������������<|�A= ^P=ڭ1=�p�< d�;$���p8D��G���)ȽB��y���<�y�轿���bԐ��p4�������<@M�<��<=DZ=�J=��=�MF���u��*��/���=پ�   �   �0���t��Ƞ��ɿ����9�V� ��/�:�9��$=���9�Ώ/�l� ��H��I���ʿ7����v���1�f%�*����1+�.������:;=n�_=hق=��=��X=`�=(1�<�!5��磼0��$/N��p�hz�Tl�H�F��Q��4��`�%;�{�<�	'=��c=}�=�y�=N�h=0.
=����ߐ���'�t���y���   �   �:��р�[���e�ӿ����.@�|�(��9�B�C��G���C��9���(����N �y�ԿH��lʁ��6<�l� �{ߢ��n8������L��=��p=H�=�{�=[��=��g=��,=h�<�6<��H	T�D���ʯ�|���Pk9� 7�P�a<XC�<��8=Z�r=�ݏ=~2�=���=�y=�J=@�"��r��ď4��|��d,���   �   ��=����	ɫ��X׿>��Ȯ���+�(X<��|G�ZkK�}G��i<�:�+����n�f~ؿ+﬿�����?����j��=������^���=�Kv=�S�=��=ڲ�=>��=إK=�=p�<�&<�KR� ߻ ��PYĻ `B:X�3<�
�<��=|�V=�=5��=���=ѩ�=*�~=�=(�3�����R�8��棾���   �   �~:��Ѐ�������ӿ�����?���(�"9�^�C���G���C�9��(����M ���Կ����Ɂ��5<�ň ��ޢ��m8�`�����L�P=��p=`H�=|�=t��=��g=��,=��<�6<���p	T�d���ʯ�����`k9� 7�p�a<hC�<�8=t�r=�ݏ=�2�=ұ�=�y=L=�"�q����4��{��$+���   �   k�0���t��Ǡ���ɿ���8�� �j�/���9��"=��9�B�/�� ��G��G��4�ʿЁ���v���1��"�n���/+���� ���== �_=�ق=0�=��X=��=T1�<�5��磼.��:/N��p�hz�`l�D�F��Q��4�� �%;�{�<�	'=J�c=��=?z�=��h=�0
=�r��ܐ���'�ɔ�����   �   n� ��`�ݓ��E���=��R�b���!�6\*��X-��"*�
8!���@���h���-����`���!�4�ھ���\���~�0���h��<��A=�_P=��1=hq�<�e�;Խ��Z8D��G���)ȽI��y���<�y�载���WԐ��p4�@�����<TN�<��<=~EZ=V�J=�= �E�6�u�~'�|-���:پ�   �   ���E��>��.��`]ɿ� ��`��%�Ȳ��4�
f�ڦ�����꿢�ȿQ���M%����E��h�6���qOi������6G� ���J�<�/=�=X�<�$!�>\-�Wn��u��9�>A��[�ݟl���q�/k���X�hA=���� �����;� �ʻ�m�<��=L9=�1�<@֜:��?�=��)�g������   �   �&��'��d`��ю���|˿d�Р��d7�
M����n~�� 俶=ʿ�5��؁_��S'�I��|�����<��
ý�]��E;-�<�3�< ׺;ز�
�v��U۽��#�}�[�{2��fl���l��.f��|-ľ�e��U����鞾�T����U����Cѽ�Ze�4�����
< L�<ش�<PW�;w�����<�;~���   �   _S���h��48�TKl�������)���Qѿܿ��߿�qۿn/пɾ�����q����hj���6�C���;��kRu���銽lĩ���;`O/<�3����}����0 �'�C������׮���Ծ
���������ä��Z��t�ۢ�mѾ�I���?��^�=������އ��Dμ��: �H<���;xf��}��ml��qv��   �   �ΐ��uӾ��W;��Bg�:������D��3�����枱��;������G���d�E9����Ѿ�1��x4��ƽH-��X��_; 5@�<�἟q�������R�7���g�ʾ< ������0���B��M�SKQ�t�L��
A�l�.������?Ǿ�n����M�������ȔѼ@�׺��;����.��%ɽ�6��   �   �	N�l욾��׾�����0��"R���o�&U������A׌����p��zem�^�O�i:.����Ծ�W��AJ�g���p�p��� �f� 	��������v�uF��xN�4�׾��v�0�X&R���o�]W��򌊿�ٌ����Ts��	jm���O�>.� ��&�Ծ�[��GJ�B�6p�@�� �g����p���*�v�'A���   �   ,����R�����?�ʾ� �|��&�0��B���M�GQ�"�L��A�~�.�R������Ǿbj��@�M���F���(�Ѽ@�ֺp��;���$�.�$)ɽ�6��А��xӾ���Y;�Fg�������=G���5��m������'>������#J��'�d��H9���Q Ѿ[5���4�#�ƽp
-�hm��_;�@����	m���   �   �{���, �ʾC�P���RӮ���Ծ=���^��K��3��W�Kq�o��gѾ�D��J;��u�=�տ���և�t,μ )�:�I< ��;pg���~��2n�xtv��U��Oj��68��Ml��������;+��-Tѿ�ܿE�߿�tۿ)2п�˾������]lj���6�����?���Wu�h�)�Щ�P�;�R/<�2�����   �   �Ų�<zv�DM۽P�#���[��.���g���g���`���'ľ0`������ 垾=P����U����9ѽ�Ie���X�
<\Y�<��<Pe�;�w�%��X<�����(�w�'��f`�)ӎ�j𭿣~˿�f�,����8�hN� ��)�����@ʿ/﬿���_�NV'�@��h�����<�`ýld� {E;�,�<�9�<��;�   �   ��<� �bO-�4f�����3�`7A���[��l���q�k���X�:=������(���+� ʻ聙<
�=�>=48�<��:0 @�R>��p�g�������+�E��?��5���^ɿ�뿾a��&� ��6�^g�(������꿰�ȿ����&��Q�E��j�����Si�^���t=G� v�$I�<X1=�=�   �   \�1=�<���; ���t*D��?��� Ƚ�~�:t��n6���轊���ː��`4�x��� �<0a�<�==KZ=f�J=��= �E���u��'��-��P;پ�� ��`��ݓ��F��z>ῊS�"���!�@]*��Y-��#*�29!���B��Ὼi��/���`�q�!���ھ������� ������<��A=@bP=�   �   �="�X=,�=�?�<��2�Hӣ����^"N��p��Yz�4l�zxF��D�(����&;�<n'=��c=U�=6|�=�h=3
= d�Wܐ���'�Ŕ��4�ﾔ�0��t��Ǡ�?�ɿ��9��� �
�/�X�9��#=�Ώ9�.�/�� ��H�+I����ʿ򂡿�v�S�1�:%�����1+�/���8��<=��_=�ڂ=�   �   }|�=<��=N�g=��,=,
�<��6<@c�H�S�\���|�������P9� �0���a<HN�<Ѕ8=��r=�ߏ=&4�=��=.�y=8N=�"��o��֍4�t{���*��t~:��Ѐ�������ӿ�����?���(�d9���C�v�G�(�C��9���(����N �~�Կ]���ʁ��6<��� ��ߢ�po8�����x�L�X=��p=`H�=�   �   ��=��=-Ŗ=2�=��M=\V=���<p��<�}j<p
S<8Wy<�Ԭ<���<:%(=�sZ={��=�F�=�J�=��=
5�=�Z�=�}Q=�R<&P7�$O���v�
ɾ2��1QQ�w��۶���pӿ������
�Ɖ�$��ƞ"�<��Ɠ�L�����3Կ�����n��3S�L���̾7&|�&��bF���<V�E=t��=Ē�=�   �   ���=M��=��=Ʒe=�.=��<��<�C< �t; �;�N�;��4<�#�<p�= \<=$vs=���=���=괯=��=9�=�P=`�`<r/�>{��kq��ž��,�M�"���૿п`����*������F�t������/�пۭ�����[O������Ǿ�bv����`�=�(i-<�D=�b�=9A�=�   �   �i�=�̅=��V=R=���<��k;�<0�<<��`�� �����d����3���;���<>n%=fe=���=겜=��=?��=8�M=�<�\�O��Yoa�HZ����
���B�dU��
���gSƿ8l�4_���r���!��u���L�}|�8�ƿ���1��1D�y<�����s�e�=V𽄍$��wV<�lB= �=��=�   �   \�j=TQ3=,��<@�[;͟�\R*�(�y�^훽}-���鴽,��������_l�<?���z�0f�;��<V_B=�;x=�q�=�ځ=��F= `�<�缨�Ƚ�H� ��M����2��Bm�����}�׼տ������	� 6��	����+O�q^տ�ж�����<�m�$�2�	+���Ψ�X�K�B�ν�S����<�J<=�x=�`�=�   �   �
=H�L<Ѝp�&F:�|ў�q1޽q��� �؅.���2���,������f�Խ��&�hZ%���<�p=J�N=��\=Դ9=�o�<0%��$"��Q)�2����/ܾu�%�Q�Hƅ�#������s׿��R�������V#��R��u�ֿ�B��Е���w����Q�����ܾ㐾V+�X���r��`�<�/=v�Q=�aB=�   �   `w";4��b	�����x� �DUM���t��剾����	�������l	���o���G�0��:8ٽ�U��xE̼��;���<P�%=.*#=���<��л�j�R����k�������Yk2�le�:U���礿"b��M˿G�տ��ؿjտ�&ʿ�M���ۣ��u��b�c�ڛ1�,��F\��pl�4��@�n�؎ �t]�< u=z�=���<�   �   W���������}J�uN��)[�� 㿾orվ� �A?���ᾃ+Ӿ
׼��㠾b���C����l��0�	� �9�P�<�� =��<�>�;ȯ���½��5�ϝ��;�Ծ�z�G<�7<h�h��$|��6�������Z����"���ʨ�PR��\쇿f�5�:�7�| Ӿ����4�9J½�$�`O];T��< f�<0x�<�4��   �   )U��	0�A�d�����Ǿ���'j�-��E##�e&�Wf"������	�-��þ�`���:^�u��F$��H � ����r�<4��<�]W<؄r��y�NI��;Y�~𢾗[���X+8���Z��=y�"r��:ۏ��8��`\��䌇�N�v�
gX���5��*��K߾ƪ���V�>���.�t�0�l�HPS<�1�<0��< ���G��   �   ����i�������ݾ�Q���&�a?��R���]�ųa�p]��qP�=	=���$�	��پLk���d�F���������0�;ඣ<85�<@�U;���_�����V�i�x���r�ݾ�N�(�&��?��R���]���a��
]�<nP��=���$��	���پ@h��x�d��B��������C�;�<�.�< �U;�������   �   �AY�6���M`����.8���Z��Ay�Qt��uݏ��:��}^��ݎ����v�%jX�D�5��,�O߾D���ZV�����t���l��OS<�6�<���<@D�X;��L���*�<�d�:���ǾǏ��f�����#��&��b"����͘	�7��{þl]��t5^�y�������� �|�,v�<���< MW<��r�x"y�lM��   �   ᠑�A�Ծ-}�'J<��?h�h��N~��z���������$���̨�T���퇿�f�`�:��8�#Ӿї����4�EM½�'� G];$��<�n�<h��< 4�,I��w��7���vJ�PJ��kV���ݿ��lվ���x9�b��N&Ӿ\Ҽ��ߠ�����+�C�>��pe����	� H�9�W�<�� =\��<P�;��K�½j�5��   �   פ�����m2��e�W���餿Gd���˿��տ �ؿ�տ�(ʿDO��Oݣ�!w��n�c�s�1�^���]���l���� �n�H� �h`�<�x=0�=	�< (#;�i�i ����� ��MM�o�t�;ቾ&�������>���\����o�9~G�ʖ�k/ٽ�N��X0̼���;h��<ƍ%=<*#=���<`ѻ`j����<�k��   �   �2ܾw���Q��ǅ��$������u׿"��j���ŗ��B%������ֿD��疢�bx���Q�����ܾ䐾t+�9Y���s��Tb�<��/=��Q=ThB=��
=0�L<hWp��5:��Ǟ�v&޽d�4� �+.��2�T�,�������ցԽԎ��l&�0%���<Zv=��N=.�\=@�9=�i�<,0���&���)�� ���   �   ,���{2��Dm�ё����t�տ�������	��6�ҿ	����dP�w_տ�Ѷ�����5�m���2��+��Ϩ���K���ν�S��t�<�L<=��x=Cc�=��j=JY3=���< �\;�����B*�4�y�[䛽+$��8ഽ3���Z󖽌Pl��1�[z����;��<�dB=�?x=�r�=ہ=��F=,Z�<���ɽ��H�7"���   �   ��
�K�B�PV������Tƿ~m��_�|� ���"��v����jL�}翳�ƿ��m�I2D��<�ỻ�{�e��U𽆌$��}V<�nB=R!�=��=l�=xυ=B�V=�Y=��<�/l;�0�X%���뼠������\���h����;���<t%=�je=X��=��=��=/��=ʯM=�<ra�
��ra�!\���   �   ��O�M��"���᫿�п8��������������������>�п׭��~��R[O�ʫ�e�Ǿ�av�:��R�=��p-<��D=�c�=TB�==��=ћ�=[�=ػe=��.=@��<̬�<HZ< �t;@;�y�;@�4<�,�<6�=V_<=�xs=���=n��=H��=��=� �=R�P=h�`<�
/�>~��(mq�ž�   �   ����QQ�bw��A���qӿ�����
���4��ƞ"�.�����&�����3Կ9���Pn��h2S����̾�$|����^F�P�<�E=&��=P��= �=�=�Ŗ=��=X�M=�V=���<��<8~j<P
S<xVy<�Ӭ<���<�$(=sZ=&��=�F�=JJ�=�=�4�=5Z�=|Q=��R<LS7�9P�b�v�
ɾ�   �   ��d�M�("���૿�пC��j����J�f����
�R����_�п���� ��ZZO���U�Ǿl`v�6����=��w-<&E=5d�=�B�=`��=䛟=d�=�e=��.=(��<���<Z<��t;`;�y�;0�4<�,�<8�=X_<=�xs=���=���=h��=��=:�=h�P=`�`< /�Q|���kq�ž�   �   ��
���B�4U�������Rƿ�k��^�X���T!�Fu�`��XK�4{��ƿ���C�p0D�>;�ܹ����e�R�N�$���V<<qB="�=�=Rl�=�υ=h�V=�Y=��<@/l;�0��%��������4��|��������;��<2t%=�je=|��=V��=��=ຎ=�M=��<z\�\��Roa�2Z���   �   {���	2��Am�����տ���F��	�H5�$�	�
��qM��\տ7϶�������m�H�2�(��R̨��K�q�νE��'�<P<=��x=�c�=d�j=�Y3=0��<@�\;����C*�R�y�k䛽?$��KഽB���f󖽜Pl��1��Zz�`��;���<feB=l@x=ss�=�ہ=��F=8c�<����Ƚ>�H�����   �   ;.ܾ(t���Q�xŅ��!�����Nr׿a��u�������E!��B��y�ֿ�@�����v���Q�
��_�ܾ�����+��R��Db���m�<��/=V�Q=�iB=r�
=��L<�Vp��5:��Ǟ��&޽s�D� �<.�"�2�`�,��������ԽҎ��R&�8/%���<0w=@ O=n�\=̷9=�t�<���s �� )�R����   �   �������i2�}�d�T���椿w`��k˿8�տ��ؿ.տ�$ʿhK���٣�t��D�c�>�1���Y���l����D�n��k ��l�<�|=��=�<@5#;�h�] ����� ��MM���t�Hቾ1�������F���d����o�=~G�ʖ�\/ٽ�N��d/̼���;l��<L�%=*.#=���<��л j����U�k��   �   �����Ծy��D<��9h����_z��;���}������i ���Ȩ�)P��_ꇿ�f�"�:��4�jӾ����X�4�C½����];���<w�<���< �3�xH�mw��:���vJ�ZJ��wV���ݿ��lվ��⾅9�k��X&ӾaҼ��ߠ�����&�C�2��7e����	� 
�9�\�<�� =���<pb�;r��m�½p�5��   �   m8Y�aX����(8���Z�6:y�0p��"ُ�p6��)Z������2�v�CcX�K�5��'�G߾��� V�x�����t��ql��tS<C�<���<��:�qL��|*�F�d�D����Ǿُ��f�����#��&��b"����Ҙ	�?��{þl]��k5^�b��%��$�� Vz��}�<���< qW< nr��y��F��   �   ����i�~�����ݾ�L�V�&�`?��R���]���a�|]�IjP�;=�@�$��	��پd����d��=�0���H��@��;�ǣ<`@�<@'V;x��������]�i�������ݾ�N�5�&��?��R���]�¯a��
]�EnP��=���$��	���پ@h��j�d��B���������_�;���<4?�< JV;��~��   �   �F���&���d�����~Ǿ܊�d����\#�_ &�o_"�$����	�m��zvþ$Y��o.^���������� �q����< ��<qW<�xr�:y�I��;Y��𢾨[���f+8���Z��=y�+r��Cۏ��8��f\��ꌇ�V�v�gX���5��*��K߾�����V�Ɍ��^�t��l�xcS<h@�<�Ĕ<���x2��   �   �>��p�����qJ��F��\R��ٿ��gվE�⾷3羞�ι Ӿ&ͼ�+۠�ٺ��<�C����9\���	� �9 k�<� =���<�_�;R��R�½��5�ӝ��I�Ծ�z�#G<�H<h�r��/|��A�������c����"���ʨ�TR��`쇿f�9�:�7�z Ӿ������4��I½"���];���<�x�<`��<��3��   �    �#;�S�W��� �佞� ��GM��t�/݉�А�����������o��vG�g���$ٽ�E��̼@H�;���<�%=�1#=��<��л�j�����k�������gk2�~e�EU��褿0b��[˿U�տ��ؿtտ'ʿ�M���ۣ��u��g�c�ޛ1�.��A\��Ql���F�n��� ��g�<�|= =��<�   �   ,�
=`M<�+p�((:������޽��.� ��x.�q�2���,�<������vԽE����%�@�$�L*�<�=�O=�\=��9=�w�<D ��q!��*)�0����/ܾu�4�Q�Qƅ�#������s׿��b���Ǖ��a#��Z��|�ֿ�B��ӕ���w����Q�����ܾ㐾&+�_W���m���g�<��/=ĳQ=NmB=�   �   ^�j=p_3=T��< R];����l5*���y��ۛ�;���ִ����aꖽ�?l��"��$z�@�;���<RmB=�Fx=�u�=�݁=��F=�e�<t�1�Ƚ҇H� ��X����2��Bm��������տ!������	�&6�
�	����1O�v^տ�ж����@�m�&�2�+���Ψ�9�K���ν\P��� �<�N<=$�x=e�=�   �   tm�=\х=$�V=�_=�<��l;�/�8��\{�`�����⼠i�������;���<�{%=6qe=*��=t��=��=/��=�M=��<~[���Loa�KZ����
���B�jU�����oSƿCl�:_���v���!��u���L��|�<�ƿ���2� 2D�z<�����`�e��U�h�$�(V<�oB=�!�=��=�   �   ���=���=b�=��e=��.=��<ĵ�<@n<@Du;�b;���;��4<L7�<D�=�c<=�|s=dÒ= ��=���=�=/�=@�P=��`<�/�{��	kq��ž��1�M�"���૿	пf����.������H�v������1�пܭ������[O������Ǿ�bv����ڙ=��l-<��D=�c�=�B�=�   �   3s�=���=/�=.�=t�=<�^=b�:=��=��=�"	= �=/&=vE=�k=���=�@�=�a�=���=�3�=b��=�ɯ=匈=��=�~:��О���+�R3��#�٬���U�����ȥ�����6�ڿ�B�����������J���ڿ7U¿�Q���ʈ��LW��?!������1�ͧ�hZz��]=�ց=�I�=���=�   �   �'�=6��=;�=�4�=L�n=b?B=�=���<`��<<��<|��<�=�%=0]O=A}=��=Ĭ�=dɺ=���=A�=t˭=�)�=^s=�] ��9����'�'��Ңܾ)���R��х����u㾿�O׿�}���������Z���v꿲d׿�%�������j���iS��2��z߾������,��ܡ�XE^��X=���=�P�=�\�=�   �   ��=�9�=bH�=� [=�5"=�8�<��j<�G�; V��@����@:���;�\�<��<��1=�Wk=P;�=Bȥ=m+�=X�=`��=�ǆ=��=�����
���0��'�Ͼm:��#G��I~�	2��ܵ��<Ϳ�߿n4뿴+��aX߿�ͿSൿ{e����H� V��,Ҿ(��Z�g���"���=�e�=�<�=�\�=�   �   ���=��s=$�4=��<P�;�+��c׼����<��pE��d7����໼�}Ի�xB<��<zF=~�=n'�=�M�=�Ϝ=(��=��$=�*�:.�_�|��Xq�J���7���	6�PGi��Ď������c�� [ο�ٿ&�ܿ��ؿ��Ϳ�����S��A���Sci�ms6�0���r��C�t�q�
��Hl�������=8s{=���=⁛=�   �    hR=T�
=�d><��[��(!�K���ば��Sӽ���'N���dnͽ�f���t����i	���<T==�b=��=Jf�=��{=��.=Q$<�� ���ݽ�M�홢����+ �RN���}�K��]���"Q��k����,ſ����R����U��\�����|��M������O5����N������)�P�;Z�$=��p=fQ�=�
�=�   �   ��< յ�p?�~�����ҽ����-,�{�D���S�wX�+�Q��A�`'�7���ƽ|�y��pټL�;���<��C=(�j=�th=�d6=|Ӛ<hе����t#$�p텾Q6žJO�׆/��X�5��k��������v��9��I��tM�������~��kW��n.�D��qľ����zv$�9맽$l��q�<�V.=2�^=�Q_=<6=�   �   PD�j%3������_
�1=�?n�1ь��ŝ��e������}I�����t���X�g�iv6�z���䦽	���?�||�<6.=�XK=�@8=��< �����X�Q��!P��
��=�ھ),��"2���S�X;q�v���M��m����⊿�X���Yo���Q��T0�����]ؾ-|��z;N�V,�\'X�Pc��t��<�V2=�JC=`�#=���<�   �   �?��8ƽ��pa��Ȓ�賾�=Ѿ�0�������6M�����| ξ>������Z�r��'��`r/�@k�� ��<�#=.^2=��= �><OѼ����H����k��ɧ���޾.��Vt'��?�(�R���^�TOb�Q�]�+)Q�H�=��f%�X�	��g۾5���,lg����e훽 ɼ��C<Z�=.�.=F�=��<����   �   钿��$#��q�t!���Ѿ ��0v� z ���)���,�K+)�|�ͩ�Ƃ��; ���:�k��F��1��T���U�:���<.�#=�>"= ��< �ӹ�?%�����#�~�q�s��
Ѿ�y��4s��v ���)�R�,�/()���2��@~��I;술�l�k�C�z,���� �:���<ԁ#=�;"=���< �׹`K%��   �   �����k�2ͧ�c�޾���]w'�b�?���R�!�^��Rb���]�U,Q��=�0i%�k�	�	k۾���pg����J񛽴	ɼ�C<6�=B�.=��=�ΰ<�W�f�?��/ƽ��a��Ē�k㳾�8Ѿ+�|���E���G������;1:��6���Z�?��� ��i/��8�����<#=N]2=P�=�><�aѼSȟ��   �   �&P����;�ھ�.��%2���S��>q�I���O��B����䊿_Z���\o�"�Q��V0�H��U`ؾ/~��Y>N�A0�F,X�pw�����<nX2=dNC=.�#=0��<����3�����4Z
��*=��7n�͌�1���a��#���E��쪛������g� q6����ݦ�V��`X?���<(
.=TYK=\?8=t��<ޝ��X�j
��   �   ��9žVQ�N�/���X��6��%�������x���:�����O��	�����~��mW�Zp.�����rľ���Lx$�|��p���o�<�W.=�^=rV_=�6=�(�< ��1�ď��Pwҽ$��0',���D���S�pX�M�Q�OA�MZ'�
2���ƽb�y�Zټ�;h��<��C=D�j=�th=c6=�ʚ<|޵��"�� '$��   �   `���>���- �nTN�V�}��L��� ���R������.ſ�������W��n���N�|�y�M�������l6��j�N�S�Ὠ�)�@
�;V�$=8�p=DS�="�=.oR=D�
=8�><�Q[�0!�����<x���Iӽ1�轐C�����dͽ�]���t����>	�8%�<�C=4"b=R�=�f�=n�{=��.=�?$<�� ���ݽ�M��   �   ��������6�jIi�!Ǝ�����d��k\ο�ٿ��ܿ�ؿ��Ϳ�����T��줎�^di�5t6����js��5�t���
��Il������ =u{=��=䃛=6��=0�s=6�4=@��<Ш�;P�+��H׼��&�<��aE��V7����Ȼ�'Ի��B<@�<�F=��=)�=�N�=М=Ƶ�=D�$=���:��_���^[q��   �   �Ͼ�;�%G�AK~��2��ݵ��=Ϳ��߿y5뿮,���$Y߿�Ϳ�ൿ�e�����H�>V�+-Ҿ0(��Z�7�����؎=�f�=�=�=l^�=��=<�=K�="'[=�<"=�H�<�k<��; ��� d���UB:7�;Dl�<��<� 2=�\k=<=�=�ɥ=^,�=��=b��=<ǆ=T�=ଫ�����2�d����   �   D�ܾ���R�T҅�:��"便aP׿K~�`���Z���ź��jv��d׿�%�������j��wiS�b2�gz߾l���r�,�ܡ��>^�nZ=p��=�Q�=�]�=	)�=w��=~<�=f6�=�n=�CB==���<���<`��<8��<�=��%=B`O=�C}=(��=���=�ɺ=��=F�=6˭=�(�=$q=k �:<��0�'�D���   �   �c��J�U�M���ȥ�>���t�ڿ�B������п���J�ڿ�T¿�Q��Aʈ�%LW�e?!�"����1�i˧�PPz��_=�ׁ=rJ�=@��=�s�=��=|�=r�=��=��^=��:=Ա=��=�"	=�=�.&="E=8k=���=�@�=Va�=f��=i3�=���='ɯ=4��=�=��:�PҞ���+�
4���   �   -�ܾV���R��х����_㾿�O׿]}�c���Y���ƹ��wu�d׿�$������j��}hS��1�>y߾����F�,�kڡ� 6^��[=ꉁ=R�=�]�=)�=���=�<�=l6�=�n=zCB=�=���<���<<��<��<ڦ=��%=<`O=�C}=*��=���=�ɺ=2��=}�=�˭=d)�=�r=�b ��:���'�z���   �   ��ϾA:�P#G�I~��1���۵�'<Ϳ0�߿�3��*��RW߿�ͿOߵ��d��T�H��T��*Ҿ�&���W���� ���=�g�=@>�=�^�=��=%<�=K�=$'[=�<"=�H�<@k<���; ����h���MB:6�;l�<��<� 2=�\k=D=�=�ɥ=�,�=*	�=ꦧ=Ȇ=��=@����
���0���   �   �󻾽��
	6�bFi�VĎ������b���YοYٿطܿq�ؿg�Ϳ6���bR�����5ai��q6����ap��̓t���
��@l������=�w{=釖=`��=x��=t�s=N�4=4��< ��;�+�I׼R��f�<��aE��V7�ʿ�\Ȼ��'Ի��B<P�<�F=��=^)�=�N�=�М=���=��$=�R�:��_���0Wq��   �   �����* ��PN���}�J��2����O������i+ſߣ������:T��ޭ��ԡ|���M��������2��,�N����X�)� C�;�$=J�p=>T�=��=�oR=��
=H�><�Q[�f!�����hx���Iӽ^�轼C�����dͽ�]���t� ���>	�l%�<DD=�"b=��=�g�=X�{=�.=0Z$<2� ���ݽ�M��   �   0셾�4žN�N�/��X��3�����E���u��P7�����K��쮐��~��hW�<l.�5���mľ1����r$�l姽XZ��l�<�\.=l�^=�X_=,6=*�< ꯹1�ۏ��xwҽ?��M',���D���S�pX�e�Q�dA�^Z'�2��ƽ\�y��Yټ���;���<��C=P�j=�wh=�g6=�ٚ<ɵ����!$��   �   
P������ھ�*�� 2�O�S��8q����L������኿�V��*Vo�j�Q��Q0�"���Yؾ�x���6N��$��X����@��<�]2=�QC=N�#=x��<0���3�����FZ
��*=��7n�"͌�H���a��5���*E������������g�q6����ݦ����L?�t��<,.=�\K=^D8=p��<`���H�X�f���   �   ����k��Ƨ���޾,���q'�L�?��R�6�^��Kb�ʱ]��%Q��=��c%���	�+c۾����Jfg�B��c曽D�ȼ0�C<֥=T�.=��=�Ұ<�O���?��/ƽ ��a��Ē��㳾�8Ѿ4+辗���^���G�� ���;=:��=���Z�>��� ��|h/��/��t��<,#=*b2=��=��><CѼ�����   �   �����#�ءq�w��VѾ-u���p��s ���)�"�,��$)�w�B���x���;񄠾ߌk��=�U$��f��@#�:��<6�#=4C"=Ľ�< �ҹ�>%�銿��#���q����$Ѿ�y��Es��v ���)�b�,�<()���;��P~��U;򈠾m�k�C�>,�� ����:T��<T�#=�B"=`��< �й�7%��   �   ԗ?�x)ƽ���ja������߳�4Ѿ+&�3������VB�������;�5��>	���Z��������[/��߁����<�#=fd2=��=�><<LѼ����H��ɥk��ɧ���޾>��jt'�'�?�=�R���^�hOb�a�]�9)Q�S�=��f%�]�	��g۾:���(lg����훽�ȼ��C<P�=D�.= �=ڰ<���   �   ���3������U
�0%=�:1n�jɌ�&����\�������@������������g��j6�����Ԧ���� �>����<.=F`K=F8=��<������X�)��!P��
��V�ھ9,��"2�׶S�r;q�����M��x����⊿�X���Yo���Q��T0�����]ؾ0|��l;N�,�2&X��R��0��<
\2=jRC=�#=�ɮ<�   �   p6�< ����%������nҽ��p!,�A�D���S� iX�J�Q��	A��S'�J,�ٗƽ�y�8=ټ��;���<��C=�j=�zh=0i6=�ؚ<H͵�4��j#$�z텾e6žYO��/��X�&5��y��������v��9��T��}M������(�~��kW��n.�H��
qľ����bv$��ꧽ�h���v�<�Z.=r�^=�Z_=:6=�   �   �tR=8�
=P�><H&[�2!�咃��o��	@ӽ��9�_�彯ZͽaT��V�s�Ă�@
	�h;�< M=�)b=��=�i�=��{= /=`Y$<�� ���ݽ�M�����'���+ �"RN���}�K��k���0Q��z���
-ſ����\����U��b�����|��M������P5����N�5�὚�)��;��$=��p=�T�=4�=�   �   ��=0�s=��4=���<`��;Ј+�00׼����}<�SE��G7�T��D�����ӻx�B< 0�<�"F=>��=�+�=�P�=PҜ=�=��$=�X�:b�_�h��	Xq�U���A���	6�aGi��Ď�ʠ���c��[ο�ٿ2�ܿ��ؿ��Ϳ�����S��E���Yci�rs6�3���r��:�t�S�
��Gl�@���P=�v{=/��=N��=�   �   ��=�=�=M�=,[=�B"=�V�<�.k<֫; ���8����D:P��;�}�<��<�2=ck=�?�=�˥=[.�=�
�=
��=�Ȇ=2�=����q
���0��2�Ͼu:��#G��I~�2��ܵ��<Ϳ�߿y4뿽+��fX߿ ͿWൿ~e����H�V��,Ҿ(���Y�#���H�6�=g�=2>�=>_�=�   �   n)�=��=X=�=~7�=��n=�FB=�=���<`��<x��<t�<��=�%=`dO=xG}=˺�=��=<˺=< �=]�=B̭=*�=t=\ ��9����'�(��עܾ,���R��х����{㾿�O׿�}���������_���v꿴d׿�%�������j���iS��2��z߾�����,��ܡ��C^��Y=B��=�Q�=�]�=�   �   �C�=���=0��=H�=��=*�=�(~=�lg=\�Y=�OV=\�]=D�n=
]�=�W�=��=f��=�A�=[�=�w�=x��=���=&�=�c=�D�<n
	�jԽ��G��`��n��I�v�J���x�����i����(���Ҿ�"¿�;��)��b���̒�L�y�p�K��r���M��L��`ݽ�9�Ho<��T=��=�ٽ=A��=�   �   l��=h��=v�=�I�=���="t�=��d=�wL=(�==��9=*�A=�2T=p�o=��=��=��=6�=�q�=�8�=D��=D#�=̤=��e=@8�<j� �ċͽ�5C�"��v�⾬h��G� �t��'���H��u;��"���&���|����1���P��O���Nu���G��t�H�op��d�G��kֽ`�to�<�W=�ӝ=�;�=O��=�   �   ��=���=��=V	�=��k=�T?=�H= ��<-�<x��<���<�=�$=��M=X�{=vB�=Dܪ=�h�=UU�=b��=�=䊣=0�j=P��<�ϼV���q^5�b����վ[�"�<��`h�.��1e��ܲ���Ȳ�Kݵ�_��������G��d���h��-=����ݿ׾�O��QM9�9½� �X��<�h]=�֜=�A�=���=�   �   ܴ�=P(�=��{=ش@=@=���<���;���@�,�0PG�`��`0� �<�i�<8�=��R=L��=x�=�i�=旹=$�=Π=6ar=��<����t���n��kC���������e,���T���{�q���qC���������F�����������W{���T��p,�.6�F�¾򇄾��"�ʳ�����<��<Z3f=���=/~�=�{�=�   �   ݉=�Z=xe= �<P�����ɼ\X+��a�Л���_��Zx}�d�V�
!�l�� �'� ��<��$=V�k=�ӑ=�P�=���=�ƛ=��y=v�=�.��,�m��f	`�fʧ��a����<��(_�7�}�C���ڑ������S��W���+�|�7^��b;�'���g��a�n��nxu��̻0?=So=N�=tC�=Z9�=�   �   C?=T.�<�̖:<V׼�K_����Ȕ׽�=���J
����������x�ν����6I��k��`��;�e�<؃O=mR�=���=֛�=��~=�*=��<���Ξɽ�l4�ʂ��$z¾m������[>�xMY�nQn�2�{������z��Em�/X��=�I��?(���=��hԉ�W 4��Bʽ�c��9 <d�#=�sv=䥎=�ގ=��|=�   �   D©<P���	-��֢� g�n���?���Y���i���n�e�g�2�U�2�:�����.��*���i���<|>=�x=Ȏ�=�v=JaE=<��<(=y���������W�횾H�ξ>�A����2� eD��O�{9S���N�D=C�� 1�m?��� ��̾���K2U��&��o��x�w�贵<BKA=ay=v�=ҍm=\�0=�   �    �.���K�~�½�.�~�H�*={�)���zm��^��翳�_D���\���/����t��B�T��	~��N�8�*�`T�<f:=`Dn=�z=L�[=��=�m�;�;�()��6�ih��9����ɾk��Rv�5���$$�'��#�����
��]�fkƾ�F��ԝc��U�R����2����;F�=��Z=�fv=,h=H�1=,g�<�   �   ()A���Ƚ�� �Jc�8ɓ�Cᴾ",Ҿ�ez�����D������,Ͼ����$d����\��e�����{3��N�ĕ�<�D=t�m=��l=��@=hS�<Е���A���Ƚ�� �3c��œ�$ݴ��'Ҿ=�ju������N?��a���(Ͼ�~��=a��;�\�2b�D��:s3� ON�М�<��D=4�m=Ҕl=h�@=�F�<�޶��   �   0����
�h��<����ɾ
���x����'$��'���#�x�� �
�{a�nƾrI��١c��X��Į� 9�P��;b�=ގZ=dhv=�h=ډ1=�v�<�t.��K��½�)�_�H�,6{�L���[i���Y������I@���X��N,����t��B�:���w��T�8�@�Ề^�<i:=|En=z=��[=Ɵ= 4�;�E��   �   ���v�W�$���ξj����f�2��gD�֜O�V<S�y�N��?C�9#1�dA�L� �&̾���`5U��(�s����w����<�JA=Xby=�w�=z�m=��0=�ө<���h�,��͢��\��h�I�?��Y���i��n���g���U���:�͙�J&�5疽�� �h�D�<� >=,x= ��=�u=N^E=䪹<H\y�X���   �   �p4�B���@}¾4�������]>�(PY�=Tn��{����u�z�YHm�_X��
=�ޛ��*���?���Չ�f4��Eʽ6g�p2 <��#=�tv=
��=���=��|=FJ?=�@�<�6�:�:׼<_������׽3��&E
����v��������νE����)I��U�� 2�;Ds�<�O=T�=d=웓=l�~=��*=��<���m�ɽ�   �   `��̧��d����"<�	+_���}�����)�������T��p����|��8^�#d;�%(��辠pa����<{u�p�̻�>=�So=8�=�D�=|;�=�߉=�Z=Dn= �<$��X�ɼTI+�,�a�����LW��xh}�~�V�~�tg�� F�,��<��$=��k=�Ց=4R�=A��=�ƛ=�y=�=`Z���m��!��   �   E��������jg,�{�T���{������D���������B�������H���.Y{���T��q,��6�!�¾����X�"���������`��<*4f=���=Z�=�}�=���=�*�=�{=��@=�H=L��<@��; K����,��!G�8�������<�z�<��=ĴR=���=�y�=9k�=���=f�=�͠=n_r=h��<$���#�����   �   �c����վ|	�s�<�rbh����f������sɲ�޵����'���OH�������h�4.=�(��<�׾.P���M9�*9½ ���<�i]=Rל=�B�=��=H�=f��=B��=��=��k=&[?=�O=ȧ�<(<�<`��<X��<��=�$="�M=�{=dD�=�ݪ=j�=V�=���=�=x��=V�j=P��<�ϼ�����`5��   �   :�����}i�q	G��t�?(��cI���;����������ϴ���1��Q��1O���Nu���G��t��G�5p����G�kֽ���q�<
W=nԝ=�<�=��=J��=l��=-w�=UK�=0��=�u�=$�d=|{L=�==4�9=��A= 6T=T�o=��=��=��=�6�=Br�=�8�=N��=#�=�ˤ=<�e=<3�<� �D�ͽQ7C��   �   �a���n�YJ��J�M�x�ȕ������)���Ҿ� "¿�;�d)��3���̒�Ԫy���K��r�M�龟���L�$_ݽN7�('o<6�T=��=Yڽ=���=�C�=ޞ�=p��=�=@��=U�=8)~=�lg=r�Y=�OV=@�]=�n=�\�=\W�=��=6��=�A�=�=�w�=&��=N��=z%�=��c=�@�<	�Խ��G��   �   g������h��G���t��'���H��>;��վ������
���;1��]P���N���Mu���G�t��F�So����G�Giֽf��u�<4W=�ԝ=�<�=8��=b��=r��=4w�=VK�=(��=�u�=�d=b{L=ª==�9=��A=6T=B�o=��=��=��=�6�=Lr�=�8�=r��=L#�= ̤=Z�e=p6�<�� ���ͽ6C��   �   �a����վ#�ǩ<�u`h�����d��P��� Ȳ��ܵ����������F�������h�r,=�����׾�N��K9��5½X�4��<l]=
؜=UC�=F��=n�={��=H��=��=t�k=
[?=�O=`��<�;�<��<���<~�=�$=�M=�{=jD�=�ݪ='j�=JV�=��=��=/��=^�j=|��<�ϼD���V^5��   �   �B��5�����e,���T���{������B������
���4�������r����U{���T�o,��4��¾5�����"�Я��𰚼���<R7f=���=��=�}�=4��=
+�=�{=j�@=�H=䕐<p��;�M����,��"G�H�� ����<dz�<��=��R=č�=z�=ik�=��=�=�Π=Lbr=��<��������ε��   �   �`�Tɧ�`�����<�)'_�f�}�8�������H��SR�������|��4^��`;�>%����ꧾ�a�����ou��p̻�D=�Wo=u�=�E�=�;�=��=�Z=2n=��<�%���ɼ�I+���a�ӓ���W���h}�вV����g�� p���<��$=��k=#֑=�R�=���=�Ǜ=f�y=V�=���<�m���   �   k4�z���]x¾���'��IY>�fKY�On���{�:���z�$Cm���W�D=���{$���:���щ�v�3��<ʽ�Z��U <$�#=yv=b��=��=��|=�J?=�@�<�4�:�;׼p<_����&�׽\3��LE
������������νk����)I��U���2�;�s�<l�O=�T�=9Ô=4��=H�~=��*=h�<����ɽ�   �   �����W�5뚾Ύξ��e����2��bD�L�O��6S���N�}:C�O1� =��� ��
̾���t-U��"�)j����w�(õ<<QA=�fy=�x�=4�m=��0=�ԩ<�����,�$΢�:]�%i�x�?�&�Y���i�7�n�ܻg��U���:���c&�I疽�� �h�T �<�!>=�x=s��=�y=FdE=4��<@+y�����   �   �$��Z��{h�7����ɾɺ�6t����1"$�l'�S~#�b��p�
�!Y�dgƾwC��8�c�jQ�J����'�p/�;0�=�Z=�lv=H!h=b�1=�x�<�s.�$�K�!�½�)���H�b6{�j���yi���Y��ƻ��b@��Y��`,����t��B�F���w��0�8����@`�<�j:=Hn=�z=��[=B�=���;~5��   �   �A�6�Ƚ	� �� c����ٴ��#Ҿ���p������m:�����k$Ͼ}z���]��0�\�6]�B���f3���M����<F�D= �m=��l=�@= V�<𐶻�A���Ƚ�� �bc��œ�Fݴ��'Ҿd龎u������l?��}���(Ͼ�~��La��M�\�<b�C���r3�`CN����<��D=��m=X�l=N�@=�\�<�d���   �   �V.�6�K���½�%�}�H�`0{��𓾣e���U������ <���T���(����t��
B���o����8�0��p�<Lp:=�Kn=�!z=��[=��=�v�;d;�3)��R��h��9��ɸɾ���hv�L���$$�,'��#�����
��]�vkƾ�F���c��U�3���J2�`��;N�=0�Z=�kv=H"h=@�1=\��<�   �    �<����,�8Ǣ��T�*d�Ɵ?�؀Y��i�=�n��g�]�U�a�:�5��n��ޖ����@h�2�<J(>=�$x=葇="{=dE=���<�9y����
����W�8횾h�ξR�X��Κ2�;eD�
�O��9S���N�V=C�!1�z?��� ��̾���S2U�x&��o����w�d��<NA=Ley=0y�=l�m=�0=�   �   �O?=�N�< R�:%׼�._�-��׽g)���?
�F��!������ھνt����I��:��Ќ�;܅�<��O=AW�=Ŕ=f��=V�~=N�*=��<8��Ğɽm4�߂��Bz¾�������([>��MY��Qn�M�{�	����z��Em�>X��=�T��N(��	>��nԉ�S 4��Bʽ�b�H? <��#=twv=l��=Q�=&�|=�   �   �=:Z=*u=(�<�ҡ�Ȓɼ <+���a�ы��EO��lX}��V����L�� Z�̹�<:�$=��k=�ؑ=�T�=y��=�ț=D�y=&�= '����m��~	`�}ʧ��a��� <��(_�R�}�Q���葒�����S��`���:�|�7^��b;�'���o��a�d���wu���̻�@=�Uo=K�=@F�=%=�=�   �   ���=�,�=�{=��@=0P=P��<�E�;����Pn,���F�p������)<��<8�=6�R=���=�|�=m�=���=*�=�Ϡ=.cr=X��<����S���s��vC�� �������e,���T���{�}���}C���������P�����������W{���T��p,�46�M�¾􇄾��"������������<N5f=U��=<��=�~�=�   �   0�=���=ض�=��=4�k=�`?=�U= ��<PJ�<��<��<��=�$=j�M=��{=�F�=�ߪ=�k�=�W�=4��=g�=؋�=f�j=̷�<<�ϼA���u^5�%b����վf�/�<�ah�7��;e��粩��Ȳ�Uݵ�e��������G��i��
�h��-=�����׾�O��NM9��8½��葡<.j]=�ל=LC�=���=�   �   ���=���=�w�=6L�=<��=w�=
 e=�~L=P�==��9=J�A=�9T=��o=u�=�=&�=�7�=Js�=�9�=*��=�#�=�̤=��e=�8�<>� ���ͽ�5C�(��~�⾳h��G��t��'���H��y;��(���+��������1���P��O���Nu���G��t�$H�op��b�G��kֽ �4p�<tW=Pԝ=�<�=:��=�   �   ��=@p�=���=�,�=,O�=���=�Μ=��=)G�=.�=v�=hG�=Fߡ=�=
O�=ܕ�=�N�=���=�E�=V]�=���=���=yk�=>�4=@��;�I�f��yQ�����.۾v=�s�1��AS�@�p�	܃�\4��෍��.���؃���p�܂S��d2������ܾﰟ��5U�h#���Y� ч9��%=E�=Lɶ=4��=hT�=�   �   b��=V��=p�=U�=5Z�=���=?�=�+�=FU�=���=�9�=%֌=�!�=��=�~�=7��=��=xa�=t��=��=�h�=kp�=�"�=0;8=�J�;�?���Z0L�Dv��&�־����.���O�u�l�����݈��U��wԈ�����
�l���O�T /��-�`wؾ0A��FP�R����O�@B�:л)=Z!�=ݏ�=���=
��=�   �   i5�=��=�=���=�E�=���=�j=�aR=�(D=>�@=B:H=�>Z=�&u=|J�=�ԝ=䑰=���=H��=���=���=�I�=�N�=��=��B=��%<b�#�Hֽ��=��鐾��ʾD����%���D���`�iKv�7��%e��X����v�.e`�%�D�P�%��9���˾�H���A���ܽ�91����;�z5=}�=ز�= ��=0��=�   �   잿=X�=BМ=7��=4�Z=�o,=�=�Z�<<��<�;�<��<���<XM=E;=(;k=�"�=2;�=��=F)�=ޝ�=e�=0�=���=��R=���<(`�!.��2�'������7��Ţ���4�4�M���a�X�n���r�^on��{a��QM��3�����񾸠�������)�
�� ��(�l<.tG=N��=Ƹ�=�w�=���=�   �   �p�=Qɏ=үf=�'=���<�<�Cu��4d�p��$����Ú��<� �ι`^<��<�9=��x=W0�=r�=7ͻ=X
�=���=F,�=L�f=���<�iy��!���?��]�������Ҿ.����z�5���G�n=S�OW�j�R��)G���4�6��X���"Ҿ;F���^�o��ݏ�Ɗ�Z�<|]=��=��=�ٸ=�=�   �   �8�=�yH=
�<�6<�W�z�
�6XT�˛��+�����E0�������D�Dy���0�Z<��=��Y=��=��=��=XЮ=�Ǟ=�{=n�=�K:R�<���ս�2�����1��%߾�2��C���)�s�3��07��}3��3)�pI��-��1ݾ蚮������1�Lս��=� �g��=Pu=��=x��=b0�=�C�=�   �   �e7=�{�<��q�����z���.��&8�c+�ӵ�����4U߽����+e�p�ܼ��:L��<(eF=ް�=,�=~�=쳞=N܇=�>>=�Ȍ<p۳��ߑ����2K����� +���Cپ'�����
�S
�o��b����	�[���#�־\Ͱ�������G��2�s뎽L'���H�<�D<=>��=���=��=�#�=8�~=�   �   �<����3�1s������* ��JA��[�n'k��p��Xi��W��<���*�����|���F�����<d#B=ră=�ؗ= V�=�j�=@�f=�U	=@��:NA�|��� �*;P��:���5���¾�ؾ3��/��u���;־>2������u���aTK� �����P���b;��=��g=���=��=*�=�6=�7=�   �   �>����<�)E��B���@���q�i���U_��X󩾿@������S�������Il��?;�ѻ�䯽�Y-� �����<�M=�U�=�X�=�Ɩ=m��=��G=�
�<p���<��=������@���q����[���奄=��N����������Dl��;;�L��tޯ�fQ-�0N����<��M=ZV�=�X�=Ɩ=ӓ�=ԽG=���<�   �   �K�
����9@P��=���8��ۢ¾�ؾI��=��Z��`?־y5��i���Ћ��3XK� ���������a;��=r�g=���=���=��=;=�7=P �<@����3�gk������V% ��DA��[�'!k��p��Ri�G�W�٢<�������ߑ������	��d��<d'B=�Ń=Jٗ=�U�=�i�=��f=ZP	=@��:�   �   7命x��"7K�>���R.��BGپ"����
�{����k����	������־�ϰ�������G�M5���0���B�<C<=��=D=��=�%�=\�~=�l7=L��< Qq��t��z�u�����(3�<&���������L߽D��Xe�t�ܼ��:x��<jF=���= -�=��=���=-ۇ=�:>=ܼ�<�볼�   �   r�ս��2�������d߾r4��E���)���3��27��3��5)�K�/��3ݾƜ�����@�1�bս�=� Hj���=�u=z��=b��=�1�=F�=P;�=ƀH=��<�`<��W�Ԃ
�HIT�䓆� �����\(��B��X�D��a𼘣�H[<v�= �Y=��=*�=��=tЮ=.Ǟ=��{=H�= �:��<��   �   ]B���]�᜞�?�Ҿ������Z�5���G�g?S�>W�;�R�/+G�Q�4�u��_���$ҾxG��o^���Dߏ�\ʊ��W�<�{]=3 �=N�=	۸=��=s�=̏=��f=�'=��<�H<`�t�d��褼D۲�ܫ����<� wɹX7^<`&�<��9=�x=l2�=��=8λ=�
�=Θ�=�+�=��f=l��<��y��%���   �   ��'������9��*��:��4���M�X�a��n�g�r��pn�/}a��RM��3�_�� �񾟡��F���ʿ)�>��j���l<4tG=���=d��=�x�=ל�=���=i�=�Ҝ=4��=�Z=Tw,=�=0l�<0	�<�M�<��<0��<�T=�K;=�@k=%�="=�=��=Z*�=���=��= �=���=4�R=䓌<k��1���   �   ��=�N됾��ʾ>����%���D�Ϙ`��Lv�����e������zv��e`���D�Ƣ%��9�i�˾I���A��ܽ�91���;f{5=f}�=[��=���=��=�6�=2!�=0�=���=H�=��=j=�gR=�.D=�@=�?H=DZ=�+u=�L�=�֝=m��=���=1��=T��=D��=�I�=�N�=�=��B=X�%<�#�HKֽ�   �   �1L�Ew��Y�־=��ٿ.�l�O�@�l�~����݈� V���Ԉ��K�l���O�e /��-�IwؾA���P����ԉO�@d�:ļ)=�!�=S��=(��=���=��=(��=d�=!V�=i[�=���=��=,-�=�V�=���=;�=a׌=#�=��=v�=���=v��=�a�=���=��=�h�=p�=�!�=J98=�4�;��?�r���   �   xQ�����x/۾�=���1�%BS���p�"܃�i4��෍��.��g؃�I�p���S�Wd2�=��M�ܾ\����4U��!����Y� ˈ9��%=�E�=�ɶ=���=�T�=��=|p�=���=�,�=TO�=���=�Μ=��=2G�=+�=f�=RG�=*ߡ=��=�N�=���=�N�=���=RE�=]�=���=F��=�j�=Ə4=Е�;��I�����   �   �0L�wv��O�־����.���O�>�l�󡁿V݈��U��"Ԉ�`���B�l��O��/�J-�.vؾ1@���P�ʦ��O�@��:�)=I"�=���=V��=���=$��=(��=`�=V�=`[�=���=��= -�=�V�=���=;�=X׌=#�=��=o�=���=z��=�a�=���=��=�h�=Qp�=^"�=�:8= C�;4�?�����   �   t�=��鐾��ʾ��;�%�7�D��`��Jv�����d������Wv��c`���D�9�%��8�O�˾iG��nA�i�ܽj41����;~5=I~�=�=��=T��=�6�=<!�=3�=�=H�=���=�j=dgR=�.D=Ұ@=�?H=�CZ=T+u=�L�=�֝=i��=���=B��=t��=z��=)J�=*O�=��=�B=�%<B�#��Gֽ�   �   �'�u����6�����*�/4�$�M�l�a��n�E�r��mn�6za��OM�q�3�:����񾸞�����`�)�1������l<�wG=���=6��=dy�=&��=���=v�=�Ҝ=)��=��Z=w,=�=�k�<��<�L�<@�<���<�T=hK;=�@k=%�="=�= ��=�*�=ʞ�=�=��=��=��R=���<�]�0-���   �   �>���]�����$�ҾB��Ğ��5��G��;S�yW���R��'G��4������= ҾD��^���8ُ�����\d�<@�]=�!�=G�=�۸=�=Cs�=!̏=��f=�'=�< G<`�t��d�x餼0ܲ�����(�<� �ɹ6^<�%�<��9=�x=z2�=*�=�λ=f�=���=-�=ȧf=���<�`y�0 ���   �   �ս��2�p���~��	߾O1�
B���)���3��.7��{3��1)�{G��+�[.ݾ'���d���o�1��
սض=� �`�~�=�u=��=v��=�2�=gF�=z;�=̀H=H�<`_<@�W�^�
��IT�/���L������(�������D�0b�����[<b�=�Y=��=��=H�=vѮ=�Ȟ=�{=��= 	:J�<��   �   �ܑ�Ո��/K������(���@پ����ֱ
�`�c��J����	�x�����־6ʰ����j�G�l/��厽����V�<.J<=��=�Û=��=I&�=
�~=�l7=,��<�Uq�u���z����+��\3�m&�߰�B���M߽z���e��ܼ��:���<fjF=첅=�-�=��=��=�݇=:A>=�ό<Lҳ��   �   �:�=�������7P��8���2��
�¾:ؾt��E�����7־�.��F}������dOK�����x����� �b;.�=Z�g=��=b��=��=X<=N7=� �<���3��k��; ���% �EA��[�d!k��p��Ri�v�W���<�������������������<(B=Fƃ=Jڗ=jW�=�k�=6�f=�Y	=�5�:�   �   ����<�t8��k�o�@��q�B|���X��K쩾�9����������v���>l�Z6;�ڳ�ׯ�`E-�@�� �<�M=�X�=�Z�=RȖ=\��=��G=p�<`���<��=������@�,�q�6���[���奄;=��n���+�������Dl��;;�b���ޯ�nQ-�@L����< �M=CW�=Z�=*Ȗ=ꖅ=v�G=�<�   �   ��<���:�3��e������! ��?A�%[�Vk��p��Li�_�W�K�<�������=����������T�<4.B=xȃ=�ۗ=#X�=�k�=��f=�V	= ��:tA����� �b;P��:���5��H�¾�ؾ^��V�龙���;־X2����������}TK������&���b;��=��g=��=��=��=�>=*7=�   �   �q7=H��< �p��j��tz�S
����罬.�n!����~���C߽�����e��ܼ i�:0��<@qF=���=|/�=��=���=m݇=�?>=ʌ<8۳��ߑ����2K�����E+���CپV�����
�j
����u����	�z���<�־pͰ�ì����G�	3�l뎽�&��`J�<F<=X�=wÛ=&�=2'�=P�~=�   �   r=�=2�H=)�<ȁ<�W�Rw
�2<T�����V	���	��t ��������D�G�t� 7[<�=8�Y=��=��=��=hҮ=ɞ=ܮ{=v�= i:L�<���ս�2�չ��S��N߾�2��C���)���3��07��}3��3)��I��-��1ݾ��������$�1�Fս~�=� �f�*�= u=���=���=43�=�G�=�   �   �t�=@Ώ=
�f=b'= �<8l<`�s���c�(Ѥ�,ò�������<� �ù�_^<�8�<��9=̮x=H5�=Y �==л=��=|��=\-�=��f=$��<�hy��!���?�D�]�ƚ����ҾB�������5���G��=S�fW�}�R��)G���4�A��b���"ҾHF���^�s�pݏ�Ŋ��[�<t}]=� �=+�=ܸ=�=�   �   ҡ�=��=�Ԝ=���=��Z=�},=D!=$|�<�<�^�<L%�<(��<�\=S;=�Gk= (�=�?�=0��=$,�=��=�=b�=v��=��R=���<�_�,.��I�'�����7������!4�I�M���a�n�n���r�qon��{a��QM���3�������à�������)�
�������l<.uG=��=�=�y�=ĝ�=�   �   N7�=,"�=t�=���=�I�="��=�j=�lR=04D=��@=xEH=�IZ=�0u=O�=�؝=\��=���=���=���=`��=�J�=�O�=:�=��B=8�%<8�#�Hֽ��=�ꐾ�ʾP����%���D���`�yKv�@��-e��_����v�7e`�-�D�V�%��9���˾�H���A���ܽL91����;�{5=�}�=���=��=���=�   �   R��=���=��=�V�=9\�=���=���=j.�=X�=P��=<�=�،=p$�=�=���=���=b��=�b�=d��=X�=�i�=�p�=�"�=x;8=L�;�?���`0L�Mv��2�־����.���O�~�l�"����݈��U��{Ԉ����l���O�W /��-�dwؾ3A��HP�L���O� I�:�)=�!�=<��=*��=���=�   �   ���=���=�B�=rC�=>�=�r�=���=�Ѯ=���=ƻ�=bJ�=�=C��=�4�=B��=�6�=�[�=&��=`y�=|D�=pz�=� �=�=��=j'=P'���nd�"����E��ʎ��Ѿ��y�e;�F�%�J6��A�A�D�*�@�m?6���%��_�1񾸿������H�X��@r����Vp=�~=�k�=���=`��=$��=�   �   ���=ZV�=���=���=��=���=Hk�=���=�7�=�A�="�=T�= -�=�d�=ܹ�=��=��=*p�=:��=�j�=6l�=���=�~�=�	�=��=`�T��;Z��z�UA����	�����l��]�"��3�{�=�52A� �=��2���"�����e��ֻ�5ތ�{�C����n2g� bԻ��=P~�=Q�=X^�=h��=���=�   �   ���=ʣ�=8~�=���=���=L��=ր�=VL�=�ֈ=���=��=Nؑ=懜=�ʩ=�{�=UN�=���=���=p��=B��=N�=K��=�Ĵ=fӊ=�>!=���:��<�v׽$t3���6����޾������/�)���3��7��3��o)������p�޾���c����5��۽�|G�@���Y=΄=;��=���=Ե�=��=�   �   f�=Ĥ�=��=�	�=T:�=�B�=�\a=��I=0z;=��7=<z?=lcQ=�Dl=��=|��=ͬ=;=h�=�&�=B"�=B�= ��=�z�=᪐=�e6=� <���_ල���[j��ߞ�<�ɾp��KM�����$��7'���#�˅�5�����ɾ8Ϟ�D�j�7�f$������;�;�,=�u�=� �=���=��=��=�   �   ���=��=4�=�}=�AK=N�=|a�<PQ�<�x~<�}j<�<�d�<�V�<8
*=�E[=��=�S�=$��=*��=��=�|�=��=��=�ޗ=`bQ=`��<�s���������CG�Z��p����Ծ����v��v?�������,�������Ӿh���^���F�W��>��\������<tJ=,��=�g�=���=
��=���=�   �   LѤ=ɚ�=�[=`;= �< ��;X����ɼ��׼����T.�� ݜ���<��<μ*=��k=Pj�=|ѫ=�f�=xy�=N~�=���= ��=��o=��=@N�N=�/gǽ�h��j`�Ժ��g����ξ�4徢u�n$��<�����A;����
I���
^�����eŽ��;��']����<"Vk=̍�=f>�=N�=�1�=JE�=�   �   J�=�[D=k�<���;��q�Z��`�Y��/����������ԗ����L�K������)��:<�="�S=���=9�=F��=@��=��=���=�ʇ=��4=X�p<�����兽l 뽯~,�S�d�����ʷ��;���+nľ�EȾp�þ�7�������ŋ��@a��1)���彅����p��0fz<��4=�߆=�(�=��=���=�a�=�=�=�   �   E>=��< ���1��l�ng��rݽ>Z�p��Z�p�M2���ս�����Z�h�ͼ@/; ��<��J=\��=6�=�E�=��=�Z�=��=��f=p=@�;8�	��T�����+�'�T�({��ڌ�ru�� ���m���<q���cw���O��O#�!���y���5����;B�
=��i=Ar�=2��=��=��=f@�=���=�   �   @�<@Rc����ʒ���ܽ���_�0���H���W���\��fV���E��,�%@���ӽs������ g�$F�<lKR=̍=�q�=t��=��=xޤ=0�=�`J=�<��b���KĒ��ܽ1����0�o�H���W���\��aV��E���,�s<�z~ӽD󉽤�� �`��O�<�NR=0͍= r�=j��= �=@ݤ=P�=`[J=�   �   �^;��	��Z����n�'��T�q-{��݌�Xx�����4����s��$hw���O��R#����Z~��PC���~�;�~
=<�i=�q�=!��=~��=��=
B�=���=2K>=/�< ���<�l��_��8wݽ�U�����U��k�.*����ս6����Z�{ͼ`�;���<�J=穉=*�=�E�=�==Z�=3�=d�f=�	=�   �   �����ꅽ�&뽎�,���d�F�������<���>qľ�HȾZ�þ]:������ǋ�Da��4)�C�������z���Wz<t�4=�ކ=h(�= �=���=3c�=�?�=���=�bD=@{�<��;��q�Ƞ���Y��(���������{͗�����K�o��X�(�p?:<��=,�S=���=��=��=~��=6��=���=ɇ=.�4=�xp<�   �   BV=�jlǽ�k��n`�#�����s�ξ�7徳x�s'����~�D;�����J��t^�õ��hŽ<�;� \]����<�Tk=���=�>�=��=�2�=�F�=vӤ=z��=x[=6C=,2�< Գ;0�������|ɼ��׼����h������ <\��<@�*=��k=`l�=ӫ=�g�=
z�=j~�=[��=��=��o=�=�iN��   �   �������GG�>��������ԾQ�������@�W�<��^��������Ӿ౮�E_����F����)���������<�J=��=h�=��=���=լ�=H��=�=�6�=:�}=�HK=@�=�r�<hc�< �~<�j<.�<�u�<Lf�<(*=�K[=r�=�U�=���=]��=��=}�=��=�=�ݗ=^_Q=���<����   �   �㶽>�i^j�eើ2�ɾ���vN�����$��8'���#�Ć���"
�?�ɾО���j�	8��%������3�;��,=�u�=� �=d��=x�=��=��=b��=��=�=�<�=�E�=ca=��I=�;=l8=Ѐ?=�iQ=4Jl=7�=���=�ά=�ξ=��=�'�=�"�=NB�=���=:z�=���=�b6=��<L���   �   {׽v3�������L�޾���{���)���3��7�ʌ3��p)��������޾���������5���۽x}G� ���2Y=D΄=���=��=h��=D�=f��=��=��=���=v��=6��=悗=~N�=�؈='��=@��=Lڑ=���=�̩=}�=�O�=���=Z��=���=���=T�=��=qĴ=�Ҋ=�<!=��:$�<��   �   }뽺A�|Ë��
���������"��3���=��2A�|�=�S�2��"�����e�׻�&ތ�N�C�=��1g�P[ԻL�=�~�=��=�^�=���=���=h��=�V�=���=���=��=���=Tl�=���=9�=�B�=0�=J�=�-�=Ke�=���=�=��=lp�=f��=�j�= l�=h��=D~�=*	�=��= �T� ?Z��   �   ����E�4ˎ�Ҿ�ez�;�x�%�>J6��A�A�D��@�I?6�V�%�r_���:���|��P�H����r�����q=�~=Fl�=ؓ�=���=X��=Ε�=���=�B�=�C�= >�=�r�=���=�Ѯ=���=ƻ�=WJ�=��=2��=�4�=��=�6�=j[�=���=8y�=HD�=6z�=� �=��=���=�%=�5��6qd��   �   X{뽘A����	�����X��7�"��3�(�=��1A���=���2�P�"����d�
ֻ�]݌��C�]���.g�KԻȉ=-�=�=�^�=���=��=p��=�V�=���=���=��=뇸=Hl�=���=9�=�B�= �=<�=�-�=@e�=���=�=��=tp�=v��=k�=<l�=���=�~�=�	�=��=��T��<Z��   �   -׽�s3������0�޾�������)���3��7�-�3�o)�-�������޾"~��9���4�5�
�۽xG� /���[=Bτ=5��=���=���=n�=���=��=��={��=h��=%��=Ђ�=aN�=�؈=��=&��=4ڑ=���=u̩=}�=�O�=���=d��=��=���=��=|��=Ŵ=yӊ=
?!= ��:D�<��   �   \߶�9��Zj��ޞ�E�ɾ3��L�����$�o6'���#��������2�ɾ�͞�w�j��4�� ��N��0_�;��,=(w�=��=��=��=&��=��=j��=��= �=�<�=�E�=�ba=:�I=��;=8=x�?=TiQ=�Il=�=���=�ά=�ξ=��=�'�= #�=�B�=���={�=8��=xf6=�	 <z���   �   ������^BG�Y ��%�����Ծ����Z��:>�������φ�������Ӿ=���<\��ЧF����; ������ܕ�<TJ=���=0i�=���=p��=��=f��=�=�6�=�}=^HK=ҏ=�q�<xb�<�~< �j<,-�<�t�<�e�<�*=ZK[=]�=�U�=���=���=�=�}�=W�=�=0ߗ=�cQ=ؾ�<8o���   �   J=�vdǽ�f�2h`�U������q�ξ2��r�!��L���
�?;����F���^�p��l`ŽJ�;�`�\�<��<@Zk=���=�?�=��=23�=4G�=�Ӥ=z��=D[=�B=H1�<�ϳ;�������~ɼ��׼����|������� <���<$�*=��k=jl�=*ӫ="h�=�z�=/�=���=˗�=\�o=��=`�M��   �   �|���ⅽ��&|,�(�d�ʫ����������jkľ�BȾ�þ�4������ Ë�$<a��-)�w��\󁽄`��(�z<��4=��=Q*�=P�=b �=�c�="@�=���=nbD=�z�<��;@�q�|��`�Y��(��􁚽{����͗�A��z�K��o����(��>:<`�=4�S=���=��=���=L��=j��=���=�ˇ=6�4=�p<�   �   �#;�	��P������'�U T��#{�D،��r��^}�������n��`^w�3�O�nK#����s��H"����;z�
=��i=Tt�= ��=���=✰=�B�=0��=LK>=�.�<@��0���l�U`���wݽV�*���U��k��*����ս����Z��{ͼ`�;���<$�J=&��=��=�F�= ��= \�=��=V�f=
=�   �   d&�<�eb�r������6�ܽ�����0��H���W���\��\V�$�E�I�,�>8�wӽ�쉽ܾ� �W�(^�<�TR=�ύ=t�=4��=��=/ߤ=��=�`J=�<��b�����Ē�u�ܽr��ݵ0���H���W�ȍ\��aV�B�E��,��<��~ӽw���� �`�P�<LOR=�͍=�r�=���=��=�ߤ=��=4dJ=�   �   �O>=:�<����	�ޮl��Y��FpݽR����FQ�fg��!����ս������Y��dͼ =;\��<J�J=���=P�=�G�=���=\�=.�=6�f=�=��;��	�8U��&��j�'�VT�j({��ڌ��u��D�������\q���cw��O��O#�[��z��6��p��;��
=@�i=�r�=,��=���=6��=bC�=���=�   �   ���=fgD=t��<�B�;@�q�t����Y�"���z���~��NƗ�����ĞK��V���(��d:<��=��S=H��=��=� �=5��=ڥ�=x��=ˇ= �4=��p<H����兽� ��~,���d�٭������g���Unľ�EȾ��þ�7�������ŋ��@a��1)��彛����p��gz<b�4=��=b)�=��=� �=od�=hA�=�   �   դ=���=�![=rI=�@�<��;���ߕ��fɼ��׼������� 8��)<ī�<��*=tl=$o�=Rի=�i�=�{�=��=���=���=d�o=��=`N�lN=�{gǽ�h��j`��������Źξ�4��u�$��a�����A;����I���
^�ĳ��eŽ��;�`%]����< Wk=���=�?�=��=�3�=<H�=�   �   ���=��=�8�=&�}=xNK=ږ=���<�s�<P�~<X�j<�?�<膶<�v�<�*=jR[=h�=LX�=�ô=2��=O�=v~�=��=d�=(ߗ= cQ=�< t��µ��D��DG�x������D�Ծ��������?� ����<������0�Ӿy���*^���F�f��K�� ������< J=���=�h�=���=ȳ�=��=�   �   ��=���=B�=��=?�=@H�=�ha=��I=<�;=�
8=H�?=�oQ=0Pl=��=,��="Ѭ=xо=3!�=�(�=�#�=fC�=��=V{�=K��=*f6=� <����ල��[j��ߞ�Z�ɾ���\M�����$��7'���#�څ�@����.�ɾFϞ�^�j�&7�r$������=�;��,=)v�=<�=���=�=���=�   �   ���=���=|��=���=؍�=͡�=���=nP�=�ڈ=C��=\��=dܑ=���=^Ω=�~�=Q�=���=~��=���=^��= �=���=ZŴ=�ӊ=L?!=@��:��<��׽>t3���K��ϱ޾�����=�)���3��7��3�p)������z�޾���k���&�5� �۽�|G�����fY=_΄=���=T��=���=��=�   �   ���=HW�=��=H��=n�=���=1m�=���=:�=D�=:�=X�=�.�=@f�=f��=��=��=q�=���=�k�=�l�=���=�~�=�	�=��=��T��;Z��z�bA����	�����s��e�"� 3���=�<2A�&�=��2��"�����e�׻�8ތ���C����n2g�PaԻ��=s~�=��=�^�=���=��=�   �   Z��=���=p�=�,�=���=L�=���=��=��=�6�=�L�=_��=b��=h,�=�^�=(w�=�y�=Dh�= 2�=X��=j �=�e�==��=܉�=��s=���<�x延�T��ֽ&�(�[k�UƗ��฾�P־Ѝ�5q��P� �G^��vv��K־
���%���Ml��Q*�J�ڽ��^��o�@#�< Th=��=[��=�v�=`�=�g�=�   �   ���=@�=���=�#�=���=���=��=B�=t~�=�պ=c�=��=z�=	�=H��=���=�'�=��=2'�=
$�=�G�=8�=
�=�r�= Qw=� =`����J�wн\]$�v�e�:����:��2Ҿ����5���Z������Ҿ�J���픾��f���%��	Խ2HT�`��R�<(
l=T��=�C�=�?�=M�=���=�   �   l��=�=�|�= �=��=F��=ա�=���=�p�=���=�
�=:��=��=�s�=���=���=�)�=Ы�=x��=$��=��=�!�=(��=��=���=
= P��6�-��弽�%�|�V����잪��9ƾ2�۾ �龝��<��Z�۾�ž�t������QCW��6�����Z5��A��s=�v=�Ҧ=[�= ��=v��=<��=�   �   $�=�^�=pu�=���=�3�=�r�=���=,��=J�=.�=�=��=DK�=�?�=���=��=�\�=��=Hx�=�8�=���=�D�=��=�2�=��=�&=�1<N  �ޞ�� ���>�'�z��������ВǾ�`Ծ��ؾsԾWǾ����������y���>��T�Մ��&,����;�=��=D��=���=<�=>[�=$<�=�   �   d�=���=.Z�=�ԡ=�Ύ=��y=��Z=hC=� 5=$}1=�8=�IJ=��d=q�=���=��=8}�=���=�l�="N�=��=�:�=���=CN�=v�=�E=Tՙ<����ڿp�dٽ� �,GV��ℾ�����������Bļ�8����鬾;ך��	��s�T�2�� ؽ8�p����4y�<��?=���=J��=3��=܉�=���=��=�   �   T��=t��=���=j�x=�|F=^4=���<�О<гr<��^<���<@z�<t��<Xv$=PU=/σ=�K�=�c�=Y��=���=b��=��=$ �=M׺=�=h=���< �ܹ~��3&��������,���Y�$���&��1����,���~���K�����iW�6�*�~����_��@-� ��`H�<p�e=�	�='�=���=b��=���=�f�=�   �   �g�=&q�=�\=�=�D�<p��;��»���(³���������X�b�`�J�h�+<��<]+=>rk=�=�A�=�ֿ=���=��=@��=u3�=���=b��=b,4=@��<�}k�L��᳽P���{'���H�m�b��,s��px��r�Y�`��,F�Ǝ$��b��r����^C���Q����<�C6=L��=ݧ=Ȑ�=.�=�B�=w��=M޺=�   �   ��=l�O=��=�I:<p%����4�9��n�/����l���S��X�e�&�-� RͼF����v<	=�;\=M]�=ze�=�=`y�=��= ��=7��=�E�=�i=��=H?<̻��"GW�%D��޲�F-��e&���3�@�7��2��=$��G��彚z����J�|l��8�0<|=en=���=jP�=XA�=�m�=��=�ƺ=��=�   �   PT=t��<��;�����g8�,z��UH��Iܽ�#񽱋��0��ݬ׽<��Dn����)�(��x<=�]=P�=<�=��=<��=(R�=J�=	�=f��=j!T=`
�<P[�;�n���\8�t���A��.ܽ,�h���*��M�׽6��i����)���� <�"=X]=��=�<�=櫿=:��=�Q�=+I�=�ު=v��=�   �   �=0#<�̫�lQW�!J������0��i&�ų3�@�7�ތ2�|A$��J�8�g��x�J�Hy��0�0<�{=dbn=��=�O�=HA�=]n�=X�=Ⱥ=:�=@�=�O=��= k:<0��l�鼄�9���n�͛��\f���M����e���-�h?ͼp����v<�= @\=�^�=�f�=��=�y�=���=���=8��=ED�=�i=�   �   �y�< �k�L�糽v��'���H���b�1s��tx��r��`��/F���$��g��r���"eC���Q�d�<$A6=e��=�ܧ=���=�.�=yC�=���=�ߺ=�i�=�s�=�\=�=U�<0�;L»�������������誼�b��]J�X�+<���<�b+=wk=��=8C�=�׿=*��=8��=��=�2�=���=ī�=�'4=�   �    �߹����*�������,�0�Y����#(��L���/������`M���!�glW���*�E���|b���1� >��C�<�e=(	�=b'�=/��=��=���=�g�=�=|��=�=<�x=x�F=�;=��<��<��r<��^<���<H��<��<�|$=U=�у=�M�=ge�=���=���=֚�=��=��=�ֺ=��=�h= ��<�   �   𭊼��p��ٽ|� �2JV�^䄾�����������/Ƽ�	����묾�ؚ���}�T�Գ��ؽ�p�����<u�<F�?=6��=9��=b��=H��=���=��=��=���=.\�=*ס=@ю=h�y= �Z=C=�5=��1=��8=PJ=L�d=�=A��=�	�=�~�=5��=�m�=�N�=��=�:�=P��=�M�=`�=�E=�̙<�   �   \% �.ួ��5?�՝z�"��"���z�Ǿ/bԾ1�ؾ�Ծ�Ǿ���������y��>��U�,���.� ��;�=u�=D��=���=��=�[�=�<�=�=�_�=�v�=q��=�5�=�t�=���=���=�L�=��=��=��=dM�=�A�=,��=Q��=�]�=��=�x�=9�=���=�D�=���=
2�=��=2�&=8"<�   �   n�-��輽F'�`�V�"������;ƾu ܾ<��ɧ�J��C�۾��žcu�������CW�$7����� �5� I�~s=�v=�Ҧ=P[�=h��=���=ƪ�=��=��=�}�=,�=e��=���=\��=���=.r�=A��=/�=���=�=u�=���=���=�*�=\��=���=`��=��=�!�=���=S�=��=�= `���   �   �J�fн�^$���e�����I;���2Ҿ�龛���Ѵ��ڙ��o��*Ҿ�J���픾��f���%��	Խ�GT� ��(S�<�
l=���=/D�=@�=jM�=V��=X��=�@�=:��=�$�=R��=���=���=�=G�=�ֺ=*�=���=(�=��=���=��=(�= ��=P'�=$�=�G�=�=�	�=or�=�Ow=� =`+���   �   ��T� �ֽƑ(�k��Ɨ�6Ḿ�P־��Qq��P� �,^��Dv�K־����%��LMl��P*�3�ڽ��^��i��%�<Uh=l��=���=(w�=��=�g�=|��=��=��=-�=���=_�=���=��=��=�6�=�L�=S��=Q��=R,�=�^�=w�=�y�=&h�=2�=0��=@ �=�e�=���=|��=��s=���<0���   �   ��J��н�]$���e�5���g:���1Ҿ��s�����������Q��!Ҿ�I���씾��f�l�%�	ԽET� ��V�<�l=���=xD�=P@�=�M�=f��=\��=�@�=6��=|$�=J��=���=���=��=8�=�ֺ="�=���=�=��=���=��=(�="��=Z'�="$�=�G�=.�=�	�=�r�=�Pw=$ =����   �   ��-��弽\%���V�����j���9ƾb�۾
�龈����$�۾��ž�s��z���tAW�5�X�{5���`v=0�v=�Ӧ=�[�=���=��=��=$��=��=�}�=%�=X��=���=H��=r��=r�=$��=�=���=�=�t�=���=���=�*�=`��=���=x��=J��=�!�=?��=��=��="= p���   �   � ��ܞ�
 ���>�יz����������Ǿ#_Ծ�ؾ�Ծ�Ǿ����9�����y���>��R�����'���;�=��=T��=��=�=\�==�=2�=�_�=�v�=]��=�5�=�t�=ғ�=v��=aL�=��=g�=��=@M�=�A�=��=:��=�]�=��=y�=D9�=��=>E�=^��=�2�=��=ڧ&=�5<�   �   8�����p�Oٽ�� �iEV��ᄾp������q���y¼�^���
謾t՚�"����T������׽*�p�����H��<$�?=���=���=A��=܊�=���=<��=��=���=\�=
ס=ю=�y=��Z=�C=>5=��1=P�8=�OJ=��d=��=$��=�	�=�~�=:��=�m�=�N�=B�=:;�=��=�N�=��=JE=�ؙ<�   �    q۹����#��_�����,�!�Y�����h$��[����*���|���I����'fW��*�'���[���%� ����Q�<F�e=�=�(�=&��=���=��=�g�=
��=t��=��=�x=�F=P;=���<���<��r<X�^<���<H��<@��<�|$=�U=�у=�M�=de�=���=���=:��=���=� �=�׺=��=�h=X��<�   �   ԋ�<�lk���K�#޳�$���x'���H� �b�)s��lx��r�j�`��(F�Y�$��\��,����UC���Q���<�H6=4��=�ާ="��=�/�=D�=��=�ߺ=�i�=�s�=��\=�=T�<0�;�Q»D ��������� ꪼ��b��fJ�`�+<��<�b+=�vk=��=SC�=ؿ=���=ҁ�=���=44�=���=^��=�.4=�   �   �= Q<|���@W��?�����P*�_b&�)�3�~�7�6�2�.:$��C���t���yJ��[��(�0<2�=�in=ޏ�=�Q�=�B�=Ro�=��=xȺ=g�=F�=�O=X�=�h:<�����V�9���n�=����f��N��~�e�B�-��@ͼ0	��x�v<^=�?\=_�=�f�=$�=Dz�=���=���=��=�F�=��i=�   �   �$T=��< ��;Xa���T8�>o��$<��ܽ��}��@��׽�/��'c��J�)��v��?<P)=�#]=���=�>�=d��=���=S�=�J�=_�=���=T!T=�	�<�V�;8p���]8�zt��B���ܽ��������׽t6��Ui��@�)�����<�"=p]=��=;=�=n��=��=�R�=�J�= �=���=�   �   ��=4�O=��=��:<���4��¶9���n����``���G���e���-��*ͼ@����w<p=�E\=Ta�=�h�=h�={�=D��=���=���=F�=:�i=h�=�=< ����GW��D��]�뽊-��e&��3���7�B�2� >$��G����z����J�m����0<�=Ten=B��=�P�=B�='o�=6�="ɺ=��=�   �   *k�=lu�=��\=d!=�a�<`K�;p	»x쁼���`����Ԫ��Xb� �I���+<P��<�i+=�|k=i�=IE�=�ٿ=���=���=L��=(4�=&��=���=d,4=Ą�<�k��L�⳽����{'�"�H���b�(-s��px�%r���`��,F��$�c������_C���Q����<�C6=���=�ݧ=r��=�/�=ID�=v��=��=�   �   8��=��=��=Ԯx=҈F=�A=���<��<��r<��^<0��<`��<p��<��$=lU=jԃ=BP�=sg�=I��=*��=��=,��=!�=�׺=`�=Rh=���< ݹ���&��	����,���Y�H���9&��W���-���~���K�����iW�Z�*������_��|-� ���H�<Ԡe=�	�=(�=���=���=r��=�h�=�   �   ��=���=�]�=�ء=cӎ=H�y=l�Z=C=�5=f�1=*�8=`VJ=@�d=�
�=¼�=��=���=۹�=�n�=�O�=��=�;�=O��=�N�=��=8E=0ՙ<d���d�p��ٽ� �fGV��ℾଛ�����@���eļ�X��� ꬾSך��	����T�N��< ؽv�p�@���\y�<��?=ӻ�=�=��=Ԋ�=4��=҆�=�   �   ��=�`�=x�=Φ�=p7�=�v�=���=̜�=�N�=�=��=I�=�O�=�C�=��=��=c_�=��=�y�=:�=���=�E�=���=�2�=��=4�&=h1<�  �<ޞ�� � ?�Z�z���������Ǿ�`Ծ��ؾ�ԾnǾ����������y���>��T��>,���;�=��=���=��=��=D\�=v=�=�   �   ���=j�=x~�=�=p��=� �=���=���=�s�=Ζ�=��=D��=��=ev�=���=���=�+�=4��=���=��=���=4"�=z��=�=��== �n�-�漽�%���V� �������9ƾK�۾�龲��P��l�۾ �ž�t������`CW��6����f5��A��s=T�v=
Ӧ=o[�=���=$��=��=�   �   ���=�@�=���=�$�=���=%��={��=��= ��=�׺=��=���=��=R�=j��=���=�(�=���=�'�=t$�=�G�=x�=>
�=s�=Qw=� =����J��нm]$���e�D����:��$2Ҿ����A���c������Ҿ�J���픾��f���%� 
Խ>HT�@��R�<P
l=r��=D�=@�=lM�=p��=�   �   ��=���=�8�=��=�Q�=���=���=Ĩ�=�8�= ��=��=�,�=���=|/�=>r�=���=���=���=�] >���=���=V��=� �=e��=��=ʆi=@��< �⺖}�����j���'-��xY��_��Eۏ�Nř�D)�����ď��S��,�Y���-����P��B�$��k����<
N`=O;�="��=��=��=z��=��=�   �   n��=��=̰�=`�="��=��=P��=�$�=���=��=���=���=`Y�=
W�=��=ƥ�=�m�=>��=8/�= q�=�F�=&��=�C�=+�=?�=`-m=`= P���c��읽�����(�k�T��D{�ތ�����x񙾯���辌��{�6�T�K)�Bq��|���C� M纨��<�Rd=~��=~P�=PE�=Vv�=���=���=�   �   ��=��=(�=(�=�`�=��=��=F��=�v�=���=��=�4�=���=���=t��= ��= ��=jv�=�x�=	�=��=��=ʣ�=���=Z��=��w=�A=���;���'=���⽈��vF��Vk��.���s�������Q�������j��&F�m��bF�	������� fh;U	=�p=�v�=�~�=D��=$��=���=,��=�   �   ���=pR�=NS�=���=r��=8r�=B{�=í=�֩=:��=�J�=p��=�z�=�`�="q�=N��=HO�=d-�=Tq�=/�=�b�=��=�"�=:��=P�=Ha�=�>(=�WR<�2���e�E�½x�	�.K0��fR�0m�F?~�����j�}�h|l��Q���/�%	��½�f�p㦼C<q##=K�=a��=D��=���=~u�=Vy�=���=�   �   �z�=@��=�J�=Uh�=�*�=H��=�4�==�j�=3�=.��=���=�s�=F�=���=��=pf�=~��=���=4��=p��=R|�=H��=�N�=��=�P�=,IG=(n�< �ڻ�"�\M���R�����2���J�u�Y���^�:4Y���I�|S1�����
�؝��� �p?ٻ|��<�`D=J8�=on�=�'�=���=�d�=]�=��=�   �   Ž�=U��=���=���=d#�=�~{=��]=�+G=t�9=@;6=6==4�M=��f=�3�=�.�=��=}�=���=��=X��=���=��=��=�,�=�=��=�.k=dO=ط
<�ԩ��T�oC��A��X��-#�JT0��4��/�;�!�]��	��Ϧ��#N��䠼�<Tb=�j=�=�d�=���=p��=�[�=Έ�=��=�   �   ��=蘭=�}�=�z=��O=q�"=�2�<D��<��<��<���<�e�<��=r@.=�\="�=���=N3�=���=(�=vy�=��=��=���=2��=^r�=�҈=<�A=��< ���߼F�]�x?[н�������^������`f̽y��D�T��μ ��:���<�]E=,��=��=a��=���=���=t2�=F��=���=�   �   ë=���=��l=0=���<X�j<�V;`�ۻhI��@c�؏:�຤� T�;���<�K�<JI<=,x=$ݗ=7�=4
�=H�=4��=��=�F�=%��=���=OF�=lv=�.(=ڢ< x'��jͼܕ=��|������X����G��4�J��n��b3�HB�� ���T��<0�/=�{=�7�=W�=�=���=�Q�=b��=l��=^e�=�   �   �J�=�i=n�!=��<�0;0�o�P�6(��E���M�<�A��E!�̏߼ �C��]�;���<u,=Z0r=��=��=���=�z�=�+�=���=�K�=���=$	�=pL�=Fi=�!=< �<��0;�{o�t=�h(��E���M�~vA��<!�0߼XzC����;��<�y,=�3r=R	�=��=u��=�z�=�+�=X��=�J�=���=��=�   �   pv=�)(=�͢<��'�4{ͼ*�=���������Ӱ��dM��v󱽷O������i3��O�� D̸$��<��/=J�{=�6�=��=��=���=�Q�=���=V��=�f�=�ī=��=��l=�0=���<��j<`�;��ۻ��H�c�Hm:��y�����;$��<W�<6N<=Dx=�ޗ=P8�=�=��=t��=ؕ�=PF�=l��=���=�D�=�   �   �A=(�<�_��߼��]�L󢽅`н1�����a�V�����j̽}���T�`�μ@�:`��<[E=,��=l��=��=��=$��=�2�=��=���=���=���=��=�=��O=�#=�@�< �<XΛ<<(�<�Ϣ<�s�<h�=@F.=�\=P	�=d��=�4�=ķ�=��=�y�=��=��=N��=n�=6q�=Lш=�   �   <K=0�
<�᩼JT��G���E罎[��0#�W0���4���/���!����ӫ�IҦ��(N� ���<�_=�j=o�=pd�=���=���=2\�=t��=��=���=ط�=t��=次=�%�=�{=��]=�1G=ĸ9=�A6=X== �M=�f=L6�=�0�=��= !�=��=��=��=��=��=���=,�=N�=��=v+k=�   �   Pf�< �ڻ�"��P���V���z�2� �J��Y�`�^��6Y���I�qU1�Z��k������ ��UٻT��<H_D=�7�=+n�=p'�=���=8e�=�]�=���=�{�=r��=L�=j�=�,�=k��=:7�=Z��=Nm�=�5�=���=���=�u�=2�=^��=��=�g�=t��=N��=���=���=Z|�=��=zN�=,�=dO�=.FG=�   �   �IR<�;��jf�e�½D�	�*M0��hR�?2m�zA~����g�}�0~l�v�Q���/�6	�8½��f�`禼�C<l"#=�J�=A��=C��=���=�u�=�y�=t��=T��=ZS�=fT�=6��=���=�s�=�|�=�ĭ=�ة=�=�L�=$��=\|�=:b�=\r�=`��=(P�=.�=�q�=p/�= c�=��=�"�=���=��=A`�=<(=�   �   0��;8���S?��o������wF��Xk�f/��_t��f����R��������j��'F���UG㽻���t���@\h;�T	=|p=�v�=�~�=t��=Z��=��=���=���=���=��=�=�a�=��=6��=t��=x�=��=7��=6�=���=���=H��=й�=���=�v�=�x�=<	�=��=���=���=v��=���=�w=�?=�   �    @ķ,f�a�
����(�o�T��E{��ތ�"��������*����{�p�T�&K)�Wq��s���C� D�L��<Sd=���=�P�=~E�=�v�=��=,��=���=j��=.��=��=���=���=��=z%�=���=��=}��=���=�Y�=xW�=�=��=�m�=d��=T/�=&q�=�F�=��=�C�=�*�=�>�=,m=�=�   �   @���S���H��A(-�-yY��_��eۏ�]ř�E)��ܴ���ď��S��ØY�J�-��������$�@�j����<�N`=�;�=h��=��=��=���=��=��=���=�8�=��=�Q�=���=���=ƨ�=�8�= ��=��=�,�=���=v/�=,r�=���=���=��=y] >p��=���=*��=� �=#��=f�=�i=(��<�   �    ���d�흽�����(�F�T�bD{��݌�`����?���l����{�8�T�J)��o�����,A�����<4Td=��=�P�=�E�=�v�=*��=>��=���=h��=,��=��=���=���=س�=j%�=���=|�=u��=x��=�Y�=pW�=��=��=�m�=j��=Z/�=4q�= G�=$��=�C�=�*�=�>�=-m=�=�   �   0��;�����<��?����quF�Vk�.���r��ꗐ�Q��<���G�j�5%F����C�찎�h��� �h;bW	=�p=Lw�=&�=���=���=B��=���=���=���=��=��=�a�=��=!��=X��=�w�= ��= ��=�5�=���=���=4��=̹�=���=�v�=�x�=P	�=�=8��=��=���=j��=��w=
B=�   �   �[R<0��"�e��½��	�J0�JeR�r.m�t=~�����Y�}�Nzl��Q�Ã/�j	�{½�f��ڦ�`C<?&#=7L�=V��=��=v��= v�= z�=���=\��=XS�=\T�=&��=���=�s�=�|�=�ĭ=Xة=� �=jL�= ��=:|�=b�=Cr�=R��=P�=.�=�q�=�/�=8c�=0�=&#�=}��=��=�a�=�?(=�   �   `q�<ЋڻJ�"�~K��qP�^��L�2���J�C�Y�w�^��1Y�I�I�'Q1������f���:� ��ٻh��<�cD=�9�=zo�=d(�=P��=�e�=�]�=��=�{�=l��=�K�=�i�=d,�=>��=7�=(��=m�=^5�=h��=ȍ�=�u�=
�=@��=i��=�g�=p��=Z��=���=���=�|�=���=NO�=W�=Q�=vJG=�   �   nQ=��
<Ω�bT��@���=��V��+#��Q0�b�4�D�/���!���u���ʦ�bN�8ؠ�p�<�f=D�j=j�=�e�=���=P��=�\�=�=��=��=ͷ�=_��=���=�%�=j�{=�]=X1G=:�9= A6=�
==��M=��f=6�=�0�=��=� �=��=��="��=4��=���=b��=-�=��=T��=20k=�   �   ��A=��<���\�޼f�]��ꢽ7Wн��N��@\��
����ea̽~t�� �T���μ Z�:Ч�<�aE=ⵉ=|��=���=��=���=j3�=`��=��=���=���=��=P=0�O=i#=�?�<�	�<͛<�&�<x΢<�r�<��=�E.=�\=/	�=J��=�4�=Ϸ�=�=8z�=H�=`�=P��=Ҁ�= s�=�ӈ=�   �   �v=�1(=�<�)'��^ͼ��=��x��-��������B��鱽�E�����<Y3��2�� $��(ʹ<�/=(�{=�9�=��=@�=���=�R�=h��=���=�f�=�ī=�=<�l=|0=\��<�j<��;��ۻ��H�  c� p:� ��@��;��<PV�<�M<=x=�ޗ=Y8�=:�=��=���=���=LG�=ҽ�=���=MG�=�   �   �M�=bi=��!=�)�<��0;�ao�t.�(��
E�R�M�$mA�V3!��m߼8ZC��ʵ;d�<�~,=x8r=@�=V�=���=|�=�,�=X��=L�=��=<	�=dL�=�i=��!=�<`u0;o� ?�H(�jE�n�M�NwA�@=!���߼�|C�Ќ�;� �<<y,=�3r=Z	�=��=���=]{�=D,�=J��=DL�=���=$
�=�   �   �ū=���=@�l=`0=���<��j<�F;0Jۻ�H�P�b�L:��8��p͚;l�<d�<�S<=$!x=���=
:�=��=��=���=Җ�=LG�=���=��=]F�=Lv=d.(=٢< �'�lͼ��=�}�����Ы��eH���7K������b3�HC�� ������<
�/=�{=�7�=��=v�=���=�R�=���=��=�g�=�   �   ���=��=���=��=>�O=4	#=�L�<��<�ۛ<H6�<�ݢ<���<� =RL.=�\=��=���=�6�=F��=0�={�=��=��=F��=���=�r�=�҈=�A=��< ��P߼�]���[н!����_���b��f̽dy��̶T��μ@��: ��<�]E=;��=@��=���=���=���=�3�=���=���=�   �   ��=���=���=���=�'�=H�{=��]=>7G=h�9=\G6=0==��M=|�f=�8�=.3�=��=�"�=q��=�=��=��=���=���=-�=[�=��=�.k=O= �
<(֩��T��C���A�+Y�.#��T0�/�4��/�o�!����U��VϦ�$N�8堼0�<>b=��j=+�=	e�=(��=��=�\�=��=��=�   �   �|�=b��= M�=bk�=.�=+��=,9�=y��=�o�=�7�=���=:��=x�=2�=0�=��=i�=���=X��=���=���=}�=Ћ�=LO�=$�=�P�= IG=�m�<��ڻ��"��M��,S���<�2�ǌJ���Y��^�l4Y��I��S1�Ъ��
����b� �0Aٻ8��<�`D=h8�=�n�=�'�=��=�e�=^�=P��=�   �   ���=
T�=8U�=5��=��=u�=i~�=uƭ=(ک=��=EN�=Җ�=�}�=�c�=�s�=���=4Q�= /�=�r�=0�=�c�=��=T#�=���=z�=Xa�=�>(=�VR<�3����e���½��	�ZK0��fR�<0m�t?~������}��|l��Q�Ʌ/�<	��½h�f��㦼�C<n##= K�=���=���=(��=v�=z�=���=�   �   ���=��=n�=��=|b�=��=.��=���=&y�=:��=[��=.7�=Ǵ�=���=.��=���=f��=|w�=fy�=�	�=Z�=x��=��=��=t��=��w=�A=@��;����W=�� �⽧��=vF�Wk��.���s�������Q�������j��&F�|��~F�$���Ԥ�� eh;U	=�p=�v�=�~�=���=���=J��=إ�=�   �   ܑ�=���=l��="�=���= ��=X��=�%�=&��=�=��=��=fZ�=�W�=z�=���=@n�=�=�/�=xq�=4G�=V��=D�=*+�=?�=h-m=N= ���c��읽����(�~�T��D{�ތ������񙾷�����{�>�T�K)�Xq������C��N纨��<�Rd=���=�P�=tE�=�v�=��=@��=�   �   K >���=x,�=lb�=��=���=P��=�B�=(n�=J-�=|��=�a�=ܒ�=r��=w�=��=� >5�>��>I>�2 >2�=���=t��=j��=�X�=�n=ds=�X <���d�E�qY����ڽ�$��P��/(�D�,�p(�Z(�x���ڽ`ߠ�X�G�D�����<��=L�g= ��=L��=f��=(��=��=���=L��=�   �   �f�=H�=N�=�)�=ҋ�=L�=�j�=��=��=��=h�=��= ~�=���=��=���=�9�=�>�>f�>F��=0��=���=FG�=�\�=V��=Ļq=�X=�e9<����zI<�_њ��xԽB���o��$�nh(���#��:��d�V^Խ�(���>� ��� q(<�=fzk=#�=,��=�B�=���=vl�=DC�=���=�   �   ���=���=���=z�=���=���=��=��=���=�^�= ��=�E�=<@�=�w�=&_�=~R�=ܤ�=��=R >B� >V�=���=��=�~�=x��=Lm�=�t|=��$=�B�<��4�J� ��������&_�F&�77��J������Ԣ�Y������ĳ!���<�8�u<O =@w=V�=�Y�=���=��=,��=���=�^�=�   �   ��=���=�(�=jB�=\�=�+�=y�=�=���=3�=���=���=~��=E�=���=�9�=b8�=`��=x��=�x�=r	�=��=h)�=Vb�=J��=�q�=���=4C;=�< �D��p�b�����b�ѽ�������M	�H�����tн�|��,�`�,��`���·<�j8=��=H��=9��=\%�=��=l��=t��=���=�   �   �3�=b��=��=�u�=+��=��=vz�=�(�=�t�=x��=&��=���=d�=B8�=��=ڈ�=���=��=l��=�=���=�^�=�7�=��=���=�@�=.��=�X=X�=P2<�]x�:	!�\P~�kا��~ǽ�x۽��O�ڽ�ƽ���6^z��z���m�t<#=p�W=ɡ�=8��=�`�=D#�=�)�=6��=$��=��=�   �   R3�=d��=ѓ�=� �=���=Mݣ=z�=���=D)�=���=>~�=*��=��=�E�=w�=B�=��=���=R��=��=*(�=Xx�=��=g�=/;�=`J�=R��=��z=3.=H´<�_:쪼`�'���o����������L�������j�h|"�pN�� ��:,�<x}0=�u{=�Y�=y�=���=�x�=��=$��=H��=���=�   �   ���=4��=俶="x�=
.�=Q�= �l=ZX=��K=]H=�kN=_]=($t=��=��=ӌ�=���=��=��=bv�=�8�=.��=<q�=��=
9�=6��=lO�=b��=��\=O
=t)�<�>�������P	�¿8��VV�ا_���S��N4��\������s:���<y�=J%a=;�=�=C�=���=l��=t��=
Y�=�@�=���=�   �   T��=�?�=���=��=�df=�>=��=��=�_�<v�<���<
�=�	#=��F=zp=�č=�T�=�{�=�,�=d��=h	�=r�=6E�=2R�=��=r��=�N�=D�=~F�=t�N=��=�ǚ<��;��	� 8���Kż�HԼ���X���޻�v�;��<F�=��U=@�=H��=��=(��=`X�=���=V3�=�]�=��=H��=�   �   �u�=�{�=c�=�R=��=���<���<�B�; �?;@v�: +l;�<��<d��<��%=[= �=�+�=���=�A�=���=x��=�j�=F�=��=��=F��=8w�=�}�=d�=~R=�=|��<���<Py�;`n@;�S�:��l;X�<x'�<���<�%=�[=�!�=8-�=���=UB�=���=���=�j�=�=���=�=D��=�   �   �B�=�D�=4�N=��=��< �;(�	��F��dZżPWԼ(��xe��`A޻�K�;��<F�=@�U=�>�=H��=��=���=X�=���=�3�=^�=���=2��=���=nA�=T��=�=�if=�>=��=�=`l�<���<��<��=�#=��F=�p=Pƍ=V�=�|�=�-�=��=�	�=��=.E�=�Q�=D�=���=�M�=�   �   ꓏=�\=�=,�<@��������W	�4�8�v^V�r�_�"�S��U4��b�����H:��<>}=�"a==�=L
�=��=p��=X��=���=`Y�=0A�=���=���=���=y��=�y�=&0�=��=�l=�X=�K=tbH=�pN=
d]=�(t=��=��=f��=��=��=t�=�v�=&9�=X��=*q�=:�=~8�=`��=LN�=�   �   ��z=|/.=���<�:������'��o�2�������������������j���"�0W���k�:<�< {0=�s{=�X�=�x�=f��=�x�=&��=l��=Ȯ�=4��=64�=~��=(��=w"�=���=@ߣ=��=���=�+�=���=t��=@��=��=�G�=�x�=ZC�=0��=���=��=���=|(�=rx�=��=�f�=�:�=�I�=5��=�   �   >�X=��=�!<�px��!�VV~��ۧ��ǽ5|۽:⽀�ڽ�ƽ�����bz��~�h�m�j<,!=�W=<��=���=�`�=:#�=�)�=r��=���=���=R4�=F��=��=�v�=���=b��=|�=v*�=lv�=E��=京=/��=��=�9�=:��=��=���=���=���=d�=���=�^�=�7�=���=��=�?�=!��=�   �   �@;= ��<�J����2�b�G���)�ѽ������
O	�SI����vн}~�� �`���鼠��ܿ�<�i8=���=
��=��=V%�= ��=���=���=4��=���=0��=�)�=ZC�=n�=�,�=Lz�=l��=��=��=8��=���=���=F�=p��=l:�=9�=���=؇�=�x�=�	�=��=J)�=b�=ě�=+q�=��=�   �   ��$=�=�<`�4��� ��������La�\'�F8��K�n�b��(���Z��a����!���<�@�u<�N =�w=V�=�Y�=���=��=T��=ʝ�=�^�=\��=���=2��=�z�=p��=t��=j�=��=|��=�_�=��=�F�= A�=Fx�=�_�=S�=N��=X��="R >R� >b�=x��=��=^~�=	��=�l�=ls|=�   �   qW=�^9<�����K<��Қ��yԽ��Kp�W$��h(�-�#�A;��d��^Խ�(���>����Pq(<�=�zk=(#�=J��=�B�=���=�l�=vC�=���=�f�=NH�=`N�=*�=4��=��=>k�=���= �=Z��=��=P�=d~�=��=X��=���=�9�=�>�>n�>L��=��=r��=G�=P\�=ᢟ=��q=�   �   �r=�T <�!��z�E�Z��|�ڽ%��P�0(�E�,�[(�0(�@��ڽ�ޠ�4�G�$�@�<e�=�g=J��=���=���=X��=6��=���=d��=K >���=�,�=tb�=��=���=T��=�B�=.n�=L-�=|��=�a�=Ғ�=l��=w�=��=� >,�>��>�H>�2 >�=���=B��=*��=jX�=n=�   �   �X=�d9< ����I<�Qњ�_xԽ��`o�]$��g(�0�#�N:�d�]Խ�'��|>�����w(<<=�{k=�#�=���= C�=��=�l�=�C�=���=�f�=HH�=\N�=*�=,��=��=2k�=v��=�=L��=��=>�=X~�=���=V��=���=�9�=�>�>t�>N��=0��=���=:G�=�\�=:��=��q=�   �   �$=�C�<p�4�^� �u���$���^�%�k6��I������Ϡ�W��������!���<���u<Q =�w=�V�=HZ�=&��=@�=���=��=_�=f��=���=*��=�z�=b��=d��=T�=h�=d��=�_�=���=�F�=�@�=6x�=�_�=�R�=D��=X��=(R >\� >~�=���=��=�~�=���=[m�=u|=�   �   �C;= �< �����&�b�D�����ѽ�������bL	��F����QrнEz����`�$�����xȷ<4m8==��=��=�%�=j��=��=���=J��=���=*��=�)�=DC�=L�=�,�=,z�=H��=Ƞ�=f�=��=���=���=�E�=P��=X:�= 9�=���=ڇ�=y�=�	�=��=�)�=�b�=u��=r�=@��=�   �    �X=��=�9<�Sx�(!��L~�2֧��{ǽ�u۽��2�ڽ� ƽ����Xz��u��tm�ȃ<l&= �W=碐=*��=�a�=�#�=h*�=���=���=���=^4�=@��=���=�v�=u��=<��=�{�=E*�=:v�=��=���=��=��=�9�=��=؉�=���=���=��=z�=���=
_�=8�=R��=��=A�=���=�   �   �z=�4.=�ƴ< :�䪼��'��o�����������飽#���&�j�\v"�tC���{�:��<��0=�x{=�Z�=z�=}��=vy�=���=̂�=��=P��=>4�=n��=
��=Z"�=���=ߣ=Z�=���=I+�=���=:��=
��=֭�=|G�=�x�=EC�=��=���=��=���=�(�=�x�=Z	�=tg�=�;�=�J�=拞=�   �   :��=��\=�=0�<�����x��hK	�Թ8�fPV��_���S��G4�V��뉼��:��<��=�(a=��=<�=K�=���=.��=(��=�Y�=lA�=���=���=n��=V��=�y�=�/�=d�=~�l=�X=t�K=�aH=tpN=�c]=P(t=ޑ�=��=H��=崻=��=x�=w�=V9�=���=�q�=��=~9�=���=P�=�   �   E�=�G�=.�N=��=�Ϛ<:�;H�	�L,���>żD;Լ\���J����ݻ0��;�(�<�=��U=�A�=���=��=,��=8Y�=V��=4�=n^�=��=J��=���=QA�=&��=��=@if=D>=ݢ=e�=�j�<0��<��<4�=>#=�F=Lp=)ƍ=�U�=�|�=�-�=(��=

�=��=�E�=�R�=F�=��=vO�=�   �   #x�=�~�=���=�R=�=���<�ʀ<��;��@; �:@�l;8�<D3�<���<�%=T#[=�#�=�.�=ꆷ=vC�=���=���=Dk�=��=d��=��=Y��=0w�=z}�=2�=R=l�=��< ��<s�;�a@;@<�: �l;��<D&�<���<��%=�[=x!�=(-�=���=fB�=(��=��= k�=��=���=`�=��=�   �   d��=}B�=���=��=`mf=>=5�=*�= w�<���<4�<T�=#=��F=(p=Lȍ=�W�=2~�=�.�=��=�
�=l�=�E�=�R�=�=���=�N�=D�=VF�=��N=�=Lƚ< �;��	��9��,MżJԼX��hY��p޻`r�; �<��=P�U= @�=D��=��=R��=�X�=��= 4�=�^�=D��=��=�   �   ���=���=�¶=c{�=�1�=x�=�l=X=��K=PgH=�uN=�h]=Z-t=4��=�!�= ��=���=J��=��=�w�=�9�=��=�q�=��=J9�=W��=mO�=J��=d�\=�	=\(�<�S��`����Q	���8��WV���_���S�|O4�J]�����T:��<*�=%a=2�=�=j�=���=���=��=�Y�=�A�=J��=�   �   �4�=R��="��=�#�=��=��=L�=���=~-�=���=���=E��=�=nI�=Hz�=�D�=r��=���=���=R��=0)�=y�=|	�=lg�=c;�=tJ�=L��=\�z=�2.=<��< ::���'���o�󇓽q�d�����٥��>�j��|"�DO�����:��<H}0=�u{=�Y�=4y�=���=y�=���=܂�=@��=̱�=�   �   �4�=���=���=�w�=���=���=�}�=�+�=�w�=ࢪ=���=�=p��=;�=���=��=���=���=���=	�=\��=T_�=<8�=H��=̍�=�@�=!��=��X=��=P0<�_x��	!�
Q~��ا��~ǽ)y۽:⽤�ڽƽe����^z�\{�(�m��r<�"=F�W=ȡ�=R��=a�=�#�=:*�=���=���=��=�   �   ��=���=,*�=D�=<�=�-�=X{�=���=��=��=n��=���=���=(G�=d��=F;�=�9�=���=f��=xy�=
�=��=�)�=�b�=c��=�q�=���= C;=x�<��0����b�������ѽW���͔��M	�'H����'uн�|����`����@��P·<�j8=��=T��=Z��=�%�=6��=ޝ�=��=���=�   �   ���=J��=���=.{�=���=��=�=B�=D��=�`�=���=tG�=�A�=�x�=b`�=�S�=̥�=Ԥ�=WR >�� >��=���=��=�~�=���=Nm�=�t|=w�$=LB�<�4��� �N���1���\_�g&�R7��J������ ���Y�������!�x�<���u<�N =8w=*V�=�Y�=���=�=z��=���=2_�=�   �   
g�=nH�=�N�=@*�=r��= �=�k�=���=~�=���=@�=��=�~�=h��=���=6��= :�=�>�>��>|��=V��=���=XG�=�\�=V��=��q=�X=he9<����I<�vњ��xԽP���o��$�~h(���#��:��d�j^Խ�(���>�L����p(<�=dzk=#�=8��=�B�=���=�l�=~C�=��=�   �   D>��>  >�}�=�^�=�`�=L��=�|�=��=���=N�==�=�{�=F��=Z��=�6 >I->(�>�O>��>5c>2��=l��=0��=�,�=�=H�=HV�=�7=p�<@�;��o����L�2��ɐ�j��j���0��V�K������q��ѥ; e�<�Y4=؂|=tl�=[�=c�=�U�=� �=@��=�v >��>�   �   ��>i� >^��=���=���=�O�=��=��=��=�w�=��=���=�C�=�z�=*(�=,��=�|>L>9�>8�>�$>4G�=���=,��=���=pٽ=X2�=n
�=��;=�}�<p��;8cR�ȥ �\�B�Fdv�����WR���u��4B��R ���S���; a�<��8=n�=n՟=[#�=���=޲�=f4�=��=�= >��>�   �   �k >�x�=,��=���=���=��=D��=���=H�=(�=�7�=(��=L��=�R�=x��=|��=���=�O>�q>��>!k>��=���=���=|t�=���=���=V�= nH=��<�v:<`4��@�м��'��;Y��wx��z��6�w��-X�B�&�8�μP���@
9<��<d.F=m�=���=W"�=غ�=<��=j�=�=n&�=�� >�   �   �=�=8��=Ɩ�=��=}�=b��=į�=2�=`��=D��=���=R��=�_�=J��=�J�=b��=���=T��= >d� >�7 >zH�=���=\�=�&�=`��=���=��=M\=�P=� �<�
:0僼���ND+��CH���Q�(_G�x�)������� �}:��<T6=�6[=bލ=�y�=��=��=>g�=���=�=���=^��=�   �   ���=��=��=^�=�G�=��=<��=�9�=n��=n �=d��=o0�=���=�j�=�)�=�3�=���=�=���=���=��=���=V}�=.��=���=bX�=³={%�=J%v=��4=D_�<0�8<� ��L���@�߼�-
�N��x����ۼ<熼��S� �C<D��<x:6=�zv=�̘=�=��=r��=�~�=���=��=~��=��=�   �   Ц�=x�=�=vD�=�a�=2�=Ll�=&��=&8�=�i�=�E�=P��=qH�=���=�M�=Bc�=�5�=d�=�M�=�]�=X��=t2�=�-�=ti�=��=���=�м=��=�'�=\�Y=^
=x;�<�%< Ӻ@.�\ ���ܓ������"��:�p6<�Y�<� =T�\=2�=�~�=x��=!�=���=���=�)�=���=���=2�=�   �   L��=(��=S��=�u�=��=e��=dğ=x�=Y�=��=�/�=���=,��=��=�=~�=���=�e�=�6�=���=@��=DQ�=̘�=�,�=���=���=��=
�=��=��=T�L=�=��<lw<�t�; 2"; �~:�o>;��<П�<�L�<�`=�Q=d�=r3�=�1�=�6�=���=�i�=3�=!�=~\�=�'�=N��=�   �   ک�=$t�=���=_�=6��=�W�=mB�=�Pt=�Qi=Nf=lxk=mx=��=�ƒ=�W�=�ڰ=�R�=_��=0��=l�=T��=X��=`��=��=|�=L��=��=�T�=�T�=+l�=�B}=�bP=h�&=	x=,��<̳�<��<8��<�Y�<ڇ= �,=��V=E��=�3�=��=P.�=���=pa�=l?�=�a�=���=�m�=���=���=�   �   ]�=�׻=���=^��=���=��d=�,G=d�0=w'#=?6=z>%=�4=ШL=�5k=	5�=<�=��=�ƾ=���=<Q�=(��=X��="9�=���=���= `�=�d�=^�=�ػ=c��=��=���=��d= 1G=�0=:,#= ;=C%=v�4=ЬL=�9k=�6�=��=��=�Ǿ=a��=�Q�=���=���=(9�=v��=���=|_�=�c�=�   �   �S�=�S�=�j�=\?}=�^P=�&=]s=h��<Щ�<��<|��<�P�<��=<�,=^�V=ޭ�=�2�=,��=�-�=$��=a�=6?�=�a�=���=n�=��=,��=���=4u�=ߡ�=��=ꗝ=xY�=mD�=�Tt=,Vi=`Rf=�|k=qx=� �=RȒ=RY�=?ܰ=�S�=<��=��=��=���=���=^��=���=$�=���=V��=�   �   	�=Ń�=M�=؉L=�=��<Yw< M�; �!;�n}: ">;p�<t��<E�<�]=�|Q=<�=�2�=�0�=J6�=@��=�i�=�2�=0!�=�\�=:(�=���=��=��=r��=w�=�=��=(Ɵ=�y�=@�=���=�1�=z��=Ѫ�=J�=q�=,�=���=�f�=�7�=��=���=bQ�=Ș�=^,�=F��=���=U��=�   �   ��=O&�=h�Y=�=�3�<��%<��Ӻ�$.�(*��d擼�&��0�"��;��6<�S�<{� =8�\=X�=�}�=���=� �=^��=x��=�)�=���=��=��=v��=B�= �=�E�=�b�=~3�=�m�=���=�9�=�k�=G�=Ϊ�=�I�==��=�N�=>d�=�6�=�=N�=P^�=���=�2�=�-�=Bi�=x��=*��=м=�   �   �$�=#v=��4=�X�<��8<@ ��ē���2
�������H�ۼ$ T���C<��<�86=|yv=̘=��=��=L��=�~�=���=J��=���=@�=��=���=ִ�=D�=�H�=<��=p��=0;�=���=��=���=�1�=З�=�k�=�*�=f4�=z��=N��=��=��=��=���=F}�=���=B��=�W�=\��=�   �   ��= K\=5N=d�< B:�냼D��� H+��GH���Q��bG���)���������Q}:ȳ�<�4=�5[= ލ=[y�=���=���=4g�=���=0�= ��=���=@>�=���=\��=«�=�}�=6��=���=$�=P��=<��=���=8��=�`�=��=.K�= ��=0��=���=* >�� >�7 >�H�=���=,�=f&�=���=,��=�   �   ��=^lH=��<�m:< H��t�мF�'��>Y�bzx��{����w��/X��&��μ����x9<t��<�-F=�l�=���=A"�=ֺ�=B��="j�="�=�&�=͝ >�k >$y�=���=l��=8��=R�=���=`��=�H�=��=H8�=���=ڕ�=tS�=���=���=���=�O>�q>��>(k>��=p��=v��=,t�=V��=t��=�   �   �	�=��;={�<`��;�iR�x� ��B��ev�����4���R���u�R5B�S ���S� ��;a�<��8=v�=x՟=j#�=���=��=�4�=0��=�= >��>��>�� >���=���=��= P�=f��=��=f��=�w�=X��=���=�C�={�=\(�=`��=�|>[>C�>A�>�$>,G�=���=��=@��=$ٽ=�1�=�   �    V�=v�7=�<��;Ȓo�$���L�J2��ɐ�j��Q������̣K�����q� ץ;�f�< Z4=d�|=�l�=��=��=�U�=� �=R��=�v >��>D>Î>  >�}�=�^�=�`�=L��=�|�=��=���=P�==�=�{�=D��=P��=�6 >C->"�>�O>��>,c> ��=Z��=��=�,�=��=�=�   �   Z
�=��;=x}�<��;�bR��� ���B��cv�v�������Q��|�u�3B�
Q �h�S����;�c�<��8=��=�՟=�#�=���=��=�4�=D��=�= >��>��>�� >���=���=���=P�=\��=��=Z��=�w�=L��=���=�C�={�=X(�=V��=�|>X>D�>@�>�$>>G�=���=$��=t��=bٽ=H2�=�   �   n�=DnH=L�<(y:<�-����м�'�:Y��ux��y����w�T+X���&�H�μ�����9<���<�/F=�m�=X��=�"�=<��=���=Vj�=B�=�&�=؝ >�k > y�=���=`��=,��=F�=���=H��=�H�=��=08�=���=ĕ�=fS�=ڝ�=���=���=�O>�q>��>4k>��=���=���=�t�=̈�=��=�   �   �=�M\=�Q=T#�<�j:�ჼ�����A+�AH���Q��[G�
�)�x������ �~:P��<�8=�8[=6ߍ=Pz�=���=���=�g�=��=b�=D��=���=F>�=���=N��=���=�}�=��=���=�=4��=��=j��=��=�`�=���=K�=��="��=���=* >�� >�7 >�H�=��=��=�&�=���=��=�   �   �%�=V&v=��4=�b�<H�8<큻������߼�)
�z��~����ۼ�߆���S�p D<H��<=6=}v=�͘=��=w�=���=P�=.��=���=���=T�=��=z��=ƴ�=2�=�H�=��=F��=;�=���=��=|��=~1�=���=�k�=~*�=N4�=h��=D��=��="��=��=ʂ�=�}�=n��=ܤ�=�X�=j³=�   �   X�=2(�=��Y=f=<@�<p�%<@�Һ�.�P��(ԓ����x�"� 9�@6<a�<A� =(�\=`�=��=J��=�!�=$��=��=R*�=��=H��=��=z��=6�=��=zE�=�b�=T3�=�m�=|��=�9�=Ok�=�F�=���=�I�=��=�N�=$d�=�6�=�=N�=`^�=���=�2�=.�=�i�=*��=��=IѼ=�   �   �
�=ą�=��=��L=U"=��<zw<���;`u"; �:@�>;�	<P��<�T�<�d=�Q=��=�4�=�2�=�7�=Z��=�j�=�3�=�!�=]�=l(�=���=��=��=R��=�v�=��=փ�=�ş=�y�=�=���=S1�=>��=���=�=M�=�=���=�f�=�7�=��=���=�Q�=$��=�,�=��=���=���=�   �   ,U�=�U�= m�=&E}=teP=��&=�{= ��<<��<м�<��<�b�<	�=��,=<�V=ᰁ=>5�=L��=S/�=���=.b�=@�=vb�=��=Vn�=@��=<��=���=u�=���=��=���=:Y�=,D�=HTt=�Ui=�Qf=|k=�px=X �=Ȓ=*Y�=ܰ=�S�=,��=��=�=Ҍ�=���=���=H��=��=���=���=�   �   �^�=~ٻ=U��=,��=ⶃ=��d=�4G=��0=60#=$?=KG%=��4=аL=H=k=R8�=�="�=�Ⱦ=V��=�R�=4��= ��=�9�=���= ��=&`�=�d�=�]�=�ػ=4��=́�=O��=�d=�0G=`�0=�+#=^:=�B%=��4=T�L=9k=r6�=t�=��=�Ǿ=^��=�Q�=���=���=�9�=���=D��=v`�=(e�=�   �   \��=�u�=Ƣ�=��=,��=�Z�=F�=TXt=�Yi=(Vf=|�k=�tx=`"�= ʒ=�Z�=�ݰ=U�=H��=ġ�=��=T��=��=��=H��=��=l��=��=xT�=�T�=�k�=dB}=4bP=��&=mw=���<���<���<���<�X�<U�=��,=H�V=��=�3�=	��=F.�=���=�a�=�?�=:b�=��=vn�=���=���=�   �   ���=ή�=H��=x�=,�=P��=�ǟ={�=��=��=:3�=��=b��=��=��=^��=���=�g�=b8�=���=&��=�Q�=H��=�,�=���=���=��=�	�=ℚ=��=�L=*=t�<xiw<@o�; '"; �~:�e>;X�<���<�K�<�`=HQ=@�=Z3�=�1�=�6�=���=j�=V3�=�!�=]�=�(�=^��=�   �   ���=��=��=wF�=�c�=�4�=o�=��=;�=�l�=�H�=4��=&K�=z��=�O�=@e�=�7�=��=�N�=�^�=��=
3�=.�=�i�=��=���=�м=��=b'�=��Y=�	=d:�<��%< )Ӻ�.��!���ݓ�����"� 4:��6<Y�<�� =�\=�=�~�=x��=$!�=���=���=8*�=2��=���="�=�   �   ���=��=r��=��=�I�=��=k��=><�=ϒ�=��=ʖ�=�2�=��=�l�=�+�=65�=4��=��=x��=���=:�= ��=�}�=h��=���=lX�=
³=_%�=%v=@�4=p^�<H�8<��x�����߼".
�������ۼ$膼@�S���C<���<::6=�zv=�̘=�=��=���=
�=��=���=��=��=�   �   �>�=��=ʗ�=F��=x~�=��=h��=��=(��=��=h��=��=�a�=���=�K�=���=���=8��=` >�� >8 >�H�= ��=��=�&�=d��=���=��=�L\=KP=H �<��:惼�����D+�dDH�f�Q��_G��)�ܯ�������}:���<6=�6[=Uލ=�y�="��=,��=dg�=̲�=d�=^��=���=�   �   �k >^y�=ަ�=���=���=��=\��=���=4I�=^�=�8�=N��=`��=�S�=Z��=J��=V��=�O>�q>ݎ>Kk>(��=���=���=�t�=���=���=D�=�mH=�<�u:<�6���м��'�8<Y�xx��z����w�,.X���&���μ�����	9<���<>.F=m�=���=["�=��=X��=8j�=@�=�&�=� >�   �   ��>�� >���= ��=.��=VP�=���=<�=���=@x�=���=&��=6D�=X{�=�(�=���=�|>p>X�>T�>�$>XG�=���=8��=���=tٽ=R2�=f
�=��;=x}�<p��;�cR�� ���B�vdv�������jR��2�u��4B��R � �S�@��; a�<z�8=k�=j՟=[#�=���=��=�4�=:��=�= >��>�   �   �>�>��>[m >x��=��=��=��=���=T��=d��=�r�=&��=��=J >�>u�>:�>�D>�>��>if>�o�=�"�=��=���=(�=yC�=���=T�g=�.0=2��<�ƌ<P�; �����@E�0Q�@���;D5�<F�<�V/=�Vf=Hٍ=1æ=Q=�=���="G�=Ԃ�=Н�=���=3>�^>�   �   �8>Ւ>�]>��=D�=4�=pQ�=�T�=�;�=��=t��=���=H\�=��=�8�='m>�>�F>o�>��>.�>LL>�k�=�R�=�=���=��=Op�=r�=�gk=�X4=�a�<���<X�< 㔹�����|뻐կ� ����<�k�<dD�<��3=�j=�e�=@�=!<�=��=���=���=.��=��=	>h>�   �   �%>�<>���=��=�"�=H��=ro�=L0�=r��=���=N��=&��=Ƅ�=`�=� �=5�=ov>��>-�>��>k >�� >^_�=���=�I�=h��=��=%�=��=غu=.�@=lP=���<�G<P�;�#��0�����z�;عK<<;�<k�=Fs@=��t=`�=���=�#�=<��=t,�=Ȁ�=���=�*�=j>�K>�   �   @c >�=�G�=���=�<�=���=j@�=��=
�=8��=��=��=�c�=��=�F�=��=���=�� >�>�>�>?z >�C�=ڽ�=2�=r��=��=HY�=#��=��=�S=
�"=�A�<Dě<��>< ��;��;�>�;8�C<���<p<�<��#=�T=�=-�=���=(��=��=i�=���=���=�Z�=�� >�� >�   �   ��=� �=���=Z�=���=L�=���=��=̕�=�4�= b�=�
�=� �=�=>��=6��=zR�=�G�=��=� >7� >���=�=���=��=v�=~Q�=d|�=�n�=�܍=4fm=�@=�=�M�<��<,��<X�~< g�<�\�<&��<�e=�/B=�o=�i�=i��=�C�=~��=�t�=�K�=�#�=��=�4�=$��=2[�=�   �   ��=�Z�=h��=(��=nm�=4��=�>�=S�=(��=T$�=j��=��=�x�=.��=��=���=H�=��=���=H|�=�4�=|��=���=�
�=�|�=��=���=A��=��=���=���=�[b=��<=�u={�=h�<�S�<�<�<0�=�3= �?=�qe=���=ȡ�=(��=3�=k��=���=���= ��=B�=���=��=��=�   �   ���=FI�=��=��=s��=���=�ɽ=i��=ʔ�=�Ҵ=#h�=x9�=��=�d�=��=
��=���=;�=�\�=���=O�=f|�=/�=�9�=z�=���=���=���=�T�=O\�=��=߃=��f=[J=<�4=�'=�x#=��(=I7=@�M=�pj=H܅=Jȗ=��=��=���=�%�=B��=��=xr�=� �=���=�W�=���=�   �   ���=��=_b�=[>�=�N�=dI�='ө=�x�=���=���=ky�=��=S �=h�=�0�="5�=�C�=���=Z��=l�=���=��=�d�=�E�=dq�=���=`��=bf�=*�=Z��=r��=V*�=c�=�~y=�g=R�[=�zX=.H]=��i=�H}=��=B��=��=�ָ=d�=���=��=l��=���=��=��=ؽ�=�E�=s�=�   �   ���=���=���=@c�=D5�=S"�=��=1�=̂�=0/�=�K�=்=���=��=��=f�=�n�=�+�=T��=TY�=b��=l��=S�=��=�;�=���=���=P��=s��=���=`d�=�6�=�#�=�=�2�=k��=�0�=VM�=a��=*��=H��=�=d�=eo�=�,�=ާ�=�Y�=���=���=S�=��=\;�=J��=��=�   �   �e�=2)�=V��==��=�(�=���=�{y=Pg=��[=HwX=�D]=��i=�E}=L�=��=��=�ո=��=T��=���="��=Ԙ�= ��=��=��=>F�=�s�=b��=��=Lc�=h?�=�O�=�J�=�ԩ=fz�=��=��=�z�=
�=��=��=�1�=6�=�D�=���=���=dl�=���=4��=�d�=�E�=$q�=h��=���=�   �   3��=	T�=D[�=p�=�݃=��f=�WJ=��4=��'=Cu#=��(= F7=f�M=6nj=*ۅ=TǗ=��=Z��=O��=h%�=���=d�=jr�=� �=���=�W�=��=P��=�I�=���=��=���=��=˽=���= ��=�Ӵ=ri�=�:�=��=�e�=���=���=���=�;�=F]�=���=TO�=�|�=/�=�9�=�y�=���=���=�   �   ���=��=���=v��= Yb=�<=�r=G�=���<xM�<�6�<G�=�0=��?=�oe=���=��=���=�2�=
��=R��=p��=��=N�=��=Z��=n��=���=4[�=��=���=Zn�=.��=�?�=i�=G��=x%�=���=���=�y�=��=���=x��=��=@��= ��=�|�=�4�=���=���=�
�=�|�=�=3��=�   �   �{�=�m�=�ۍ=dm=�@==H�<��<<��<��~<�a�<|W�<~��<�c=�-B=o=i�=ꛤ=WC�=/��=�t�=�K�=�#�=��=�4�=X��=�[�=���=T�=n��=�Z�=d��=�L�=���=n��=���=�5�=c�=��=��=��=��=Ң�=�R�=�G�=��=3� >M� >���= �=r��=Ҩ�=�u�= Q�=�   �   �X�=v��=�=2�S=��"=l=�<���<ض><���;޳;P,�;(|C<$��<F9�<�#=��T=��=�,�=v��=��=��=�h�=��=���=�Z�=�� >� >ic >`�=:H�=F��=(=�=R��=A�=���=�
�=���=���=��=�d�=���=G�=��=��=�� >�>7�>�>Dz >�C�=���=�1�=��=���=�   �   ��=���=��u=č@=�N=T��<��G< �;��#��K� X��o�;��K<<9�<��=�r@=$�t=*�=b��=�#�=*��=r,�=ʀ�=���=�*�=}>�K>�%>�<>��=f��=�"�=���=�o�=�0�=���=>��=���=���=,��=��=@!�=T5�=�v>��>?�>��>p >�� >P_�=���=�I�=(��=���=�   �    p�=�q�=�fk=�W4=t_�<x��<�< d��������� ۯ� �� �<�j�<�C�<԰3=tj=�e�==�="<�=��=���=���=>��=��=>v>�8>�>�]>L��=6D�=l�=�Q�=.U�=4<�=��=���= ��=v\�=B��=�8�=8m>�>�F>w�>��>4�>JL>�k�=�R�=��=P��=���=�   �   JC�=���=��g=N.0=R��<ƌ<���;@#�����HE��O�@ �P��; 6�<�F�<
W/=FWf=xٍ=\æ=m=�=���=:G�=��=��=���=#3>�^>�>�>�>^m >|��=��=��=��=���=X��=d��=�r�= ��=��=J >>q�>7�>�D>�>��>bf>�o�=�"�=���=}��=�=�   �   Dp�=�q�=�gk=�X4=�a�<���<��< ���Ї���v�`ί� ����<�m�<ZF�<�3=Zj=6f�=��=\<�=;��=���=���=R��=.��=>x>�8>�>�]>J��=0D�=d�=�Q�=$U�=,<�=��=���=���=l\�=4��=�8�=7m>�>�F>x�>��>9�>QL>�k�=�R�=�=x��=��=�   �   9�=/��="�u=��@=�P=,��<��G<���; �"� �������;�K<\>�<��=�t@=��t=��=���="$�=���=�,�=���= ��=�*�=�>�K>�%>�<>ތ�=^��=�"�=���=�o�=�0�=���=(��=���=���=��=��=8!�=R5�=�v>��>B�>��>y >�� >p_�=
��=�I�=z��='��=�   �   wY�=f��=<�=��S=�"=4D�<<Ǜ<�><���;@�;@O�;،C<쿞<z@�<��#=��T=��=�-�=K��=���=�=\i�=>��=���=�Z�=�� >
� >jc >^�=.H�=6��==�=<��=�@�=|��=�
�=���=���=|�=ld�=���=�F�=��=ܧ�=�� >�>7�>>Tz >�C�=���=(2�=���=;��=�   �   �|�= o�=Tݍ=Vgm=H@=L =\Q�<� �<���<�~<,l�<�a�<��<8h=�1B=�o=�j�=(��=^D�=��=`u�=VL�=*$�=��=5�=z��=�[�=���=J�=^��=�Z�=N��=�L�=x��=N��=���=n5�=�b�=��=��=��=β�=���=�R�=�G�=��=:� >W� >ޅ�=<�=���=:��=Jv�=�Q�=�   �   ���=A�=��=P��=<]b=��<=�w=��=�
�<hY�<�B�<��=Q6=��?=te=���=���=���=�3�=���=��=���=���=��=��=x��=���=���=,[�=��=ܘ�=8n�=��=�?�==�=��=J%�=`��=̰�=�y�=���=h��=f��=��=8��= ��=�|�=5�=Ĳ�=���=(�="}�=��=��=�   �   W��=jU�=�\�=h�=�߃=��f=b]J=��4=��'=�{#=��(=�K7=�M=dsj=�݅=dɗ=��=֧�=���=d&�=���=�=�r�=0�=��=$X�=��=N��=�I�=���=���=^��=���=�ʽ=��=�=�Ӵ=Bi�=�:�=��=�e�=���=���=f��=�;�=@]�=��=rO�=�|�=J/�=�9�=^z�=>��=��=�   �   �f�=�*�=��==��=B+�=n�=.�y=2g=�[=�}X=K]=��i=\K}=��=v��=��=�׸=5�=���=���=��=p��=p��=Z��=@��=bF�=�s�=^��=��=&c�=@?�=�O�=J�=Tԩ=(z�=ϩ�=Ƥ�=�z�=�	�=i�=l�=�1�=�5�=�D�=���=���=ll�=���=`��= e�=$F�=�q�= ��=���=�   �   ʶ�= ��=���=-e�=~7�=�$�=-�=�3�=���=42�=�N�=Ĳ�=���=���=8�=j�=Qp�=N-�=���=RZ�=(��= ��=nS�=�=�;�=���=���=F��=W��=���=4d�=`6�=�#�=��=`2�=(��=�0�=M�=(��=���=��=��=>�=Jo�=v,�=֧�=�Y�=���=���=LS�=�=�;�= ��=��=�   �   ؐ�=(	�=�c�=+@�=�P�=�K�=�թ=�{�=H��=J��=,|�=]�=��=��=�2�= 7�=�E�=V��=z��=�l�=X��=���=@e�="F�=�q�=���=d��=Tf�=�)�=2��=D��="*�=&�=L~y=g=��[=zX=�G]=T�i=,H}=d�=��=��=�ָ=U�=���=��=���=(��=N��=P��=V��=�F�= t�=�   �   ���=vJ�=v��=���=U��=ñ�=̽=ĥ�=<��=�Դ=�j�=�;�=��=�f�=���=���=@��=D<�=�]�=x��=�O�=�|�=`/�=�9�=@z�=��=���=���=�T�= \�=x�=�ރ=l�f=�ZJ=��4=��'=x#=n�(=�H7=ʫM=\pj=܅=*ȗ=��=僚=���=�%�=Z��=��=�r�="�=��=PX�=j��=�   �   ���=�[�=���=���=
o�=���=�@�=R�=:��=n&�=���=��=�z�=���=T��=0��=��=ʀ�=���=�|�=P5�=��=��="�=}�=��=���=*��=��=Z��=r��=<[b=L�<=2u=��=f�<�R�<�;�<��=-3=��?=\qe=���=���=��=3�=h��=���=���=R��=��=$��=���=���=�   �   ���=��=���=:[�=���=rM�=L��=0��=x��=\6�=�c�=v�=b�=��=���=d��=�S�=dH�=^�=e� >t� >��=N�=���=(��=v�=wQ�=N|�=�n�=�܍=�em=�@=K=�L�<��<H��<`�~<<f�<�[�<\��<�e=t/B=bo=�i�=U��=�C�=y��=�t�=L�=�#�=��=5�=���=�[�=�   �   �c >��=�H�=���=�=�=���=�A�=&��=V�=���=T��=(�=e�=,��=�G�=b �=T��=� >�>X�> >ez >�C�=���=2�=t��=��=8Y�=
��=��=��S=��"=A�<�Û<�>< ��;�;�;�;؂C<(��<�;�<��#=��T=��=�,�=���="��=��=i�=��=���=�Z�=�� >� >�   �   &>�<>��=���=F#�=���=:p�=1�=J��=���=&��=���=���=�=�!�=�5�=�v>��>[�>��>� >�� >�_�=��=�I�=p��=��=�=��=��u=��@=6P=(��< �G<��;�(#��4���y�;�K<�:�<I�=,s@=��t=P�=���=�#�=<��=�,�=܀�=���=�*�=�>�K>�   �   �8>�>�]>l��=TD�=��=�Q�=^U�=`<�=�=���=0��=�\�=n��=�8�=Jm>�>�F>��>��>>�>XL>l�=�R�=�=���=
��=Kp�=�q�=|gk=�X4=@a�<`��<�< ������� ~�p֯� �`�<Xk�<8D�<�3=tj=�e�=8�=<�=��=���=���=>��=,��=>|>�   �    Y>|�>�
>��>G� > ��=d��=���=���=H��=>I�=L��=.��=�} >��>"/>�b>�G>��>��>�>�>0��=rR�=އ�=���=x�=j��=c�=�~�=h��=�zv=^�T=��7=ZU!=B`=`�=��=~�!=� 8=`�T=fqv=c�=���=y>�=Nt�=�#�=Z��=0��=BO�=N��=�>�K>�0>�   �   �>��>�>(p>H& >t��=|��=�A�=l�=LU�=���=
a�=�a�=B��=zQ>��>��>��>�j>�H>�e>B�>���=�t�=���=h�=��='Q�=J�=���=��=��y=:.X=��;=��%=$�='=�=`�%=$<=ĎX=��y=j؎=.A�=�L�=�R�=^��=�|�=��=~�=���=	}>�(>`�>�   �   �>>��>{k>� >z4�=Hz�=�,�=�}�=^��=xn�=�#�=���=��= ��=6��=�T>	�>�>f�>!�>�>�h>j��=���=��=�\�=���=F��= �=�+�=X�=���=T�b=(G=��1=��$=T4 =��$=�2=l�G=Lec=@��=� �=��=g�=���=���=��=��=Z�=��=�L>.�>J]>�   �   ��>�� >X��=(��=��=��=7�=�;�=(�=���=��=rf�=���=���=�{�=8�=x� >�1>A.>�>�6>�>���=hu�=��=�~�=���=�s�=n��=���=���=��=�~s=�kY=�|E=\	9=n�4=��9= `F=��Z=��t=|��=L��=�Ӫ=�\�=|��=
�=h�=���=���=���=�� >�>`Z>�   �   . >0�=Pt�="L�=:�=,8�=���=L��=�+�=���=���=���=���=O�=�y�=���=>�=���=�J>v><5>�u>H��=69�= ��=�B�=��=�h�=��= �=�<�=Tڒ=���=�qq=T_=`�S=�P=WT=L`=s=��=���=��=܋�=A��=mH�=\H�=���=x��=��=��=5� >�->^� >�   �   ���="��=6��={�=�K�=L��=���=n��=���=�{�=*{�=Z��=�>�=��=���=���=�9�=��=T��=BQ >�� >�� >�D�=V�=���=8|�=�:�=�B�=d��=�Ǻ=*c�=�q�=���=�Ԇ=�&}=��r=<�o=��s=,�~=Hׇ=�Ӓ=���=Fr�=���=���=��=�3�=�!�=J �=��=���=���=] >ڎ�=�   �   0T�=���=`��=(H�=���=h�=j3�=��=h�=
��=��=k��=t��=�$�=�3�=X��=+�=j6�=�i�=@m�=Z��=��=���=���=(��=b��=�(�=ʯ�=p��=�Y�=���=�+�=�ڟ=�A�=9��=X��=�%�=���=V�=�z�=�F�=ר�=&��=1��=]��=�i�=|��=�
�=���=�D�=���=P��=:k�=ޗ�=�   �   `k�=���=���=��=$:�=�.�=�?�=���=�'�=�u�=�þ=���=���=�'�=�g�=�5�=V�=d��=^>�=���=,��=v��=L0�=��=��=J��=�B�=�_�=F?�=�V�=�2�=�i�=Z��=?�=���= �=� �=ĩ�=���=Υ�=�:�=0�=��=��=���=���=v�=�
�=/�=\c�=N��=8��=$e�=%�=�   �   p�=��=�O�=4��=���=1�=$�=Ű=���=Φ�=�!�=,�=�=w�=x��=a��=�C�=tR�=F��=���=~��=��=p_�=�2�=��=��=�Q�=��=���=~P�=���=t��=�1�=,�=+ư=���=觬=�"�=7�=夷=Z	�=B��=��=tD�=�R�=���=
��=���=<��=v_�=�2�=��=��=�Q�=�   �   _�=�>�=(V�=�1�=�h�=U��=�=�=f��=��=���=���=|��=Ѥ�=�9�=P/�=^��=l��=(��=@��="�=T
�=�.�=Rc�=V��=^��=\e�=x%�=�k�=.��=���=���=�:�=�/�=�@�=���=�(�=�v�=�ľ=���=���=\(�=�h�=\6�=��=ڗ�=�>�=���=^��=���=N0�=��=n�=��=�B�=�   �   J��=���=Y�=ꌷ=�*�=�ٟ=�@�=��=4��=�$�=p��=J��=�y�=�E�=��=z��=���=���=i�=0��=�
�=p��=�D�=���=l��=pk�=,��=�T�=z��=���=�H�=���=6�=H4�=̏�=i�=���=t�=N��=H��=�%�=t4�=���=�+�=�6�="j�=�m�=���=4��= ��=���=���=��=6(�=�   �   0B�=���=*Ǻ=eb�=�p�=Ƭ�=�ӆ=�$}=��r=�o=|�s=8�~=`և=�Ғ=A��=�q�=��=K��=���=F3�=v!�=* �=��=���=���=v >��=��=���=���=�{�=BL�=���=~��=2��=f��=b|�=�{�= ��=�?�=���=,��=X��=F:�=~��=���=`Q >� >�� >�D�=>�=���=�{�=�:�=�   �   xh�=]��=_�=:<�=�ْ=Լ�=�oq=x_=l�S=�P=LUT=TJ`=� s=X��=�=+�=j��=���=#H�= H�=v��=`��=���=��=@� >�->}� >S >\0�=�t�=�L�=��=�8�=*��=��=.,�=\��=v��=f��=���=�O�=Jz�=F��=��=��=�J>�>L5>�u>>��= 9�=���=JB�=���=�   �   )s�=���=��=�=-�=t}s=hjY={E=�9=��4=z�9=�^F=H�Z=t�t=���=���=kӪ=u\�=J��=��=�g�=��=���=���=�� >�>vZ>��>�� >���=���=�=~��=x7�=r<�=��=F��=���=�f�=��= ��=.|�=��=�� >�1>[.>!�>�6>�>���=Tu�=Z�=b~�=@��=�   �   ���=��=e+�=��=&��=D�b= G=h�1=`�$=;3 =��$=�~2=��G=�dc=���=� �=��=�f�=���=h��=��=��=X�="��=�L><�>X]>�>>>�k>� >�4�=�z�=0-�=�}�=���=�n�=$�=��=T��=D��=v��=�T>%�>�>u�>+�>
�>�h>d��=���=İ�=Z\�=t��=�   �   �P�=�=m��=k�=ޫy=�-X=�;=߈%=y�=r&=:=�%=�<=��X=��y=V؎=$A�=�L�=�R�=\��=�|�=��=~�=���=}>�(>j�>�>�>�>;p>Z& >���=���=�A�=Hl�=|U�=���=2a�=�a�=f��=�Q>ŷ>��>��>�j>�H>�e>?�>���=�t�=���=B�=��=�   �   J��=H�=�~�=F��=�zv=*�T=x�7=4U!=.`=X�=�=��!=8=��T=�qv=2c�= �=�>�=jt�=�#�=n��=@��=PO�=X��=�>�K>�0>Y>�>�
>��>I� >"��=b��=��=���=J��=@I�=L��=*��=�} >��>#/>�b>�G>��>��>�>�>(��=hR�=̇�=���=�w�=�   �   $Q�=E�=���=��=��y=X.X=؄;=҉%=u�=}'=8=�%=�<=d�X=p�y=�؎=pA�=M�=S�=���=�|�=��=~�=���=}>�(>l�>�> �>�>;p>X& >���=���=�A�=@l�=rU�=���=,a�=�a�=\��=�Q>��>��>��>�j>�H>�e>I�>���=�t�=���=d�=��=�   �   Y��=�=�+�=��=؇�=Եb=�G=@�1=M�$=;5 =��$=�2=`�G=Jfc=���=n!�=P�=Vg�=$��=���=*�=��=��=>��=M>B�>_]>�>>>�k>� >�4�=�z�=$-�=�}�=���=�n�=�#�=��=B��=8��=j��=�T> �>�>x�>-�>�>�h>z��=��=��=�\�=���=�   �   �s�=���=���=إ�=4�=�s=�lY=�}E=�
9=��4=J�9=�aF=ȌZ=ڧt=��=���=AԪ="]�=���=P�=Xh�=8��=���=���=�� >�>|Z>��>�� >���=z��=��=h��=f7�=X<�=��=0��=x��=�f�=��=
��=|�=��=�� >�1>Z.>$�>�6>>ƿ�=�u�=��=�~�=���=�   �   i�=(��=M�=V=�=�ڒ=:��=�rq=�_=вS=fP=�XT=�M`=�s=̙�=D��=X�=p��=���=�H�=�H�=��=���=B��=T��=Q� >�->�� >S >V0�=�t�=�L�=��=�8�=��=ԍ�=,�=<��=X��=D��=p��=�O�=2z�=:��=��=
��=�J>�>U5>�u>h��=\9�=��=�B�=��=�   �   �B�=���=8Ⱥ=�c�=@r�=X��=BՆ=`(}=d�r=�o=d�s=��~=(؇=jԒ=�=�r�=?��=>��=d��=�3�=�!�=� �=��=���=��=� >(��=
��=���=���=�{�=*L�=��=\��=��=D��=8|�=�{�=���=�?�=p��=��=N��=6:�=n��=���=bQ >� >�� >�D�=��=��=h|�=0;�=�   �   ��=���=4Z�=A��=T,�=T۟=�B�=
��=:��=�&�=}��=I�=�{�={G�=���=���=֞�=���=�i�=��=8�=��=.E�=$��=���=�k�=<��=�T�=h��=���=�H�=���=�=4�=���=�h�=���=L�=&��= ��=v%�=X4�=ޯ�=x+�=�6�=j�=�m�=���=P��=0��=���=X��=���=�(�=�   �   �_�=�?�=RW�= 3�=<j�=��=�?�=e��=� �=��=���=��=���=s;�=�0�=���=���=2��=��=��=�
�=p/�=�c�=���=���=xe�=~%�=�k�=��=~��=���=�:�=X/�=�@�=���=i(�=�v�=lľ=���=Z��=3(�=�h�=B6�=��=Η�=�>�=���=p��=���=�0�=N��=��=���=,C�=�   �   @	�=��=�P�=���=��=�2�=��=�ư=���=ר�=�#�=$�=˥�=-
�=��=���=E�=zS�=(��=r��=��=���=�_�= 3�=��= �=�Q�=��=���=^P�=���=P��=�1�=��=�Ű=o��=���=f"�=�=���=/	�="��=���=VD�=�R�=���=��=���=^��=�_�=3�=��=*�=6R�=�   �   (l�=���=��=Z��=�;�=,0�=�A�=���=l)�=�w�=wž=���=R��=)�=ti�=�6�=|�=X��=0?�=V��=���=���=�0�=L��=��=`��=�B�=�_�=(?�=�V�=n2�=oi�=)��=�>�=N��=��=y �=���=Z��=���=n:�=�/�=���=���=���=���=t�=�
�=</�=�c�=���=���=�e�=�%�=�   �   �T�=���=`��=TI�=8��=��=�4�=���=�i�=���=<	�=��=��=D&�=5�=���=,�=F7�=�j�=�m�=���=x��=D��=���=D��=r��=�(�=���=Z��=�Y�=���=�+�=vڟ=�A�=���=#��=�%�=T��=$�=�z�=pF�=���=��=��=O��=vi�=|��=�
�=���=E�=��=���=�k�=v��=�   �   X��=���=��=|�=�L�=���=��=Җ�=��=}�=�|�=���=F@�=$��=���=���=�:�=���= ��=�Q >)� >�� >�D�=~�= ��=B|�=�:�=�B�=K��=�Ǻ=c�=�q�=���=aԆ=z&}=T�r=ƺo=(�s=̨~=ׇ=nӒ=ښ�=*r�=���=���=��=�3�=�!�=^ �=��=���=&��=� >\��=�   �   p >�0�=u�=�L�=,�=09�=���=v��=�,�=���= ��=��=��=P�=�z�=���=��=f��=K>�>i5>�u>z��=T9�=��=�B�=��=�h�=ϱ�=��=�<�=0ڒ=���=2qq=�_= �S=�P=�VT=�K`=�s=昅=p��=��=Ƌ�=0��=bH�=XH�=���=���=$��=F��=T� >�->�� >�   �   �>�� >���=Ћ�=X�=���=�7�=�<�=�=���=���=Tg�=���=~��=�|�=��=�� >�1>y.>>�>�6>>п�=�u�=��=�~�=���=�s�=Z��=��=t��=��=�~s=�kY=`|E=	9=(�4=��9=�_F=<�Z=P�t=c��=6��=�Ӫ=�\�=t��=�=h�=
��=���=���=�� >�>�Z>�   �   �>>֊>�k>� >�4�=�z�=p-�= ~�=���=o�=H$�=Z��=���=���=���=U>>�>/�>��>C�>�>�h>���=
��=��=�\�=���=@��=��=�+�=F�=���= �b=�G=V�1=P�$=4 =��$=�2=2�G=(ec=1��=� �=��=�f�=���=~��=��=��=j�=6��=M>I�>h]>�   �   �>	�>*�>Gp>g& >���=���=B�=hl�=�U�=���=Ta�=�a�=���=�Q>ҷ>��>��>�j>�H>�e>K�>���=�t�=���=d�=��=$Q�=D�=���=��=p�y=.X=|�;=n�%=��=�&=�=J�%=<=��X=��y=b؎=&A�=�L�=�R�=\��=�|�=��=~�=���=}>�(>r�>�   �   �>jY>��>��>�>= >
> >^�=4��=>��=�0�=� >l� >�>��>T�>��>Lh>d�>��>c�>{>|d>�#�=L�=�f�=l�=�:�=��="\�=���="�=LК=63�=T��=VO�=�Ƀ=�g�=�	�=�a�=\��=",�=�h�=j�=��=���=P}�=E�=���=
��=3� >��>��>ڑ>�   �   Uy>�>\`>4x>d>�� >N��=<k�=���=ҵ�=�8�=G�=|g >Y>Be>�t>�i>i$>��>k>/�>�k>,c>.>�=48�=��=��=t��=���= *�= u�=�2�=3 �=N~�=~@�= ��=2=�=�׆=Go�=D��=�-�=�G�==d�=~�=M�=x�=���=ʢ�=N��=P��=ܓ >܈>k�>�i>�   �   ��>P>fu>�k>DU >Ğ�=���=���=���=���=8X�=4z�=� �=� >~;>Qg>�|>QZ>��>��>�h>�=>�^>���=���=<��=�!�= f�=���=\��=�5�=U�=*~�=�K�=�K�=��=��=�=^��=��=�Ɵ=.��=�F�=Gj�=tl�=���=�_�=���=n��=�.�=� >e>]}>�>�   �   ��>Z>�� >\m�=���=�~�=�}�=��=�-�=x�=��=��=���=��=x��=�� >#�>D>C�>�>��>��>�U>���=���=..�=P-�=8 �=��=S�=^��=0[�=z�=�`�=)=���=�M�=�ґ=@�=`̜=膥=��=��=�l�=D��=r��=>��=�f�=���=���=�� >�)>|�>�.>�   �   �s>W >X��=2��=V��=���=�}�=N��=b��=*��=-�=f��=@��=�r�=���=Թ�=b��=lQ>�c>�>�>��>^D>��=��=�#�=|��=tq�=�%�=8X�=�u�=���=Gr�=�_�=�>�=s�=�<�=��=:��=��={�=��=���=E��=�P�=�b�=H��=��=�L�=��=« >B�>�N>�%>�   �   օ�=,}�=��=t�=&W�= ��=��=\��= ��=�_�=^�=��=hI�=�v�= �=R��= ��=�W�=�� >�>&'>� >z&>�!�=��=�p�=|�=���=~,�=�R�=ie�=nٽ=�*�=&ԭ=tE�=7ؤ=�ƣ=�"�=,Ѩ=���=d�=�=1�=x��=��=
��=��=(2�= �=�f�=� >�h>Nt>� >�   �   Ҝ�=���=f*�=�{�=X��=���=PG�=V��=�'�=���=X��=D��=���=(I�=���=�F�=���=�]�=X1�=� >M	>�Z>�� >ҹ�=�
�= ��=<��=Z�=���=@��=��=Ƌ�=ʾ=�>�=�M�={F�=�\�=���=,��=4"�=*Կ=���=�$�=���=҈�=���=V��=��=P��=�E�=:� >i� >�q >4��=�   �   �F�=LI�=���=4#�=���=ذ�=���=,e�=ƈ�=��=��=,@�=^��=�$�=�F�=���=�p�=T��=���=���=���=�� >�� >�! >H��= ��=�>�=���=��=���=P'�=���=��=e!�=]Ѿ=�1�=;o�=s��=���=�&�=>�=��=�u�=~)�=8��=ĵ�=d��=>��=е�=- >� >?B >��=�w�=�   �   0��=��=���= F�=���=H��= �=NR�=��=fz�=؃�=7!�=�$�=M�=|K�=��=0n�=>��=���= ��=���=��=l >�Z >X�=�$�=���=���=J��=��=�F�=0��=���=��=S�=R�=/{�=���=�!�=q%�=�M�=L�=���=�n�=���="��=Z��=���=
��=l >�Z ><�=�$�=f��=�   �   ���=���=j��=�&�=��=Z��=� �=�о=
1�=qn�=���=ꍿ=�%�=��=��=@u�=)�=޲�=x��=$��=��=���=( >� >KB >��=�w�=8G�=�I�=r��=�#�=���=x��=H��=�e�=~��=��=���=�@�=��=�%�=2G�=.��=�p�=���=J��=ʣ�=Č�=� >�� >�! >*��=Ҏ�=N>�=�   �   �=L��=���=�=��=eɾ=>�=�L�=�E�=�[�=�=u�=�!�=�ӿ=���=x$�=d��=|��=l��=��=��=6��=�E�==� >t� >	r >l��= ��=R��=�*�=8|�=���=���=�G�=���=�(�=B��=���=��=2��=�I�=��=*G�=��=.^�=�1�=� >`	>[>�� >Ĺ�=�
�=���=���=�   �   ���= ,�=R�=�d�=�ؽ=�)�=tӭ=�D�=�פ=@ƣ="�=�Ш=䏮=��=n��=�0�=��=���=���=|�=2�=�=�f�=� >�h>_t>*� >��=z}�=x��=��=�W�=~��=L�=���=���=Z`�=��=���=�I�=w�=t�=���=Z��=�W�=� >(�>5'>� >y&>�!�=��=�p�=>�=�   �   *q�=^%�=�W�=du�=;��=�q�=_�=M>�=nr�= <�=i��=���=0�=�=���=|��=��=XP�=zb�=��=ě�=�L�=؍�=ë >J�>�N>�%>t>2W >���=���=���=4��=N~�=ĺ�=ط�=���=�-�=ڞ�=���=,s�=܁�=(��=���=�Q>�c>>>��>_D>��=f�=�#�=H��=�   �   ���=���=�R�=���=�Z�=�=`�=���=6��=:M�=Bґ=��=�˜=���=���=k�=�l�=��=H��=��=�f�=���=���=�� >�)>��>�.>��>w>�� >�m�=<��=6�=$~�=�=J.�=��=f��=l��=���=H�=���=�� >@�>Z>W�>�>��>��>�U>���=���=.�= -�=�   �   �e�=^��=��=u5�=�T�=�}�=ZK�=bK�=@�=>�=��=��=Ж�=EƟ=���=�F�="j�=Wl�=���=�_�=��=l��=�.�=� >e>h}>�>��>P>wu>�k>^U >���=���=2��=4��=���=zX�=pz�=!�=� >�;>hg>�|>aZ>�>��>�h>�=>�^>���=���="��=�!�=�   �   T��=���=�)�=�t�=�2�=���=~�=H@�=ɼ�=�<�=�׆=#o�="��=�-�=�G�=0d�=r�=�L�=t�=���=Ģ�=P��=P��=� >ވ>n�>�i>]y>�>f`>Dx>r>� >j��=Zk�=���=���=�8�=8G�=�g >(Y>Me>�t>�i>q$>��>k>3�>�k>,c>(>�= 8�=���=��=�   �   �:�=��=\�=���=�!�=>К=&3�=J��=RO�=�Ƀ=�g�=
�=�a�=l��=2,�=i�=~�=��=΁�=V}�=E�=���=��=6� >�>��>ۑ>�>mY>��>��>�>> >> > ^�=6��=>��=�0�=� >i� >�>��>S�>��>Lh>d�>��>b�> {>zd>�#�=<�=�f�=l�=�   �   t��=���=�)�=!u�=�2�=B �=a~�=�@�=��=T=�=؆=wo�=s��=�-�=�G�=jd�=��=+M�=��=���=ޢ�=d��=d��=� >�>s�>�i>ay>�>g`>Ax>n>� >h��=Tk�=���=��=�8�=.G�=�g >&Y>Je>�t>�i>o$>��>k>2�>�k>1c>0>�=28�=��=��=�   �   f�=���=m��=�5�==U�=T~�=�K�=�K�=��=��=V�=���=d��=�Ɵ=v��=G�=�j�=�l�=��=�_�=��=���=�.�=%� >$e>l}>�>��>P>xu>�k>[U >���=���="��=*��=���=nX�=dz�=!�=� >�;>cg>�|>`Z>�>��>�h>�=>�^>���=���=F��=�!�=�   �   R �=9��=BS�=���=l[�=��=�`�=�=��="N�=.ӑ=��=�̜=P��=p��=�=(m�=���=���=n��=g�=���= ��=�� >�)>��>�.>��>q>�� >�m�=,��=(�=~�=��=6.�=��=R��=X��=��=:�=���=�� >9�>X>U�>�>��>��>�U>���=���=D.�=h-�=�   �   �q�=�%�=lX�="v�=��=�r�=`�=\?�=�s�="=�=���=Į�=:�=��=���=K��=���=�P�=�b�=���=��=�L�=��=֫ >V�>�N>�%>t>-W >���=~��=���=��=4~�=���=���=���=p-�=�=���=s�=΁�=��=���=�Q>�c>>>��>lD>4��=��=�#�=���=�   �   (��=�,�=�R�=�e�=�ٽ=�*�=�ԭ=�E�=�ؤ=�ǣ=W#�=�Ѩ=��=��=r��=�1�=���=\��=\��=��=f2�=T�=�f�=1� >�h>it>0� >��=p}�=h��=��=�W�=f��=.�=���=r��=8`�=��=|��=�I�=�v�=Z�=���=J��=�W�=� >'�>>'>� >�&>�!�=��=�p�=��=�   �   ��=���=���=�=.��=�ʾ=Q?�=HN�=G�=0]�=O��=���=�"�=�Կ=��=t%�=D��=2��=��=���=�=���=�E�=S� >�� >r >r��=��=F��=�*�=(|�=���=l��=�G�=ԯ�=d(�=��=ܝ�=�=��=�I�=��=G�=���=^�=�1�=� >f	>[>�� >���=�=J��=l��=�   �   $��=8��=8��=�'�=��=���=�!�=�Ѿ=l2�=�o�=��=D��="'�=��=���=@v�=�)�=���=��=���=~��=��=H >*� >ZB >$��=�w�=2G�=�I�=Z��=�#�=h��=V��=$��=�e�=V��=Y�=���=�@�=޶�=p%�=G�=��=�p�=���=F��=ȣ�=Ԍ�=� >�� >
" >p��=4��=�>�=�   �   £�=���=l��=G�=���=h��=<�=�S�=��=�{�=8��=�"�=	&�=JN�=�L�=��=o�=���=t��=���=���=D��=4l >�Z >t�=�$�=���=~��=6��= ��=�F�=��=���=��=�R�=&�={�=p��=�!�=K%�=�M�=�K�=���=�n�=���=��=\��=���="��=+l >�Z >��=%�=���=�   �   tG�=�I�=���=$�=��=��=΄�=ff�=��=�=d��=pA�=���=&�=�G�=���=Vq�=��=���=��=��=(� >û >" >`��=��=�>�=���=ޡ�=���=<'�=s��=���=;!�=/Ѿ=�1�=o�=G��=|��=f&�=�=���=�u�=l)�=.��=���=\��=H��=��=@ >(� >bB >D��=&x�=�   �   X��=���=+�=�|�=H��=���=dH�=t��=)�=���=���=l��=���=(J�=v��=�G�=h��=|^�=�1�=  >}	>[>�� >���=�=*��=:��=N�=���="��=��=���=�ɾ=�>�=�M�=OF�=k\�=���=��="�=	Կ=i��=�$�=���=Ĉ�=���=T��=��=d��=�E�=Q� >�� >"r >���=�   �   H��=�}�=���=0�=�W�=���=��=Z��=��=�`�=f�=��=ZJ�=xw�=��=��=���=DX�=:� >@�>N'>� >�&>�!�=��=�p�=z�=��=n,�=bR�=Re�=Kٽ=r*�=�ӭ=FE�=ؤ=�ƣ=�"�=Ѩ=a��=A�=յ�=
1�=d��=���= ��=��=02�=*�=�f�=/� > i>st>B� >�   �   t>JW >���=���=��=���=�~�=$��=6��=��=�-�=>��=
��=�s�=2��=r��=���=�Q>�c>'>>��>rD>2��=��=�#�=x��=hq�=�%�= X�=�u�=���='r�={_�=�>�=�r�=z<�=⮚=��=��=^�=��=���=5��=�P�=�b�=B��=��=�L�=���=ҫ >X�>�N>�%>�   �   ��>�>�� >�m�=p��=v�=l~�=T�=�.�=$�=���=���=D��=��= ��=İ >\�>s>i�>�>��>�>�U>���=���=2.�=L-�=0 �=��=S�=J��=[�=`�=j`�==���=�M�=�ґ=$�=B̜=Ά�=���=��=�l�=8��=j��=:��=�f�=���=��=�� >�)>��>�.>�   �   ��>$P>�u>�k>uU >$��=���=f��=h��=���=�X�=�z�=H!�=� >�;>zg>�|>uZ>�>��>�h>�=>�^>���=���=@��=�!�=�e�=���=Q��=�5�=U�=~�=�K�=�K�=��=��=��=L��= ��=vƟ=$��=�F�=:j�=ll�=���=�_�=���=r��=�.�=!� >%e>l}>�>�   �   ey>�>o`>Kx>|>� >���=zk�=���=��=�8�=PG�=�g >4Y>Ye>�t>�i>x$>�>k><�>�k>3c>0>�=68�=��=��=t��=���=�)�=u�=�2�=+ �=C~�=t@�=���= =�=�׆=:o�=8��=�-�=�G�=8d�=v�=�L�=v�=���=Ģ�=T��=X��=� >�>u�>�i>�   �   ��>Xu>��>�Q>��>��> d>� >M� >[� >�� >yG>^�>?�>@H>�	>��>�:>�y>\^>��>��>@>U) >��=\��=���=`��=�_�=Z��=���=�b�=ǻ=S]�=B��=���=̀�=���=���=���=D�=�t�=���=�i�=T�=Hd�=�#�=��=@0�=�F�=��>�(>�">�>�   �   x�>�C>�>q>�U>�>J>�� >�] >�U >� >3� >Հ>�5>e�>�>|>�>dP>�>>D�>��>�?>~3 >A�=&�=r�=�<�=<��=��=�k�=j�=���=:9�=�k�=�p�=�t�=���=P��=He�=i��=�3�=�k�=���=d��=���=Tx�=�]�=^�=<a�=��>r >`>�>�   �   �>��>�>xF>�w>�� >~ >� �=��=(��=J��=���=�� >�D>
>:�>3�>q>r�>��>�>΢>�>>P >��=4��=���=�[�=�3�=0��=�I�=d6�=d�=���=$�=4�=5B�=�M�=rE�=���=�!�=od�=p`�=��=z�=��=^r�=l�=|��=��=+�>>>8�>L+>�   �   0V>"�>7�>,># >�V�=\��=V��=��=���=�j�=�\�=���=\y�=մ >�>-�>�{>n>�H>m>�l>�9>�z ><f�=<��=4`�= *�=�f�=,W�=dJ�=���==��=�̼=�_�=��=���=Wĵ= ��=i�=���=���=}��=Hs�=0^�=���=�=�O�=$��= >к>I�>hx>*�>�   �   �P>�z>_o >��=.N�=D4�=to�= �=X^�=�8�=���=��=�X�=�U�=<��=,��=1&>�/>��>wy>��>B>M->� >�M�=h<�=BE�=���=�S�=���=�G�=��=��=v(�=(	�=\~�=¯�=ڨ�=�X�=N��=��=Ï�=���=n�=�z�=0��=��=���=���=�U >��>�>/�>X�>�   �   6>���=Z5�=h�=��=.%�=�	�=�y�=��=6]�=���=*�=���= C�=���=��=&��=�� >!�>x>j�>9�>>S� >[�=���=���=Ds�=z��=��=@�=:z�=���=N��=��=�t�=��=���=�'�=T�=x#�=(�=���=`p�=3�=@��=��=v��=��=� >�>�K>T>1�>�   �   6�=VH�=T�=(��=~P�=,R�=���=(��=���=L��=b+�=��=��=�h�=>��=���=L�=��=�- >cJ>� >>>��>�>�~�=L��=��=��=���=(��=�b�=^v�=j�=/��=�<�=D,�=8��=j�=F��=k?�=F��=@�=�'�=G�=�W�=��=�P�=���= ]�=5� >��>l�>K�>/� >�   �   ���=zZ�=c�=hV�=Vo�=��=���=���=�g�=B�=���=U�=���=h��=���=���=���=�w�= �=���=�>:�>*�>�R>IT >���=Ҿ�=|�=��=J��=�=j��=��= �=��=�I�=���=׏�=���=D��=���=���=V��=xb�=*��=���=�5�=���= _ >CD>i�>�l>&� >��=�   �   (��=�1�=D�=`��=�0�=��=6��=�=:w�=�	�=���=z��=\h�=�=`?�= ��=��=j'�=�k�=z�=� >�>��>�}>�� >��=Rt�=h��=�1�=��=���=1�=f�=���=��=�w�=0
�=R��=���=�h�=��=�?�=`��=6��=�'�=�k�=��=� >�>��>�}>�� >���=(t�=�   �   >�=���=��=��=���=��=��=h�=8I�=p��=L��=��=���=F��="��=���=$b�=��=���=^5�=���=�^ >>D>l�>�l>8� >��=���=�Z�=rc�=�V�=�o�=���=��=:��=8h�=��=@��=�U�=��=���= ��=Z��=��=.x�=L �=���=�>B�>+�>�R>?T >~��=���=�   �   ���=���=Д�=Rb�=�u�=��=���=s<�=�+�=���=�i�=ʱ�=�>�=���=�?�=^'�=�F�=�W�=t�=�P�=���=�\�=0� >��>t�>Y�>D� >J6�=�H�=��=~��=�P�=�R�=X��=���=r��=Ĕ�=�+�=���=���=�h�=���=H��=XL�=R��=�- >uJ>� >>> �>�>|~�=*��=T�=�   �   s�=6��=���=��=�y�=#��=و�=���=*t�=f��=���=L'�=��=#�=��=���=p�=�2�=��=��=\��=��=� >�>�K>'T>D�>O>&��=�5�=Rh�=v��=�%�=
�=�y�=|��=�]�=���=��=��=zC�=D��=d��=j��=� >9�>x>w�>?�>>Q� >�Z�=���=���=�   �   Ɛ�=`S�=h��=�G�=.�=���=(�=��=�}�=V��=s��=3X�=��=p�=u��=n��=4�=�z�=��=d�=���=���=�U >��>�>7�>f�>�P>�z>|o >(��=vN�=�4�=�o�=\ �=�^�=L9�=Z��=j��=>Y�= V�=~��=l��=P&>�/>��>�y>�>G>K->� >�M�=H<�=E�=�   �   �)�=�f�=�V�=#J�=f��=��=�̼=�_�=¢�=T��=�õ=՜�="�=W��=`��=D��=s�=^�=���=��=zO�=��= >Һ>M�>ox>8�>AV>2�>N�>G>@ >W�=���=���=��=���=�j�=�\�=п�=�y�=� >,�>C�>�{>|>�H>u>�l>�9>�z >"f�=&��=`�=�   �   �[�=�3�=���=aI�=(6�=.�=i��=��=�3�=�A�={M�==E�=���=l!�=Ld�=M`�= ��=`�=��=Hr�=b�=|��=��=-�>A>?�>T+>�>ͯ>>�F>�w>ֳ >� >!�=��=Z��=z��=(��=�� >�D>>L�>E�>)q>{�>��>�>Ң>�>>P >ֲ�="��=���=�   �   �<�=$��=��=�k�=C�=���=9�=~k�=�p�=�t�=���=:��=3e�=Q��=�3�=�k�=���=`��=���=Px�=�]�=^�=@a�=��>s >f>�>~�>�C>��>x>�U>�>Q>�� >�] >�U >�� >?� >��>�5>m�>!�>|>�>kP>�>>I�>��>�?>z3 >�@�=�=b�=�   �   R��=�_�=N��=���=�b�=ǻ=I]�==��=���=π�=���=���=���=H�=u�=���=j�=`�=Rd�=�#�=��=H0�=�F�=��>�(>�">�>��>Xu>��>�Q>��>��>�c>� >N� >[� >�� >yG>^�>?�>?H>�	>��>�:>�y>[^>��>��>@>T) >��=T��=���=�   �   �<�=<��=��=�k�=r�=��=J9�=�k�=q�=u�=ȅ�=p��=ee�=���=�3�=l�=���=|��=���=bx�=�]�=^�=Ha�=��>u >h>�>}�>�C>��>w>�U>�>O>�� >�] >�U >�� ><� >܀>�5>j�> �>|>�>kP>�>>H�>�>�?>3 >A�=(�=r�=�   �   �[�=
4�=8��=�I�=u6�=��=ɿ�=F�=,4�=cB�=�M�=�E�=���=�!�=�d�=�`�=F��=��= �=tr�=��=���= ��=4�>D>B�>X+>�>ͯ>>�F>�w>ӳ >� >!�=��=N��=n��= ��=�� >�D>>L�>D�>(q>y�>��>�>Ԣ>�>>P >��=:��=���=�   �   4*�= g�=HW�=�J�=ݚ�=h��=ͼ=+`�=X��=���=�ĵ=h��=��=���=���=���=|s�=^^�=���=(�=�O�=>��= >ۺ>T�>ux>9�>@V>3�>K�>B>: >W�=���=���=��=���=�j�=�\�=¿�=�y�=� >&�>@�>�{>|>�H>x>�l>�9>�z >Ff�=N��=D`�=�   �   ��=�S�=���=H�=��=B��=�(�=p	�=�~�=��=0��=�X�=���=�=��=���=��= {�=^��=��=���=���=�U >��>%�>?�>k�>�P>�z>wo > ��=jN�=�4�=�o�=H �=�^�=89�=B��=T��=*Y�=�U�=r��=\��=J&>�/>��>�y>	�>M>T->�� >�M�=�<�=dE�=�   �   hs�=���=F��=|�=yz�=Ո�=���=R��=u�=B��=^��=(�=��=�#�=|�=F��=�p�=P3�=x��=<��=���=��=�� >�>�K>0T>I�>M>��=�5�=Fh�=`��=x%�=
�=�y�=d��=�]�=���=z�=���=fC�=6��=Z��=^��=� >6�>x>|�>G�>>a� >,[�=��=։�=�   �   ��=���=X��=�b�=�v�=��=���=P=�=�,�=���=~j�=���=�?�=���=`@�=
(�=XG�="X�=��=�P�=���=(]�=H� >��>}�>b�>G� >@6�=�H�=��=p��=�P�=zR�=:��=|��=T��=���=�+�=d��=h��=�h�=���=4��=HL�=F��=�- >tJ>� >%>>�>�>�~�=p��=��=�   �   ��=:��=���=H�=���=L�=|�=L�=J�=d��=A��=���=���=��=��=���=�b�=h��=���=�5�= ��=_ >VD>|�>�l>?� >��=���=�Z�=\c�=�V�=�o�=p��=���=��=h�=��=��=xU�= ��=���=��=D��=���= x�=@ �=���=>M�>:�>�R>[T >Ħ�=���=�   �   ���=2�=��=��=T1�=��=��= �=&x�=�
�=���=f��=8i�=��= @�=���=���=�'�=l�=��=� >�>Ǌ>�}>�� >��=Xt�=`��=�1�=��=���=�0�=H�=���=��=�w�=

�=.��=ޘ�=�h�=t�=�?�=J��=&��=�'�=�k�=��=� >�>��>�}>�� >*��=�t�=�   �   " �=�Z�=�c�=W�=p�=���=p��=���=�h�=&�=���=�U�=v��=*��=V��=���=T��=hx�=� �=���=>V�>@�>�R>ST >���=Ծ�=t�=���=2��=��=P��=��=�=��=�I�=���=���=h��=(��=���=t��=B��=hb�=��=���=�5�=���=_ >OD>|�>�l>I� >�=�   �   r6�=�H�=��=���=,Q�=�R�=���=���=���=��=6,�=ؓ�=ڳ�=Ji�=��=���=�L�=���=�- >�J>� >1>>�>�>�~�=V��=��=֭�=���=��=�b�=Fv�=N�=��=�<�=",�=��=�i�=$��=M?�=(��=�?�=�'�=�F�=�W�=��=�P�=���=]�=B� >��>��>k�>X� >�   �   d>T��=�5�=�h�=���=�%�=h
�=Nz�=̐�=�]�=H��=��=P��=�C�=���=���=���=*� >N�>*x>��>Q�>>_� >[�=���=���=<s�=l��=��=.�="z�=r��=0��=���=�t�=¼�=ܨ�=�'�=:�=^#�=�=��=Vp�=3�=6��=��=~��=��=� >�>�K>9T>X�>�   �   �P>�z>�o >\��=�N�=�4�=p�=� �=�^�=�9�=���=���=�Y�=<V�=���=���=i&>0>��>�y>�>V>Z->�� >�M�=h<�=BE�=��=�S�=���=�G�=v�=��=\(�=
	�=@~�=���=���=yX�=4��=��=���=���=b�=�z�=&��=��=���=���=�U >��>(�>E�>w�>�   �   LV>D�>]�>Y>U >@W�=���=ʹ�=�=��=.k�= ]�= ��=�y�=� >?�>U�>�{>�>�H>�>�l>�9>�z >>f�=>��=0`�=*�=�f�= W�=TJ�=���='��=�̼=�_�=��=���==ĵ=
��=Q�=���=���=m��=:s�=(^�=���=�=�O�=&��= >ں>V�>{x>B�>�   �   �>د>>�F>�w>� >� >>!�=:��=���=���=P��=�� >E>)>Y�>N�>2q>��>��>�>آ>�>>P >��=6��=���=�[�=�3�="��=�I�=T6�=X�=���=�=�3�=#B�=�M�=fE�=���=�!�=id�=h`�=��=p�=��=Zr�=l�=���=��=3�>G>C�>_+>�   �   ��>�C>�>�>�U>%�>[>�� >�] >�U >� >F� >�>�5>u�>'�>|>�>pP>�>>J�>�>�?>3 >A�=$�=n�=�<�=6��=��=�k�=b�=���=29�=�k�=�p�=�t�=���=F��=>e�=_��=�3�=�k�=���=`��=���=Tx�=�]�=^�=Ba�=��>u >j>��>�   �   M�>�[>��>��>�>Ճ>r>k�>��> �>�>��>_>��>�l>��>hv>5�>�>��>Ӎ>��>��>�*><��=� �=���=b<�=�A�=��=��=\M�=�$�=J��=ȕ�=���=��=��=���=���=�B�=\b�=��=h�=��=���=���=
��=���=o� >]U>:l>�!>~>�   �   �n>�6>��>T>��>�G>��>	�>�N>uF>i>��>�>1�>�5>Z�>�J>/�>��>��>->��>�>�1>��=�)�=6�=؀�=X��=��=�{�=��=j��=vg�=�0�=4�=��=�C�=gL�= ��=h��=���=��=�t�=�p�=�C�=n��=���=6�=i� >W>jf><>�h>�   �   [>��>]R>}�>�(>��>�>Ⱥ >.� >{z >� >�� >Rc>9�>�>�4>��>�B>��>!�>1S>
�>��>^F>���=��=���=ZK�=���=$��=6��=:�=.A�=��=%��=!
�=Fi�=��=!�=@D�=Xn�=�`�=���=P��=�t�=Z�=Bn�=(A�=Vx�=<� >i[>pT>J�>(>�   �   o�>\>e�>m�>�>�v >���=���=`w�=�^�=|��=^�==1 >�� >݉>�E>��>�>n�> +>�	><�>Ӭ>�e>,t�=�e�=���="��="�=�l�=���= ��=X��=:��=���=&��=�g�=��="�=`�=�	�=��=��=���=R�= |�=,��=B�=��=�$>�_>�4>�>��>�   �   :�>g.>j>� >Lv�=4��=Ɠ�=z��=��=���=d:�=��=�*�=���=% >�>+�>�>�9>U�>	�>�U>ɤ>G�>� >�h�=t�=PF�=�!�=(��=:��=J��=L,�=�q�=��=���=�a�=N
�=��=ڻ�=$��=D��=.��=��=�D�=�N�=6�=f7�= ��=�V>�a>>�G>�/>�   �   ��>+>  >2�=��=�6�=���=~�=���=ĥ�=��=���=z>�=f��=,��=~��=�� >�x>�F>��>W >�>p�>��>�q >���=��=�U�=Ҟ�=���=>��=DW�=�:�=���="6�=:��=j%�=���=�y�=b&�=���=���=�T�=B�=t��=��=���=`��=sY >�>�^>��>z�>X|>�   �   �� >fu�=d�=N��=j/�=P �=�+�=���=T��=���=X6�=�8�=��=���=���=�m�=���=M! >F+><�>r�>?�>"}>��>�� >6��=���=���=�m�=��= ��=��= ��=ا�=�Q�=\��=�w�=�=��=@�=rG�=�
�=�/�=&��=x��=���=���=j�=�� ><�>�T>�z>->>ک>�   �   R:�=Ƒ�=ڰ�=x��=���=e�=�C�=F��=ܹ�=By�=���=x�=���=��=Գ�=Č�=�w�=pL�=���=L>t�>�H>~[>Z>�L>�1 >��=b(�=�o�=���=��=���=���=T��=
��=�z�=��=��=��=P�=�0�=���=nH�=�#�=���=Ȗ�=���=K >QU>E�>�B>�>��>*� >�   �   ���=N��=�#�=P��=�y�=���=B�=�B�=b(�=���=�[�=���=ԟ�=N/�=�.�=ft�=N��=~)�=�C�=���=>��>+1>�(>��>�� >6��=$��=���=�#�=���=�y�=���=��=C�=�(�=��=\�=��=(��=�/�=�.�=�t�=���=�)�=�C�=���=*>��>+1>�(>��>�� >��=�   �   4(�=�o�=~��=���=���=���=���=���=rz�=Z�=���=��=�O�=�0�=D��=*H�=�#�=���=���=\��=	K >IU>B�>�B>�>Ú><� >�:�=���=��=���=.��=^e�=>D�=���=:��=�y�=��=��=���=
�=��=
��=(x�=�L�=���=\>��>�H>~[>Z>�L>�1 >ȇ�=�   �   f��=rm�=��=��=Ȁ�=���=���=JQ�= ��=Dw�=��=���=��=&G�=�
�=b/�=��=L��=j��=l��=R�=~� >7�>�T>�z>7>>�>�� >�u�=��=���=�/�=� �=(,�=���=���=���=�6�=�8�=f��=���=���=n�=��=d! >\+>K�>~�>G�>&}>��>�� >��=ڏ�=�   �   �U�=���=n��= ��=�V�=P:�=>��=�5�=��=%�=���=Ly�=&�=<��=H��=�T�=�=L��=��=���=L��=kY >�>�^>��>��>f|>��>?>6 >f�=�=&7�=Ч�=X~�= ��=��=>�=��=�>�=���=h��=���=ȃ >�x>�F>��>d >�>p�>��>�q >���=з�=�   �   *F�=�!�=���=��=��=
,�=�q�=Ҥ�=���=�a�=
�=���=���=��=��=���=��=�D�=bN�=�=T7�=���=�V>�a>!>�G>�/>I�>x.>0j>,� >~v�=t��=��=���=��=���=�:�=��=�*�=ޠ�=7% >�>C�>�>�9>_�>�>�U>Ȥ>C�>� >�h�=\�=�   �   ��= �=xl�=|��=��=$��=��=���=���=�g�=L�=� �=/�=�	�=���=��=h��=>�=�{�=��=.�=��=�$>�_>�4>�>��>{�>j>r�>��>�>�v >���= ��=�w�=�^�=���=D^�=T1 >�� >�>	F>��>+�>v�>+>�	>?�>լ>�e> t�=�e�=���=�   �   BK�=���=��=��=�9�=A�=��=���= 
�=i�=��=��=D�=4n�=�`�=���=@��=�t�=J�=8n�="A�=Rx�=:� >l[>qT>O�>�(>b>��>fR>��>�(>��>>׺ >?� >�z >� >�� >`c>H�>�>�4>��>�B>��>(�>6S>�>��>ZF>���=���=p��=�   �   Ȁ�=L��=��=�{�=���=U��=]g�=d0�=�3�=ڌ�=�C�=XL�=��=X��=���=؅�=�t�=�p�=�C�=h��=���=4�=j� >W>kf>@>�h> o>�6>��>T>��>H>��>�>�N>�F>i>��>�>:�>�5>a�>�J>4�>��>��>2>��>�>�1>ܡ�=�)�=.�=�   �   Z<�=�A�=��=��=TM�=�$�=E��=ƕ�=~��=��=��=���=���=�B�=\b�=��=n�=��=���=���=��=���=q� >_U>:l>�!>~>M�>�[>��>��>�>׃>r>h�>��>�>�>��>	_>��>�l>��>hv>4�>�>��>֍>��>��>�*>2��=� �=���=�   �   ؀�=\��=��=|�=��=v��=~g�=�0�=4�=��=�C�=�L�=7��=w��=���=���=�t�=�p�=�C�=v��=���=<�=n� >"W>nf>A>�h>�n>�6>��>T>��>H>��>�>�N>}F>i>��>�>6�>�5>`�>�J>1�>��>��>4>��>�>�1>��=�)�=:�=�   �   bK�=���=,��=H��=&:�=@A�=��=3��=?
�=bi�=��=F�=VD�=rn�=�`�=���=n��=�t�=l�=Tn�=8A�=`x�=A� >q[>tT>N�>�(>c>��>dR>��>�(>��>>Ѻ >;� >�z > � >�� >\c>D�>�>�4>��>�B>��>(�>:S>�>��>bF>���=��=���=�   �   4��=8�=�l�=���=<��=v��=]��=���=J��=�g�=��=V�=��=�	�=D��=��=���=p�=|�=>��=T�=��=%>�_>�4>�>��>|�>i>o�>|�>�>�v >���=��=�w�=�^�=���=8^�=M1 >�� >�>F>��>+�>w�>+>�	>E�>ڬ>�e>4t�=f�=���=�   �   fF�="�=B��=X��=n��=t,�=(r�=F��=*��=/b�=�
�=P��=
��=T��=r��=\��=�=�D�=�N�=P�=�7�=��= W>�a>&>�G>�/>J�>t.>*j>(� >vv�=f��=��=���=��=���=�:�=��=�*�=Р�=2% >�>>�>�>�9>`�>�>�U>Ф>P�>� >�h�=��=�   �   �U�=���=ƿ�=h��=pW�=�:�=���=T6�=r��=�%�=,��=�y�=�&�=���=���=�T�=t�=���=��=���=���=Y >��>�^>��>��>i|>��>=>1 >Z�=��=7�=���=D~�=���=���=.�=���=�>�=���=X��=���=ă >�x>�F>��>g >�>{�>��>�q >��=��=�   �   ���=�m�=�=R��=J��=T��=��=�Q�=���=�w�=T�=T��=��=�G�=:�=�/�=X��=���=���=���=��=�� >H�>�T>�z>=>>�>�� >�u�=��=���=�/�=� �=,�=���=���=���=�6�=�8�=R��=��=���=�m�=���=_! >W+>J�>��>N�>.}>��>�� >R��=��=�   �   �(�=p�=��=��=*��=2��=���=N��={�=�=4��=(�=DP�=.1�=̒�=�H�=$�=��=��=���='K >]U>Q�>�B>�>Ț>?� >~:�=��=��=���=��=He�=&D�=���= ��=�y�=���=��=���=��=��=���=x�=�L�=���=]>��>�H>�[>i>�L>2 >��=�   �   F��=���=$�=Ȼ�=$z�=(��=��=^C�=)�=P��=L\�=N��=l��=�/�=/�=�t�=���=�)�=D�=���=9>��>;1>�(>��>�� >:��=��=t��=�#�=���=�y�=؊�=��=C�=�(�=���=�[�=��=��=�/�=�.�=�t�=|��=�)�=�C�=���=+>��>71>�(>��>�� >X��=�   �   �:�="��=>��=���=d��=�e�=zD�=ܭ�=x��=�y�=B��=�=��=D�=X��=@��=\x�=�L�=���=n>��>�H>�[>e>�L>�1 >��=\(�=�o�=���=ҥ�=���=���=<��=��=�z�=��=Щ�=��=�O�=�0�=~��=bH�=�#�=���=���=|��=K >UU>N�>�B>�>њ>L� >�   �   � >�u�=��=���=�/�=� �=b,�=6��=���=��=�6�=<9�=���=*��=���=>n�=0��=w! >n+>[�>��>S�>1}>��>�� >>��=���=���=�m�=��=��= ��=��=���=�Q�=B��=�w�=��=���=*�=ZG�=�
�=�/�=��=p��=���=���=p�=�� >G�>�T>�z>C>>��>�   �   ��>P>H >��=:�=T7�=��=�~�=8��=H��=v�=D��=�>�=���=���=���=߃ >�x>�F>��>n >�>|�>��>�q >���=��=�U�=Ȟ�=���=0��=8W�=�:�=v��=
6�=$��=T%�=���=�y�=L&�=j��=v��=�T�=8�=n��=��=���=d��=vY >�>�^>��>��>u|>�   �   W�>�.>Aj>>� >�v�=���=0��=��=�=���=�:�=�=+�=��=L% >�>R�>��>�9>m�>�>�U>Ӥ>K�>� >�h�=t�=JF�=�!�=��=,��=:��=6,�=�q�=��=���=�a�=8
�= ��=���=��=4��= ��=��=�D�=~N�=4�=h7�=��=�V>�a>*>�G>�/>�   �   ��>w>��>��>�>�v >���=D��=�w�=�^�=ح�=h^�=g1 >�� > �>F>��>:�>��>+>�	>F�>۬>�e>4t�=�e�=���=��=�=�l�=���=��=H��=(��=���=��=�g�=t�=�=T�=�	�=��=��=~��=L�=�{�=(��=@�=��=%>�_>�4>�>��>�   �   k>��>oR>��>�(>ǖ>>� >M� >�z >� >�� >mc>T�>��>�4>��>�B>��>0�><S>�>��>bF>���=��=���=TK�=���=��=0��=:�= A�=��=��=
�=4i�=��=�=0D�=Fn�=�`�=���=N��=�t�=X�=@n�=(A�=Zx�=@� >n[>wT>R�>�(>�   �   o>�6>��>T>��>H>��>�>�N>�F>i>��>�>=�>�5>e�>�J>7�>��>��>5>��>�>�1>��=�)�=2�=Ԁ�=V��=��=�{�=��=h��=jg�=u0�=
4�=��=�C�=aL�=��=d��=���=ޅ�=�t�=�p�=�C�=n��=���=8�=n� >W>mf>B>�h>�   �   �I>�%>.�>(�>)>g�>u>�3>	>�>�>�F>x�>��>OM>5�>*>�J>l><`>E>��>�>^�>*Z >ns�=:��=��=�t�=~"�=���=D��=d�=|t�=fA�=R��=�t�=���=hT�=���=}�=��=b��=�'�=�o�=���=���=�T�=�G >d�>��>P}>c�>�@>�   �   �4>�>�>Kf>>�>�F>�>��>��>m�>�>�a>;>�%>֌>u�>�0>~W>Q>r>��>(�>F�>d >H��=��=���=��=�f�=�3�=NC�=���=��=���=�Q�=��=�\�=��=���=���=R[�=�D�=�n�=��=���=,��=�t�=aR >է>�>�x>��>C1>�   �   ��>{�>�f>��>�>�><�>u>zH>�<>�R>ֈ>/�>�?>O�>�$>��>��>e>�#>��>�>	�>��>*� >D��=l]�=>y�=�^�=�1�=b�=B�=���=���=��=*��=�!�=��=���=j�=���=ra�=�2�=�A�=�d�=�t�=�O�=���=r >�>�>zj>��>o>�   �   K�>4@>;�>-Q>�>�M>�� >� >�[ >�M >�f >(� >�� >*r>��>H{>��>�g>ҵ>��>��>j>��>y�>� >�v�=�=Nf�=�y�=�y�=6��=���=.��=H��=���=J��=�'�=���=���=� �=&��=�=T��=P��=���=Hm�=��=i�=i� >��>��>�Q>#�>�>�   �   >��>�>j>�� >�6 >Xo�=.��=�:�=��=$R�=f��=��=j] >� >��>�2>��>�+>in>z>HD>��>r�>�� >@3�=H�=���=���=n1�= �=.�=���=V�=�h�=�:�=H��=�M�= ��=���=B �=Z;�=���=D\�= �=���=� �=*0�=~� >�>�>u->^>rM>�   �   ,Y>��>�>�N >� �=���=��=V��=�2�=J�= L�=���=��=t�=^|�=�} >�;>d�>*>��>L> >ӽ>�>�6>�
 >�I�=�#�=f��=�F�=���=z��=���=8V�=̋�=0t�=x�=P��=p��=̎�=���=���=��=J��=.��=F�=F_�= >q4>h>.�>2�>�>,�>�   �   ��>Y� >���=�=JN�=4��=[�=�W�=*��=��=���=��=���=�
�=���=�q�=n >\� >��>YM>l�>��>;�>�?>�>։ >���=6��=��=���=T��=̏�=��=ʹ�=��=��=��=�/�=&E�=���=(8�=&��=|��=���=L�=n�=���=l� >��>�;>��>{�>��>�->�   �   U� > z�=f�=�E�=r8�=r]�=���=��=T��=���=��=��=l�=
��=��=h��=\��=v��=�� >"�>�3>Q�>C�>~_>��>�>�
 >Ъ�=,��=Z/�=�a�=b��=`X�=*]�=l��=���=ķ�=b�=j�=���=���=��=��= ��=hE�= ��=�  >:>��>A_>��>i{>X>��>�   �   ���=�?�=T��=W�=$��=6��=^�=���=���=���=X�=���=�c�=�5�=�Z�=���=�'�=:��=Z��=� >��>�8>=>|{>Z->H�>�� >���=�?�=���=<W�=`��=r��=��=.��=���=���=��="��=&d�=�5�=�Z�=4��=�'�=b��=z��=!� >�>�8>=>|{>U->@�>�� >�   �   ���=��=,/�=fa�=*��= X�=�\�=*��=b��=|��= �=,�=t��=���=t�=���=���=FE�=���=�  >0>��>?_>��>n{>a>ŀ>f� >Dz�=>f�=�E�=�8�=�]�=���=R��=���=��=8�=@��=��=J��=D��=���=���=���=�� >,�>�3>X�>D�>�_>��>�>�
 >�   �   ��=���=���=(��=���=���=���=��=��=���=l/�=�D�=R��=�7�=���=L��=���=,�=N�=���=c� >��>�;>��>~�>��>�->�>j� >��=D�=|N�=h��=<[�= X�=h��=2��=0��=X��=֢�=$�=ƭ�=�q�=� >o� >��>dM>w�>��>>�>�?>�>Ή >���=�   �   �#�=J��=�F�=X��=B��=���= V�=���=�s�=<�=��=>��=���=b��=���=��=$��=��=F�=,_�=� >k4>f>/�>3�>�>7�>9Y>��>>�N > !�=���= ��=���=&3�=~�=XL�=���=6��=��=�|�=�} >�;>r�>9>��>U>>Խ>�>�6>�
 >�I�=�   �   ���=���=J1�=�~�=�=���=�U�=�h�=�:�=��=pM�=ҋ�=b��= �=2;�=Ա�=$\�=��=޷�=� �=0�=y� >
�>�>y->^>|M>>��>�> j>� >�6 >�o�=X��=�:�=��=VR�=���=J��=�] >/� >̖>�2>�>�+>rn>z>LD>��>p�>�� >.3�=<�=�   �   :f�=fy�=�y�=��=���=��=$��=���= ��=�'�=���=���=� �=��=��=2��=8��=|��=8m�=v�=i�=d� >��>��>�Q>&�>�>V�>B@>G�>;Q>�>�M>� >$� >�[ >
N >�f >:� >�� >:r>��>X{>��>�g>ٵ>��>��>j>��>z�>� >�v�=�=�   �   ,y�=�^�=�1�=N�=�A�=h��=���=���=��=�!�=Λ�=���=R�=���=Xa�=�2�=�A�=�d�=�t�=�O�=���=r >�>�>yj>��>t>��>��>�f>��>%�>�>F�>$u>�H>�<>�R>�>;�>�?>Z�>�$>��>��>j>�#>��>�>	�>��>%� >:��=b]�=�   �   ���=���=�f�=�3�=<C�=���=��=���=�Q�=���=�\�=ܽ�=���=���=H[�=�D�=�n�=��=���="��=�t�=_R >֧>�>�x>��>G1>�4>�>�>Mf>>��>�F>�>��>��>u�>�>�a>Ծ>�%>܌>x�>�0>�W>!Q>v>��>&�>E�>�c >D��=��=�   �   ��=�t�=x"�=���=@��=d�=vt�=dA�=N��=�t�=���=jT�=���=}�=��=`��=�'�=�o�=���=���=�T�=�G >c�>��>L}>c�>�@>�I>�%>/�>)�>)>g�> u>�3>	>�>�>�F>u�>��>LM>6�>,>�J>
l>;`>F>��>�>_�>$Z >js�=8��=�   �   ���=��=�f�=�3�=RC�=���="��=ĩ�=�Q�=��=�\�=���=
��=���=\[�=�D�=�n�=��=���=,��=�t�=cR >ۧ>�>�x>��>I1>�4>�>�>Mf>>��>�F>�>��>��>t�>�>�a>Ѿ>�%>݌>v�>�0>�W>Q>s>��>'�>G�>d >J��=��=�   �   @y�=�^�=�1�=p�=$B�=���=���=$��=<��="�= ��=���=|�=���=�a�=�2�=
B�=�d�=u�=�O�=���=r >�>	�>}j>��>v>��>��>�f>��>!�>�>E�>!u>�H>�<>�R>�>8�>�?>W�>�$>��>��>j>�#>��>�>�>��>+� >J��=v]�=�   �   Zf�=�y�=�y�=L��=���=J��=`��=���=`��=(�=ܞ�=���=� �=@��=�=f��=j��=���=Zm�=��= i�=p� >��>��>�Q>'�>�>U�>=@>F�>9Q>�>�M>� >� >�[ >N >�f >6� >�� >4r>��>T{>��>�g>ٵ>��>��>$j>��>��>� >�v�=(�=�   �   ���=���=�1�=�=H�=���=.V�=�h�=�:�=l��=�M�=(��=���=^ �=z;�=��=^\�=�=��=� �=>0�=�� >�>��>|->^>|M>>��>�>j>� >�6 >to�=P��=�:�=��=FR�=���=<��=z] >)� >ɖ>�2>�>�+>sn>z>PD>��>w�>�� >L3�=\�=�   �   �#�=���=�F�=���=���=޻�=\V�=��=Tt�=��=z��=���=��=���=���=��=j��=J��=:F�=X_�= >x4>r>7�>7�>�>6�>9Y>��>�>�N >!�=���=��=z��=3�=l�=LL�=���=&��=��=~|�=�} >�;>q�>6>��>Y>
>۽>�>�6>�
 >J�=�   �   P��=.��=Σ�=x��=��=B��=���=�=�=>��=�/�=TE�=���=L8�=L��=���=���=l�=��=���=w� >��>�;>
�>��>��>�->�>e� >��=@�=tN�=\��=&[�=
X�=T��=��= ��=H��=¢�=�=���=�q�= >l� >��>dM>z�>��>F�>@>�>�� >���=�   �   ��=H��=r/�=�a�=���=�X�=T]�=���=���=��=��=��=ޣ�=��=��=��=D��=�E�=��=�  >E>��>L_>��>q{>d>ǀ>c� ><z�=,f�=�E�=�8�=�]�=���=<��=���=Ҿ�="�=0��=��=8��=<��=���=~��=���=�� >-�>�3>_�>M�>�_>��>�>�
 >�   �   ڊ�=@�=���=`W�=���=���=��=X��=��=��=��=R��=Vd�=6�="[�=X��=�'�=���=���=/� >�>�8>H>�{>]->L�>�� >���=�?�=p��=.W�=P��=b��=��=��=���=���=��=��=d�=�5�=�Z�=&��=�'�=X��=z��=!� >�>�8>E>�{>b->T�>�� >�   �   r� >`z�=Vf�=�E�=�8�=�]�=��=|��=���=��=d�=r��=��=n��=p��=ħ�=���=���=�� >;�>�3>`�>N�>�_>��>�>�
 >Ȫ�= ��=J/�=�a�=V��=JX�=]�=V��=���=���=L�=X�=���=���=��=��=��=`E�=���=�  >;>��>K_>��>u{>k>р>�   �   �>y� >8��=d�=�N�=���=d[�=HX�=���=\��=\��=���=���=H�=��=�q�=� >{� >��>oM>��>��>F�> @>
�>׉ >���=2��=��=���=L��=���=��=���=��=��=���=�/�=E�=x��=8�=��=r��=���=F�=h�=���=m� >��>�;>	�>��>��>�->�   �   DY>��>>�N >@!�=��=B��=���=L3�=��=~L�=��=V��=��=�|�=�} >�;>�>D>��>\>>۽>�>�6>�
 >�I�=�#�=^��=�F�=x��=j��=���=&V�=���=&t�=b�=<��=^��=���=���=���=��=@��=&��=F�=B_�= >t4>n>8�>9�>�>A�>�   �   $>Ĕ>	>0j>� >�6 >�o�=���=;�=�=tR�=���=h��=�] >?� >ؖ>�2>�>�+>xn> z>SD>��>t�>�� >@3�=J�=���=���=d1�=�~�="�=���= V�=�h�=�:�=2��=�M�=��=x��=0 �=N;�=���=<\�=��=���=� �=20�=�� >�>��>�-> ^>�M>�   �   Z�>J@>P�>EQ>)�>N>� >3� >�[ >N >�f >H� >�� >Dr>��>`{>
�>�g>ߵ>��>��>"j>��>|�>� >�v�=�=Ff�=vy�=�y�=.��=���=&��=8��=���=@��=�'�=���=���=� �=��=��=H��=J��=���=Dm�=��=i�=l� >��>��>�Q>+�>"�>�   �   ��>��>�f>��>/�>�>P�>.u>�H>�<>�R>�>C�>�?>b�>�$>��>��>q>�#>��>�>�>��>+� >F��=p]�=6y�=�^�=�1�=\�=B�=z��=���=��=$��=�!�=��=���=`�=���=la�=�2�=�A�=�d�=�t�=�O�=���=r >�>�>j>��>{>�   �   �4>�>�>Rf>>��>�F>�>��>��>y�>�>�a>վ>�%>ߌ>y�>�0>�W>"Q>v>��>)�>F�>d >J��=��=���= ��=�f�=�3�=FC�=���=��=���=�Q�= ��=�\�=��=���=���=N[�=�D�=�n�=��=���=(��=�t�=bR >٧>�>�x>��>K1>�   �   9>��>η>�u>Y+>+�>ĝ>Eg>OB>�1>�7>�R>C>��>v�>>>>=z>��>@�>��>R�>33>(�>��>8� >��=��=�,�=p+�=H�=�%�=nb�=P��=���=�e�=tv�=�'�=*}�=@r�=��=z�=.{�=>B�=�?�=�S�=\^�=�D�=<��=}!>">$�>�r>�>�>�   �   :�>��>�>b\>E>��>}>E>[>�>>�0>c_>�>~�>S&>�e>��>��>��>��>�/>f�>r�>�� >&��=b%�=�Q�=�V�=P�=6]�=D��=�1�=�.�=���=D��=jr�=F��=���=�@�=rG�=^��=z�=�q�=�~�=���=pa�=* >J(>>��>�n>�>��>�   �   q�>y�>�`>�> �>�g>�>��>p�>��>�>��>3>&D>��>_�>n(>�c>�>4�>�q>0&>
�>��>�>���=b|�=l��=���=���=�=S�=���=���=F��=���=�N�=P��=���=F�=�	�=Bm�=n�=�=^��=���=2��=i  >f<>�'>v�>�a>j�>u�>�   �   v~>�E>~�>�>B4>��>*�>�=>�>�� >z	>c->Uh>n�>@>$k>��>/>>E>�]>�O>�>��>�	>
6>P2 >	�=l�=6��=r��=B�=�v�=�+�=�E�=���=���=.��=(�=$��=RZ�=D�=���=�*�=��=���=R��=d>�=TR >!\>�5>E�>�K>�>��>�   �   �>#�>�c>��>x|>�>�� >�a >�0 >� >G* >�T >�� >c� >K]>��>�9>�>��>�>� >
�>�>� >�d>�x >��=<V�=f��=x�=�s�=���=4��=�=@��=���=F��=R��=.��=V�=���=X�=|��="0�=j��=f|�=���=� >��>�F>q�>�,><R>I>�   �   ƙ>�.>]�>$%>�� >C >�S�=B��=�:�=2�=l1�=
��=�8�=� >#� >�>a�>�	>r>½>��>��>��>�;>��>z� >���=�q�=��=��=B&�=���=���=�=���=p�=Z��=��=���=0�=���=���=>�=��=�&�=���=t��=q� >�>�Y>��>�>�>��>�   �   >|>�� >]9 >�,�=���= �=�<�=@��=���=��=2�=���=���=��=�% >]� >�`>u�>�T>a�>W�>��>�X>��>�,> T >"��=���=�M�=|�=���=l�=p��=2V�=X��=�b�=T��=c�=,��=�&�=
�=<$�=�\�=P��=��=�] >U9>0�>)m>&�>�>;�>�r>�   �   sb>ն >t��=m�=���=P��=�t�=*��=t�=b��=*�=,��=�n�=���=���=6W�=���=�� >0O>q�>RJ>��>V�>Du>>�>�� >� >�&�=�'�=�'�=�?�=���=b�=��=�_�=x(�=�d�=��=�&�=$��=�I�=:.�=<+�=�'�=� >�� >�> ">>��>��>#]>5�>�   �   � >��=|�=�L�=
��=�=`��=���=B9�=.�=z;�="��=8��=�=v��=xF�=��=*��=� >�_>[�>/X>9�>�>S]>�>i> � >$��=��=�L�=2��=4�=���=���=t9�=^�=�;�=R��=b��=D�=���=�F�=�=D��=�� >�_>b�>5X>:�>�>O]>�>i>�   �   � >�&�=�'�=l'�=�?�=^��=4�=x�=�_�=F(�=�d�=��=�&�=���=�I�=.�=+�=f'�=� >�� >��>">�~>��>��>']><�>�b>� >���=6m�= ��=v��=�t�=Z��=��=���=X�=Z��=o�=Ǝ�=���=ZW�=���=�� ><O>z�>YJ>��>W�>Bu>>�>�� >�   �   
��=���=�M�=^�=���=H�=B��=V�=,��=�b�=*��=�b�=��=�&�=�	�=$�=�\�=:��=���=�] >M9>)�>%m>'�>�>@�>�r>>%|>� >o9 >�,�= �=< �=�<�=l��=Е�=@��=@2�=���=��=��=�% >j� >a>�>�T>e�>^�>��>�X>��>�,>�S >�   �   �q�=l�=��=$&�=���=���=��=~��=B�=2��=z�=���=�/�=���=���=�=�=���=�&�=n��=^��=l� >�>�Y>��>�>�>��>Й>�.>h�>3%>�� >U >T�=f��=�:�=\�=�1�=2��=�8�=� >3� >�>p�>�	>!r>ͽ>��>��>�>�;>��>t� >��=�   �   *V�=L��=^�=~s�=���=��=� �=��=���="��=4��=��=4�=���=<�=^��=0�=X��=T|�=���=� >}�>�F>q�>�,>BR>I>�>.�>�c>��>�|>�>� >�a >�0 >� >Y* >�T >� >v� >X]>��>�9>�>��>�>� >�>�>� >�d>�x >��=�   �   l�=(��=\��=.�=lv�=�+�=rE�=���=���=��=�=��=:Z�=�C�=t��=�*�=���=���=D��=T>�=QR >\>�5>F�>�K>�>��>�~>�E>��>��>N4>��>6�>�=>�>�� >�	>q->ah>}�>K>0k>��>6>FE>�]>�O>�>��>�	>6>M2 >	�=�   �   ^��=���=v��=��=�R�=���=���=(��=���=�N�=:��=���=2�=�	�=4m�=`�=�=R��=���=(��=f  >c<>�'>u�>�a>l�>u�>s�>~�>�`>�>�>�g>�>��>x�>��>�>��>;>/D>��>h�>t(>�c>�>8�>�q>3&>�>��>�>���=\|�=�   �   zQ�=�V�=
P�=,]�=8��=�1�=�.�=z��=:��=^r�=@��=���=�@�=lG�=T��=z�=�q�=�~�=|��=la�=' >H(>>��>�n>�>��><�>��>�>g\>G>��>}>"E>^>�>>�0>d_>�>~�>X&>�e>��>��>��>��>�/>h�>r�>�� > ��=d%�=�   �   �,�=n+�=D�=�%�=jb�=V��=���=�e�=nv�=�'�=0}�=Dr�=��=x�=.{�=<B�=�?�=�S�=Z^�=�D�=>��=}!>!>%�>�r>�>�>;>��>ͷ>�u>Y+>-�>>Eg>QB>�1>�7>�R>B>��>t�>?>><z>��>A�>��>R�>63>,�>��>6� >��=��=�   �   �Q�=�V�=P�=<]�=D��=�1�=�.�=���=F��=rr�=N��=���=�@�=xG�=f��=z�=�q�=�~�=���=ta�=+ >L(>!>��>�n>�>��><�>��>�>g\>D>��>}>#E>^>�>>�0>__>�>��>V&>�e>��>��>��>��>�/>h�>u�>�� >"��=h%�=�   �   p��=���=���=�=S�=���=���=H��=���=�N�=\��=���=J�=
�=Nm�=x�=$�=f��=��=6��=n  >h<>�'>x�>�a>k�>x�>v�>�>�`>�>�>�g>�>��>w�>��>�>��>9>.D>��>i�>q(>�c>�>7�>�q>1&>�>��>�>���=j|�=�   �   "l�=F��=x��=N�=�v�=�+�=�E�=���=���=@��=6�=B��=\Z�=D�=���=�*�=��=���=`��=l>�=YR >%\>�5>I�>�K>�>��>�~>�E>��>��>I4>��>2�>�=>�>�� >�	>m->[h>x�>G>-k>��>7>EE>�]>P>�>��>�	>6>U2 >(	�=�   �   HV�=t��=��=�s�=���=H��=�=N��=���=Z��=l��=J��=l�=���=r�=���=60�=z��=t|�=���=%� >��>�F>u�>�,>BR>I>�>)�>�c>��>�|>�>� >�a >�0 >� >S* >�T >� >q� >T]>��>�9>�>��>�>� >�>��>� >�d>�x >��=�   �   �q�=��=,��=X&�=��=��=6�=���=��=v��=��=���=20�=���=���=8>�=,��='�=���=���=w� >#�>�Y>��>�>�>��>љ>�.>d�>/%>�� >O >�S�=Z��=�:�=J�=�1�=&��=�8�=� >0� >�>n�>�	>r>˽>��>��>��>�;>��>�� >
��=�   �   6��=���=�M�=��=���=��=���=LV�=t��=�b�=t��=<c�=F��=�&�= 
�=X$�=]�=f��=$��=�] >[9>5�>/m>,�>�>D�> s>>!|>� >l9 >�,�=
 �=( �=�<�=^��=�=8��=22�=���=��=��=�% >h� >a>}�>�T>h�>a�>��>�X>��>�,>T >�   �   � >�&�=(�=�'�= @�=���=|�=��=�_�=�(�=�d�=��=�&�=@��=�I�=T.�=X+�=�'�=� >�� >�>%">>��>��>)]><�>b>ݶ >���=0m�=��=l��=�t�=F��=��=���=J�=L��=�n�=���=���=TW�=���=�� >:O>{�>\J>�>^�>Ku>>��>�� >�   �   )� ><��=��=M�=P��=V�=���=���=�9�=��=�;�=v��=���=`�=���=�F�=.�=Z��=� >	`>k�><X>A�>�>V]>
�>i>� >��=��=�L�=(��=(�=|��=���=h9�=L�=�;�=B��=R��=4�=���=�F�=
�=@��=�� >�_>d�>8X>@�>�>Z]>�>i>�   �   �b>� >���=Rm�=:��=���=�t�=t��=��=���=x�=z��= o�=��=���=|W�=��=�� >EO>��>bJ>�>^�>Gu>
>��>�� >� >�&�=�'�=�'�=�?�=v��=T�=��=�_�=b(�=�d�=��=�&�=��=�I�=4.�=6+�=z'�=� >�� >�>"">>��>��>/]>F�>�   �   >.|>� >~9 >�,�=2 �=T �=�<�=���=��=^��=^2�=���=(��=��=�% >y� >a>��>�T>p�>`�>��>�X>��>�,> T > ��=���=�M�=v�=���=`�=`��="V�=L��=�b�=J��=c�=��=�&�=�	�=6$�=�\�=N��=��=�] >W9>2�>.m>.�>�>G�>s>�   �   ٙ>�.>o�>@%>�� >^ >T�=���=�:�=v�=�1�=N��=�8�=� >A� >�>x�>
>*r>ҽ>��>��>��>�;>��>z� >���=�q�=|�=��=:&�=���=���=�=���=f�=J��=��=���=0�=���=���=>�=��=�&�=���=r��=s� >!�>�Y>��>�>�>��>�   �   �>6�>�c>��>�|>�>� >�a >�0 > >c* >�T >�� >}� >d]>��>�9>��>��>�>� >�>��>� >�d>�x >��=6V�=^��=p�=�s�=���=*��=� �=2��=���=4��=L��=$��=F�=���=N�=r��=0�=d��=f|�=���=!� >��>�F>v�>�,>FR>"I>�   �   �~>�E>��>��>S4>��>?�>�=>�>�� >�	>{->hh>��>U>4k>��>:>GE>�]>P>�>��>�	>6>Q2 >	�=l�=0��=l��=8�=~v�=�+�=�E�=���=���="��=�= ��=FZ�=�C�=���=�*�=���=���=R��=`>�=VR >#\>�5>G�>�K>�>��>�   �   v�>��>�`>�>�>�g>�>��>��>��>�>��>C>7D>��>m�>u(>�c>�>:�>�q>5&>�>��>�>���=b|�=j��=���=|��= �=S�=���=���=:��=���=�N�=L��=���=<�=�	�=>m�=l�=�=X��=���=2��=l  >h<>�'>w�>�a>n�>}�>�   �   <�>��>�>j\>K>��>}>(E>a>�>>�0>i_>�>��>Z&>�e>��>��>��>��>�/>f�>r�>�� >&��=`%�=�Q�=�V�=P�=4]�=>��=�1�=�.�=���=@��=`r�=D��=���=�@�=pG�=^��=z�=�q�=�~�=���=pa�=( >K(> >��>�n>�>��>�   �   ��>:�>b�>�Y>>.�>��>�r>�K>a2>[(>�->�@>	_>��>�>I�>3�>0>.�>��>��>�O>��>u0>Gm >V�=*�=��=��=���=��=ni�=��=���=O�=��=�R�=���=��=,��=<�=�2�=�Q�=4��=���=���=9� >��>c>��>q\>��>��>�   �   Z�>��>�~>2H>}
>�>9�>�[>�3>�>>5>�+>�K>s>��>��>:�>��>��>��>�>�P>��>�6> v >�/�=�E�=�=�=\,�=T'�=�D�="��=�3�=~(�=��=�K�=��=T/�=L@�=���=>e�=FX�=�r�=V��=���=j��=c� >8�>�c>�>X>#�>��>�   �   8�>�~>zO>?>!�>�>�L>�>��>��>R�>��>��>�>�>>\o>"�>4�>��>��>��>��>�S>5�>�H>ԏ >�r�=���=J��=���=���=���=�!�=���=h��=��=���=>�=4��=���=<0�=���=���=b��=���=�
�=� >� >q�>)f>��>K>�>Q�>�   �   )c>�;>%>%�>Cp>�$>��>�>{>�a>�[>Xh>A�>M�>D�>�">d\>��>��>j�>�>��>5X>*�>\f>�� >j��=��=�7�=�G�=L`�=&��=� �=��=���=��=���=��=̯�=^��=P�=���=�x�=�q�=�x�=vx�=�. >�>��>�i>t�>�5>�d>zr>�   �   �>V�>P�>!E>��>j�>�K>�>� >� >�� >~� >� >(0>�q>�>>�C>xx>a�>9�>b�>�]>{>m�>b� >R7 >���=��=82�=�c�=X��=R,�=<��=���=^�=�(�=nY�=���=���=�"�=��=�g�=D�=�+�=.
�=�f >2>��>Km>Y�>>7>55>�   �   p�>�n>G>�>iL>>� >+� >�O >) >I >� >4 >M >� >H� >�7>��>(�>�.>rd>Q�>��>+d>�!>2�>4>k� >d��=0��=�M�=���=�=2��=�f�=4��=.��=º�=��=�n�=�N�=j|�=R��=̇�=*A�=��=<��=I� >�_>��>�p>=�>��>5�>��>�   �   �H>��>r}>>R� >�# >"��=���=H��=zR�= Y�=��=�
�=���=P5 >$� >v>�x>��>�$>�Y>Ir>j>�>>r�>�>~� >�G >��=܎�=��=���=�6�=D�=�@�=J��=ʃ�=���=$�=���=�=T�= ��=^�=���=W> >{� >ˑ>>�r>�>��>��>��>�   �   ��>Y>B� >8M >:��=���=���=��=X��=Bn�=�|�=���=�S�=6�=��=���=K} >Y� >&w>��>,>�]>�n>']>�'>$�>=Y>&� >�# >j��=���=$.�=��=���=n&�=
��=.r�=��=(��=X��=���=��=*�=؎�=>��=(� >�A>
�>\->�s>s�>2�>(q>>->�   �   	L>q� ><& >r�=��=8��=���=R�=r��=�q�=n��= ��=r��=�`�=i�=���=0��=6~ >�>��>�>�F>Wr>�z>x_>�!>G�>L>{� >G& >��=.��=X��=���=v�=���=r�=���=<��=���=�`�=0i�=���=H��=A~ >�>Ő>�>�F>Ur>�z>s_>�!>B�>�   �   � >�# >R��=z��=.�=���=���=J&�=��=r�=��=
��=<��=l��=���=*�=���=2��=!� >�A>�>Y->�s>s�>4�>+q>C->��>'Y>M� >EM >V��=̑�=ƹ�=��=~��=fn�=�|�=���=T�=X�=6��=���=V} >`� >/w>��>,>�]>�n>']>�'> �>:Y>�   �   �G >��=�=��=���=�6�=(�=�@�=*��=���=r��=�#�=���=��= T�=��=�]�=���=M> >v� >Ƒ>>�r>�>��>��>�>�H>��>z}>>`� >�# >>��=���=f��=�R�=@Y�=��=�
�=ک�=Z5 >1� >�>�x>��>�$>Z>Lr>j>�>>m�>�>x� >�   �   T��=$��=�M�=���=��=��=�f�=��=��=���=���=�n�=�N�=R|�=<��=���=A�=��=0��=@� >�_>��>�p>;�>��>7�>�>x�>�n>M>�>sL>J� >7� >�O >8 >W > >A >$M >'� >T� >�7>��>0�>�.>wd>U�>��>-d>�!>-�>}4>g� >�   �   ���=��=$2�=�c�=B��=>,�=(��=���=�]�=�(�=\Y�=���=���=�"�= ��=pg�=�C�=�+�="
�=�f >2>��>Im>Z�>!>7>95>�>Y�>Z�>(E>��>v�>�K>�>"� >+� >�� >�� >*� >60>�q>��>>�C>x>b�>>�>e�>�]>z>g�>]� >N7 >�   �   ��=�7�=�G�=<`�=��=� �=���=��=��=���=��=���=N��=>�=v��=�x�=�q�=�x�=hx�=�. >�>��>�i>t�>�5>�d>}r>/c>�;>*>+�>Kp>�$>��>�>"{>b>�[>`h>I�>W�>K�>�">k\>��>��>o�> �>��>4X>)�>Xf>�� >f��=�   �   ��=>��=���=���=���=�!�=~��=L��=��=���=0�=&��=n��=.0�=���=���=Z��=���=�
�=� >� >o�>*f>��>K>�>R�>;�>�~>}O>B>'�>#�>�L>�>��>��>X�>��>��>�>�>>co>(�>8�>��>��>��>��>�S>6�>�H>я >�r�=�   �   �E�=�=�=X,�=N'�=�D�=��=�3�=p(�=��=�K�=��=L/�=H@�=���=8e�=BX�=�r�=V��=���=b��=`� >9�>�c>�>X>$�>��>]�>��>�~>2H>
>�>:�>�[>�3>�>$>8>�+>�K>s>��>�>@�>��>��>��>�>�P>��>�6>�u >�/�=�   �   *�=��=��=���=��=ti�=��=���=O�=��=�R�=���=��=(��=<�=�2�=�Q�=6��=���=���=8� >��>c>��>o\>��>��>��>;�>a�>�Y>>.�>��>�r>�K>`2>[(>�->�@>_>��>�>F�>6�>0>/�>��>��>�O>��>q0>Hm >V�=�   �   �E�=�=�=Z,�=V'�=�D�=,��=�3�=t(�=��=�K�=���=Z/�=L@�=���=De�=JX�=�r�=^��=���=h��=a� >:�>�c>�>X>$�>��>_�>��>�~>5H>|
>�>:�>�[>�3>�>$>6>�+>�K>!s>��>�>=�>��>��>��>�>�P>��>�6>�u >�/�=�   �   ���=N��=���=���=���=�!�=���=f��=��=���=J�=B��=���=@0�=���=���=n��=���=�
�=� >�� >q�>*f>��>
K>�>R�><�>�~>|O>@>&�> �>�L>�>��>��>V�>��>��>�>�>>ao>&�>;�>��>��>��>��>�S>7�>�H>ԏ >�r�=�   �   ��=�7�=�G�=R`�=0��=� �=��=��=��=���=��=ޯ�=j��=X�=���=y�=�q�=�x�=zx�=�. >�>��>�i>w�>�5>�d>}r>/c>�;>'>,�>Hp>�$>��>�> {>b>�[>^h>F�>S�>I�>�">l\>��>��>m�>!�>��>8X>-�>\f>�� >t��=�   �   ���=��=B2�=�c�=b��=b,�=J��=���=^�=�(�=~Y�=���=���=�"�=(��=�g�=D�=�+�=:
�=�f >2>��>Om>^�>">7>;5>�>Z�>S�>'E>��>r�>�K>�> � >&� >�� >�� >%� >00>�q>��>>�C>~x>d�>A�>h�>�]>~>m�>f� >W7 >�   �   n��=B��=�M�=���=�=H��=�f�=@��=>��=Ժ�=��=�n�=�N�=x|�=h��=އ�=>A�=��=J��=L� >�_>��>�p>?�>��>8�>�>v�>�n>K>�>qL>G� >4� >�O >3 >P >� >= > M >"� >R� >�7>��>3�>�.>xd>X�>��>2d>�!>5�>�4>p� >�   �   �G >��=��=��=Ҋ�=�6�=Z�=�@�=\��=ރ�=���=0$�=���= �=,T�=2��=^�=���=\> >�� >ё>>�r> �>��>��>�>�H>��>z}>>_� >�# >2��=���=^��=�R�=:Y�=��=�
�=ҩ�=X5 >/� >>�x>��>�$>Z>Qr>j>�>>v�>�>�� >�   �   ,� >�# >t��=���=6.�=$��=���=�&�= ��=Fr�=��=B��=j��=���=&��=2*�=��=N��=/� >�A>�>`->�s>w�>6�>.q>E->��>%Y>G� >CM >R��=���=���=��=r��=Xn�=�|�=���=T�=P�=.��=���=U} >a� >-w>��>,>�]>o>-]>�'>+�>DY>�   �   L>�� >P& >��=B��=n��=���=��=���="r�=���=Z��=���=a�=Hi�=���=^��=H~ >�>ː>�>�F>Zr>�z>x_>�!>I�>L>x� >C& >��=(��=L��=���=j�=���=�q�=���=6��=���=�`�=&i�=���=D��=>~ >�>Đ>�>�F>[r>�z>y_>�!>N�>�   �   ��>/Y>R� >PM >n��=���=޹�=��=���=zn�=}�=���=&T�=d�=L��=��=a} >e� >7w>��>,>�]>o>*]>�'>&�>?Y>#� >�# >`��=���=.�=��=���=b&�=��=r�=���=��=P��=���=��=*�=֎�=>��=(� >�A>�>`->�s>x�>7�>2q>I->�   �   �H>��>�}>%>j� >�# >T��=���=~��=�R�=VY�=(��=�
�=��=d5 >9� >�>�x>��>�$>Z>Or>j>�>>t�>�>~� >�G >��=Ԏ�=��=���=�6�=:�=�@�=B��=���=���=$�=���=�=T�=��=�]�=���=S> >{� >ϑ>	>�r>!�>��>��>�>�   �   }�>�n>S> �>|L>Q� >@� >�O >A >a >	 >L >+M >/� >_� >�7>��>7�>�.>|d>Y�>��>/d>�!>1�>�4>l� >b��=0��=�M�=���=�=,��=�f�=(��=(��=���= ��=�n�=�N�=`|�=P��=ȇ�=(A�=��=<��=I� >�_>��>�p>A�>��><�>�>�   �   �>_�>]�>/E>��>{�>�K>�>*� >4� >�� >�� >0� >80>r>��>>�C>�x>h�>C�>i�>�]>}>k�>b� >S7 >���=��=22�=�c�=P��=J,�=2��=���=�]�=�(�=hY�=���=���=�"�=��=�g�=D�=�+�=,
�=�f >2>��>Qm>]�>">7>?5>�   �   4c>�;>.>1�>Np>�$>��>��>({>b>�[>eh>O�>[�>T�>�">q\>��>��>o�>"�>��>7X>+�>\f>�� >l��=��=�7�=�G�=H`�=��=� �=��=��=��=���=��=ȯ�=X��=H�=���=�x�=�q�=�x�=rx�=�. >�>��>�i>u�>�5>�d>~r>�   �   >�>�~>�O>F>+�>$�>�L>�>��>��>[�>��>�>�>�>>ao>*�>=�>��>��>��>��>�S>9�>�H>ԏ >�r�=��=F��=���=���=���=�!�=���=`��=��=���=:�=4��=x��=:0�=���=���=`��=���=�
�=� >�� >r�>.f>��>K>��>U�>�   �   _�>��>�~>5H>�
>�><�>�[>�3>�>%>:>�+>�K>!s>��>��><�>��>��>��>�>�P>��>�6>�u >�/�=�E�=�=�=Z,�=P'�=�D�= ��=�3�=t(�=��=�K�=��=N/�=J@�=���=@e�=DX�=�r�=X��=���=j��=c� >:�>�c>�>
X>&�>��>�   �   u�>��>)n>B>�>4�>��>hg>z8>2>��>��>��>��>��>��>!>�">�,>?,>{>��>1�>Ā>� >�� >r >d
�=<��=`m�=x�=��=���=���=(+�=���=V��=��=�.�=���=N��=��=t�=���=�u�=���=�� >�j>W>��>7�>E>�z>.�>�   �   �>��>0b>5>��>f�>S�>�W>�(>�>��>��>��>��>��>�>
>)>�'>)>2>@�>��>ބ>[&>�� >�( >  �=���=���=�<�=��=��= �=8N�=���=��=���=�N�=��=B�=�0�=v��=� �=���= >�� >m>�>^�>�>X@>Pt>G�>�   �   dw>+c>�>>N>�>��>�_>)>��>t�>1�>�>��>"�>'�>��>C�>	>�> >�>��>W�>ڐ>}7>�� >D >`�=�!�=��=ړ�=�`�=�L�=ze�=���=�F�=��=dA�=H��=�a�=�S�=\{�=v��=�9�=@��= >u� >�s>J>t�>�>Q2>ua>�w>�   �   &J>U/>�>��>�>R>�>v�>�>��>tp>�e>h>v>��>;�>l�>�>�>�>�>Y>W�>=�>BS>�� >!p >t��=��=�Z�=!�=D��=
��=~	�=�\�=���=���=��=�H�=���=���=���=�7�=8��=���=4 >�� >
>v
>>M�>]>�B>�Q>�   �   �>�>B�>�x>=5>R�>��>.t>D>� >�>�>R>
$>\D>�k>j�>�>��>��>=
>q>��>�>Xx>>� >�( >�3�=��=���=���=��=���=�<�=���=b��=���=H�=ڵ�=؍�=>��=���=��=�c�=�Z >$� >��>>�u>��><�>>�>�   �   }�>m�>KU>n>��>Mw>�0>�� >�� >�� >�� >>� >\� >k� >�� >>�T>��>��>��>��>�>��>�>�>V>�� >�{ >���=���=���=F��=��=���=L�=��=��=X��=��=���=Lh�=r\�=jt�=���=^��=�� >�>��>�>Vj>��>��>��>T�>�   �   Aj>C.>�>b�>p>>�� >�� >_ >�- >i >3  >B > >�H >:� >�� >>�N>��>��>3�>+>�>��>�>E�>�A>�� >_c >���=���=&��=0��=\�=��=N�=J��=f��=F1�=���=�_�=�;�=�8�=2J�=�1 >� >r=>ʰ>h> \>Ҏ>�>��>͔>�   �   .
>��>�i>(>!� >R >D  >�x�=��=���=���=���=�#�=D��= >m\ >#� >�
>u^>��>��>>�$>c$>\>��>�>�=>�� >d >@��=���=P�=�a�=���=fc�=�-�=P.�=ne�=���=`j�=�+�=�
�=<��=�y >3� >�a>�>�>^K>jm>Ew>�h>�C>�   �   Ȥ>�K>�� >�} >g >b�=Z��=z#�=ȼ�=x��={�=ȣ�=j��=�}�=V#�=F��=YY >�� >�(>Ņ>|�>(>�8>�I>tB>|#>�>Ѥ>�K>�� >�} >s >(b�=p��=�#�=��=���=4{�=ܣ�=x��=�}�=f#�=\��=_Y >� >)>Ʌ>�>*>�8>�I>qB>x#>�>�   �   �=>�� >d >.��=r��=:�=�a�=���=Pc�=�-�=6.�=^e�=h��=Nj�=�+�=�
�=2��=�y >-� >�a>�>�>_K>jm>Hw> i>�C>6
> �>�i>/>,� >R >O  >�x�=��=���=���=���=$�=X��= >w\ >,� >�
>~^>��>��>>�$>c$>Y>��>�>�   �   �� >Xc >���=���=��=��=J�=��=6�=2��=T��=21�=��=�_�=�;�=v8�= J�=�1 >�� >p=>ư>e>\>Ԏ>�>��>Ӕ>Kj>J.>�>k�>y>>�� >�� >_ >�- >s ><  >K >  >�H >A� >�� >>�N>��>��>6�>->�>��>�>A�>�A>�   �   �{ >���=���=���=2��=���=���=�K�= ��=���=J��=��=x��=:h�=\\�=Xt�=~��=V��=�� >�>��>�>Uj>��>��>��>V�>��>r�>PU>u>��>Vw>�0>�� >�� >	� >�� >G� >g� >s� >�� >#>�T>��>��>��>��>�>��>�>�>�U>�� >�   �   �( >�3�=��=���=���=���=���=�<�=���=R��=���=:�=ε�=ʍ�=.��=���=��=�c�=�Z > � >��>>�u>��>@�>!>�>�>�>E�>�x>B5>[�>��>7t>#D>� >�>�>X>$>cD>�k>p�>�>��>��>A
>s>��>�>Tx>�> � >�   �   l��=���=�Z�=!�=4��=���=n	�=�\�=���=���=���=�H�=���=���=���=~7�=0��=���=4 >�� >>u
>>M�>`>�B>�Q>+J>Z/>�>��>�>�R>�>}�>	�>��>}p>�e>h>%v>��>A�>n�>
�>�>�>�>]>V�>>�>?S>�� >p >�   �    `�=�!�=��=֓�=�`�=�L�=pe�=���=�F�=��=\A�=<��=�a�=�S�=X{�=j��=�9�=>��= >s� >�s>J>r�>�>O2>ya>�w>kw>+c>�>>Q>�>��>�_>)> �>y�>6�>��>��>*�>$�>��>G�>		>�> >�>��>Z�>ِ>z7>�� >D >�   �   ��=���=���=�<�=��=��= �=2N�=���=
��=���=�N�=��=8�=�0�=p��=� �=���= >�� >m>�>\�>"�>Z@>St>J�>�>�>1b>5>��>l�>S�>�W>�(>�> �>��>��>��>��>	�>
>+>�'> )>7>?�>��>܄>W&>�� >�( >�   �   `
�=@��=\m�=t�=��=���=���="+�=���=\��=��=�.�=���=H��=x�=
t�=���=�u�=���=�� >�j>T>��>7�>E>�z>.�>u�>��>&n>B>�>5�>��>gg>{8>3>��>��>��>��>��>��> >�">�,>=,>|>��>2�>ǀ>� >�� >s >�   �   ��=���=���=�<�=��=��= �=<N�=���=��=���=�N�=��=@�=�0�=v��=� �=���=
 >�� >m>�>\�>!�>Y@>Rt>G�>�>��>1b>5>��>j�>R�>�W>�(>�> �>��>��>��>��>	�>
>)>�'>)>7>B�>��>��>X&>�� >�( >�   �   
`�=�!�=��=���=�`�=�L�=~e�=���=�F�=��=lA�=J��=�a�=�S�=n{�=|��=�9�=D��= >x� >�s>L>t�>�>R2>va>�w>jw>.c>�>>R>�>��>�_>)> �>u�>6�>�>��>&�>%�>��>K�>		>�> >�>��>Z�>ܐ>~7>�� >D >�   �   |��=��=�Z�=!�=L��=��=�	�=�\�=���=���=��=�H�=���=���=���=�7�=D��=���=	4 >�� >>y
>>N�>_>�B>�Q>*J>Y/>�>��>�>�R>�>z�>�>��>zp>�e>h>!v>��>C�>q�>�>�>�>�>_>Y�>>�>@S>�� >%p >�   �   �( >�3�=��=��=���=��=���=�<�=���=p��=���=X�=��=ލ�=L��=���=��=�c�=�Z >%� >��>>�u>��>A�>#>�>�>�>C�>�x>D5>Y�>��>5t>$D>� >�>�>U>$>aD>�k>r�>�>��> �>B
>u>��>�>Yx>>� >�   �   �{ >
��=���=���=P��=��=���=L�=$��=��=l��=��=���=Vh�=|\�=xt�=���=j��=�� >�>��>�>Yj>��>��>��>W�>��>q�>NU>u>��>Tw>�0>�� >�� >� >�� >F� >b� >s� >�� >!>�T>��>��>��>��>�>��>�>�>V>�� >�   �   �� >ec >���=���=4��=>��=j�=��=^�=X��=t��=X1�=��=�_�=�;�=�8�=@J�=�1 >	� >w=>ΰ>k>#\>؎>�>��>Ҕ>Ij>G.>�>j�>w>>�� >�� >_ >�- >n >:  >H > >�H >@� >�� >>�N>��>��>:�>4>�>��>�>H�>�A>�   �   �=>�� >d >L��=���=`�=�a�=��=vc�=�-�=b.�=�e�=���=jj�=�+�=�
�=L��=�y >8� >�a>�>�>bK>lm>Iw>i>�C>4
>��>�i>/>'� >R >L  >�x�=��=���=���=���=$�=V��= >z\ >.� >�
>z^>��>��>>�$>h$>^>��>�>�   �   դ>�K>�� >�} >x >4b�=���=�#�=��=���=F{�=��=���=�}�=x#�=j��=jY >
� >)>̅>��>.>�8>�I>uB>}#>�>Τ>�K>�� >�} >n >b�=d��=�#�=ڼ�=���=*{�=أ�=t��=�}�=f#�=\��=bY >� >)>ʅ>��>/>�8>�I>wB>�#>�>�   �   :
>�>�i>9>2� >%R >X  >�x�=��=��=���=���=$�=f��= >\ >4� >�
>�^>��>��>>�$>g$>]>��>�>�=>�� >d ><��=���=L�=�a�=���=bc�=�-�=J.�=le�=x��=^j�=�+�=�
�=>��=�y >4� >�a>�>�>dK>om>Lw>i>�C>�   �   Nj>N.>�>q�>�>>�� >�� >_ >�- >{ >D  >R >$ >�H >J� >�� >>�N>��>��>;�>0>�>��>�>D�>�A>�� >]c >���=���=��=&��=R�=��=J�=B��=b��=@1�=��=�_�=�;�=�8�=,J�=�1 >� >t=>ΰ>l>%\>َ>�>��>֔>�   �   ��>x�>RU>}>��>\w>�0>�� >�� >� >�� >O� >j� >x� >�� >)>�T>��>��>��>��>�>��>�>�>V>�� >�{ >���=���=���=B��= ��=���=L�=��=
��=T��=��=���=Fh�=p\�=jt�=���=b��=�� >�>��>�>Yj>��>��>��>]�>�   �   �>�>J�>�x>F5>_�>��>>t>*D>� >�>�>\>$>jD>�k>u�>�>��>�>C
>s>��>
�>Xx>>� >�( >�3�=��=���=���=
��=���=�<�=���=\��=���=B�=Ե�=ҍ�=:��=���=��=�c�=�Z >$� >��>>�u>��>C�>(>�>�   �   -J>_/>�>��>�>�R>�>��>�>��>p>�e>h>'v>��>E�>u�>�>�>�>�>\>Z�><�>BS>�� >#p >r��=���=�Z�=!�=>��=���=v	�=�\�=���=���=��=�H�=���=���=���=�7�=8��=���=4 >�� >
>x
>>N�>b>�B>�Q>�   �   kw>/c>�>>U>�>��>�_>!)>�>|�>9�>��>��>+�>)�>��>J�>		>�># >�>��>[�>ܐ>}7>�� >D >`�=�!�=��=ړ�=�`�=�L�=te�=���=�F�=��=dA�=@��=�a�=�S�=`{�=x��=�9�=>��=	 >v� >�s>M>u�>�>T2>za>�w>�   �   �>�>4b>	5>��>l�>T�>�W>�(>�>�>��>��>��>��>�>
>,>�'>#)>5>=�>��>ۄ>Y&>�� >�( >��=���=���=�<�=��=��= �=6N�=���=
��=���=�N�=��=>�=�0�=t��=� �=���=	 >�� >m>�>^�>!�>Z@>Tt>K�>�   �   ?�>�t>Z>H2>n >y�>��>�L>~>_�>S�>M|>-[>8C>q4>�->�,>�/>4>�6>x4>C+>�>a� >�� >� >8X >�
 >pj�=̴�=t��=(L�=Ʃ�=$�=��=Do�=6V�=l�=v��=�(�=���=ғ�=�{�= z�=�B >�� >`O>��>�>>¡>%�>4>�`>z>�   �   x> l>�P>x(>5�>	�>�>?B>M>��>�>�s>dS>}<>�.>)>y)>�->23>�6>46>5.>�>� >�� >`� >�` >
 >(~�=���=@�=�b�=���=>6�=���=z��=\k�=
��=���=.9�=z��=��=���=���=�E >� >�O>��>3<>X�>��>�.>MZ>�r>�   �   `>R>�4>\>
�><�>�`>M#>��>V�>��>UZ>�<>�(>�>�>�>�'>�0>f8>N;>�6>)>�>}� >� >�x >�. >
��=��=�S�=���=H�=�z�=��=>��=:��=0��=t��=>j�=��=h��=��=��=!M >�� >�O>/�>L5>�>D�>@>&G>�\>�   �   �8>�'>�>��>�>�k>].>�>��>�>U>%1>u>&>�>�>�>�>�,>�:>mC>�D>�<>�(>z>�� >;� >,Z >�
 > k�=f��=��=�s�=���=,|�=�1�=f�=6�=�S�=��=>J�=r��=���=(��=GY >*� >�O>��>*>i�>{�>�>(>�9>�   �   &>q�>��>ƛ>|d>(>��>��>$t>B>�>n� >G� >Y� >�� >�� >� >>r'>C=>CN>�W>�V>BJ>�0>D	>�� >�� >lI >r��=&H�=��=��=�}�=��=��=b��=
��=���=�$�=ڧ�=�N�=��=���=ji >4� >P>��>�>�l>��>��>��>�	>�   �   ��>[�>�>/M>�>��>��>FY>@">1� >_� >ش >�� >o� >�� >�� >�� >�� >� >�@>O[>Bn>�v>�r>a>aA>�>�� >є >�H >���=�P�=���=�0�=P��=6n�=�?�=�8�=:[�=*��=��=��=�`�=� >�| >�� >�O>İ>~>�P>Ɗ>��>b�>c�>�   �   Ny>�W>*>��>�>�t>�4>�� >�� >r� >�x >�e >M` >h >D| >ٚ >4� >h� >>	D>�i>��>=�>�>��>��>�Z>(>� >k� >�W >�
 >���=��=$��=:2�=��=X��=b��=;�=���=��=,��=�4 >�� >�� >�N>�>.�>�0>a>��>�>B�>�   �   (>��>��>��>N>:>�� >P� >�\ >�4 >� > >8 >�# >�B >�l >�� >2� >E>tG>2y>g�><�>��>	�>$�>3�>R|>GE>�>!� >�t >- >��=pa�=��=<��=���=���=���=�'�=<��= >�W >h� >w� >�L>f�>S�> >3>�H>�M>�B>�   �   ��>��>�h>L'>�� >�� >�Z >h  >"��=d��=pp�=�g�=Z��=n��=~ >�< >| >�� >�>vJ>��>��>�>=>�>�	>y�>��>��>�h>R'>�� >�� >�Z >q  >2��=v��=zp�=�g�=b��=x��=� >�< >| >�� >�>yJ>��>��>�><>�>�	>u�>�   �   K|>@E>�>� >�t >- >���=`a�=��=,��=���=���=���=�'�=4��= >�W >g� >t� >�L>d�>R�>>3>�H>�M>�B>(>��>��>��>"N>@>�� >Y� >�\ >5 >� > >< >�# >�B >�l >�� >2� >L>tG>2y>g�>9�>��>�>#�>1�>�   �   (>�� >c� >�W >�
 >���=��=��=*2�=��=L��=V��=
;�=���=��=��=�4 >�� >�� >�N>�>+�>�0>
a>��>�>E�>Vy>�W>*>��>�>�t>�4>�� >�� >y� >�x >�e >T` > h >G| >� >8� >i� >>D>�i>��>>�>�>��>��>�Z>�   �   �� >͔ >�H >���=�P�=���=�0�=<��=(n�=�?�=�8�=2[�= ��=��=��=�`�=� >�| >�� >�O>ð>|>�P>Ȋ>��>c�>f�>��>^�>�>4M>�>��>ĕ>LY>F">7� >g� >ߴ >�� >s� >�� >�� >�� >�� >� >�@>S[>?n>�v>�r>a>]A>�>�   �   � >fI >l��=H�=���=��=�}�=��=���=X��=���=���=�$�=Χ�=�N�=��=���=ki >2� >P>��>�>�l>��>��>��>�	>*>u�>��>ʛ>�d>(>��>��>*t>B>�>t� >J� >_� >�� >�� >� >
>u'>E=>EN>�W>�V>BJ>�0>@	>�� >�   �   'Z >�
 >k�=\��=��=zs�=���=|�=�1�=`�=*�=�S�=޹�=4J�=h��=���=$��=GY >'� >�O>��>*>h�>}�>�>(>�9>�8>�'>�>��>�>l>_.>�>��>�>U>*1>y>*>�>�>�>�>�,>�:>qC>�D>�<>�(>w>�� >9� >�   �   �. >��=��=�S�=���=F�=�z�=��=:��=4��=(��=j��=6j�=~�=b��=��=��= M >�� >�O>/�>M5>�>E�>=>*G>�\>`>R>�4>^>
�>>�>�`>L#>��>[�>��>WZ>�<>�(>�>�>�>�'>�0>g8>N;>�6>)>�>w� >� >�x >�   �    >&~�=���=>�=�b�=���=@6�=���=n��=Xk�=��=���=(9�=t��=��=���=���=�E >� >�O>��>3<>Z�>��>�.>MZ>�r>x>!l>�P>w(>6�>
�>�>@B>N>��>�>�s>hS>|<>�.>)>y)>�->33>�6>46>7.>�>� >�� >_� >�` >�   �   �
 >rj�=ʴ�=v��=&L�=̩�=�=��=Bo�=8V�=l�=r��=�(�=���=Г�=�{�=z�=�B >�� >`O>��>�>>��>%�>4>�`>z>?�>�t>Z>H2>n >{�>��>�L>~>`�>S�>L|>-[>;C>o4>�->�,>�/>4>�6>}4>C+>�>e� >�� >� >;X >�   �    >*~�=���=D�=�b�=���=F6�=���=t��=Zk�=��=���=*9�=~��=��=���=ā�=�E >� >�O>��>4<>Z�>��>�.>PZ>�r>x> l>�P>z(>5�>	�>�>AB>N>��>�>�s>eS>}<>�.>�(>y)>�->43>�6>56>9.>�>� >�� >a� >�` >�   �   �. >��=��=�S�=���=N�=�z�=��=B��=@��=4��=t��=<j�=��=n��=��=��=#M >�� >�O>2�>N5>�>F�>?>'G>�\>`>R>�4>_>
�>>�>�`>M#>��>W�>��>VZ>�<>�(>�>�>�>�'>�0>l8>R;>�6>)>�>|� >� >�x >�   �   .Z >�
 >"k�=l��=��=�s�=���=0|�=�1�=r�=<�=�S�=��=BJ�=v��=���=0��=LY >,� >�O>��>*>h�>�>�>(>�9>�8>�'>�>��>�>l>_.>�>��>�>U>,1>y>)>�>�>�>�>�,>�:>qC>�D>�<>�(>z>�� >>� >�   �   �� >oI >v��=0H�=��=��=�}�=��=��=n��=��=���=�$�=ާ�=�N�=��=���=oi >8� >P>��>�>�l>�>��>��>�	>*>t�>��>ʛ>�d>(>��>��>)t>B>�>t� >I� >]� >�� >�� >� >>v'>H=>FN>�W>�V>DJ>�0>E	>�� >�   �   �� >Ք >�H >���=�P�=���=�0�=R��=Bn�=�?�=�8�=H[�=2��=��= ��=�`�=� >�| >�� >�O>Ȱ>~>�P>Ȋ>��>e�>f�>��>_�>�>3M>�>��>Õ>JY>G">3� >e� >� >�� >t� >�� >�� >�� >�� >� >�@>W[>Fn>�v>�r>a>dA>�>�   �   (>� >l� >�W >�
 >ȁ�=&��=.��=D2�=��=b��=n��= ;�=���=��=8��=�4 >�� >�� >�N>�>0�>�0>a>��>�>G�>Ty>�W>*>��>�>�t>�4>�� >�� >x� >�x >�e >R` > h >K| >� >;� >l� >>D>�i>��>C�>
�>��>��>�Z>�   �   X|>KE>�>&� >�t >- >��=|a�=��=H��=��=���= ��=�'�=H��= >�W >m� >{� >M>i�>V�>>3>�H>N>�B>(>��>��>��>N>?>�� >U� >�\ > 5 >� > >< >�# >�B >m >�� >5� >K>uG>7y>p�>E�>��>�>)�>9�>�   �   ��>�>�h>W'>� >�� >[ >t  >>��=���=�p�=h�=l��=���=� >�< >| >�� >�>|J>��>ý>	�>?>�>�	>x�>��>��>�h>R'>�� >�� >�Z >n  >4��=r��=|p�=�g�=b��=z��=� >�< >| >�� >�>zJ>��>Ƚ>�>B>�>�	>~�>�   �   (>��>��>��>'N>E>�� >[� >�\ >5 >� > >A >�# >�B >m >�� >5� >O>wG>8y>m�>>�>��>
�>(�>6�>R|>DE>�>!� >�t >- >��=na�=��=2��=���=���=���=�'�=@��= >�W >l� >y� >�L>j�>X�>>3>�H>N>�B>�   �   Xy>�W>*>��>�>�t>�4>�� >�� >~� >�x >�e >U` >"h >O| >� >@� >k� >>D>�i>��>?�>�>��>��>�Z>(> � >h� >�W >�
 >���=��=$��=:2�=��=X��=`��=;�=���=��=.��=�4 >�� >�� >�N>�>1�>�0>a>��>�>K�>�   �   ��>c�>	�>9M> >��>ɕ>PY>K">;� >i� >� >�� >y� >�� >�� >�� >�� >� >�@>U[>En>�v>�r>a>bA>�>�� >ϔ >�H >���=�P�=���=�0�=H��=<n�=�?�=�8�=:[�=(��=��=��=�`�=� >�| >�� >�O>ʰ>�>�P>̊>��>h�>k�>�   �   ,>y�>��>͛>�d> (>��>�>/t>B>�>y� >L� >_� >�� >�� >� >>y'>H=>DN>�W>�V>BJ>�0>B	>�� >� >hI >n��="H�=��=��=�}�=��=���=`��=��=���=�$�=ԧ�=�N�=��=���=ni >7� >P>��>�>�l>�>��>��>�	>�   �   �8>�'>�>��>�>l>b.>�>��>#�>U>,1>}>,>�>�>�>�>�,>�:>rC>�D>�<>�(>|>�� >=� >*Z >�
 >k�=d��=��=�s�=���=(|�=�1�=j�=2�=�S�=��=>J�=p��=���=*��=KY >,� >�O>��>*>m�>~�>�>(>�9>�   �   `>R>�4>_>�>A�>�`>P#>��>\�>��>[Z>�<>�(>�>�>�>�'>�0>l8>Q;>�6>)> >{� >� >�x >�. >��=��=�S�=���=L�=�z�=��=@��=8��=.��=r��=>j�=��=f��=��=��=!M >�� >�O>2�>O5>�>H�>C>,G>�\>�   �   x>!l>�P>|(>:�>�>�>CB>O>��>�>�s>gS>{<>�.>)>w)>�->23> 7>56>5.>�>� >�� >_� >�` > >,~�=���=@�=�b�=���=>6�=���=t��=Pk�=��=���=(9�=|��=��=���=���=�E >� >�O>��>5<>]�>��>�.>OZ>�r>�   �   mt>�k>^S>",>��>��>0q>�#>��>�>5>� >b� >!r >�D >�" >� >� >���=� >Y >� >�. >< >�E >�I >cG >�= >- >� >
��=v��=�w�=l=�=�=$��=���=��=��=D�=П�=_ >�R >ģ >�� >dW>R�>>�d>��>��>O,>WT>�l>�   �   �l>d>�K>�$>|�>��>|j>�>��>~>�0>�� >ҧ >�p >D ><# >= > >c >:
 >y >�% >H5 >,C >M >�Q >�O >F >l5 >d >l >���=j��=�K�=t�=T��=���=��=�=0I�=��=� >WR >M� >3� >4T>N�>W
>d_>��>V�>n%>.M>/e>�   �   OV>OM>�4>>��>ڜ>�V>>>�>%o>$>p� >j� >�k >qB >�$ >� >W >v >� >�% >7 >�H >@X >�c >i >�g >�^ >VN >c7 >1 >���=x��=w�=.A�="�=��=X�=� �=XX�=.��=� >Q >� >4� >�J>��>w�>�O>!�>N�>!>�7>$O>�   �   �1>>(>�>��>V�>�z>�6>\�>š>W>�>�� >\� >|d >�? >�& >� >1 >� >�+ >U> >PS >"h >Ez >և >�� >ڎ >�� >�v >�_ >C >Y" >���= ��=���=&S�=�6�=
0�=�B�=q�=V��=K >�N >,� >�� >Y;>D�>��>�5>�~>r�>/�>A><+>�   �   	 >P�>�>��>��>�L>B>��>}>�6>�� >Ƿ > � >�Z >e< >* >R# >1' >�3 >wG >|_ ><y >+� >Ч >+� >~� >� >� >t� >�� >.x >=V >�1 >| >^��=2��=�z�=di�=fp�=R��=���=� >�K >�� >�� >�&>Tw>�>>X>��>��>h�>��>�   �   ��>J�>2�>�|>M>�>5�>��>rP>
>|� >� >bp >�N >-8 >�- >
/ >�: >�N >4i >�� >�� >�� >�� >u� >�� >�>=� >�� >n� >B� >�� >�m >0F >�  >���=���= ��=���=��=���=t >rH >Ƃ >?� >'>�W>��>��>�(>�`>I�>O�>��>�   �   P~>Qs>a[>�7>
>��>X�>G[>0>�� >� >&~ >�Y >�@ >�3 >92 >`< >�P >m >e� >ϴ >�� >�� >>%4>YC>I>�D>�6>�>| >� >�� >8� >\ >�5 > >���=���=V��=� >� >�D >v >6� >-� >d3>�v>��>��>�%>�N>�k>�{>�   �   �2>�&>>��>�>B�>�V>�>� >q� >� >�\ >nA >�1 >{. >7 >�J >zh >ō >S� >G� >�>.;>�^>�z> �>I�>ђ>��>Wn>N>�&>� >�� >�� >Lo >�H >;* > >� >, >3# >h@ >Zh >,� >�� >�>(H>t�>�>��>�
>'$>�1>�   �   �>��>,�>Ý>(t>{D>%>�� >o� >�| >FV >[9 >�' >" >�( >�; >�Y >� >Q� >J� >�>vJ>�y>̢>��>�>��>!�>��>2�>ȝ>,t>�D>'>�� >t� >�| >JV >]9 >�' >" >�( >�; >�Y >� >P� >K� >�>uJ>�y>ʢ>��>�>��>�   �   ̒>��>Rn>N>�&>
� >�� >�� >Ko >�H >7* > >� >* >3# >e@ >\h >0� >�� >�>*H>v�>�>��>�
>+$>�1>�2>�&>$>��>�>H�>�V>�>� >w� >� >�\ >qA >�1 >|. >	7 >�J >wh >ƍ >Q� >E� >�>);>�^>�z>�>G�>�   �   �D>�6>�>w >� >�� >5� >\ >�5 >� >���=���=P��=� >� >�D >v >8� >-� >f3>�v>��>��>�%>�N>�k>�{>X~>Ws>b[>�7>#
>��>^�>K[>5>�� >� >)~ >�Y >�@ >�3 >:2 >a< >�P >m >b� >δ >�� >�� >{>4>VC>�H>�   �   7� >�� >j� >?� >�� >�m >*F >�  >���=���=��=���=��=���=s >rH >Ƃ >B� >(>�W>��>��>�(>�`>M�>T�>��>��>L�>4�>�|>M>�>9�>��>tP>>�� >� >cp >�N >,8 >�- >/ >�: >�N >2i >�� >�� >�� >�� >p� >}� >�>�   �   � >o� >|� >,x >:V >�1 >w >P��=,��=�z�=bi�=jp�=J��=���=� >�K >�� >�� >�&>Tw>�>>X>��>��>m�>��> >U�>�>��>��>M>G>��>}>�6>�� >ȷ >!� >�Z >e< >* >U# >/' >�3 >uG >{_ >=y >(� >Χ >%� >y� >� >�   �   �� >�v >�_ >C >S" >���=���=���=S�=|6�=0�=�B�=q�=R��=H >�N >-� >�� >W;>F�>��>�5>�~>u�>0�>C>@+>�1>C(>�>��>Y�>�z>�6>_�>ǡ>W>�>�� >[� >{d >�? >�& >� >/ >� >�+ >S> >QS >h >Ez >ч >�� >َ >�   �   �^ >TN >`7 >0 >���=p��=w�=$A�=�=��=X�=� �=VX�=*��=� >Q >� >7� >�J>��>w�>�O>!�>P�> >�7>(O>OV>PM>�4>>��>ڜ>�V>@>�>'o>$>o� >l� >�k >nB >�$ >� >U >v >� >�% >7 >�H >@X >�c >i >�g >�   �   F >l5 >b >m >���=l��=�K�=j�=R��=���=��=�=,I�=��=� >SR >O� >4� >2T>L�>U
>d_>��>X�>q%>.M>0e>�l>d>�K>�$>z�>��>~j>�>��>
~>�0>�� >ҧ >�p >D >@# >< > >b >8
 >{ >�% >H5 >,C >M >�Q >�O >�   �   �= >- >� >��=n��=�w�=j=�=��= ��=���=��=��=D�=̟�=\ >�R >ģ >�� >bW>Q�>>�d>�>��>N,>WT>�l>qt>�k>[S>#,>��>��>1q>�#>��>�>5>� >c� >%r >�D >�" >� >� >���=� >[ >� >�. >< >|E >�I >cG >�   �   F >j5 >e >o >���=p��=�K�=n�=T��=���=��=�=(I�=��=� >UR >M� >8� >3T>M�>W
>f_>��>W�>p%>2M>1e>�l>d>�K>�$>{�>��>}j>�>��>~>�0>�� >ϧ >�p >D >@# >> > >c >:
 >z >�% >L5 >,C >M >�Q >�O >�   �   �^ >ZN >c7 >2 >���=x��=w�=0A�=&�=��=Z�=� �=XX�=0��=� >Q >� >7� >�J>��>z�>�O>"�>N�> >�7>%O>SV>OM>�4>>��>ڜ>�V>A>�>(o>$>r� >k� >�k >qB >�$ >� >X >w >� >�% >7 >�H >CX >�c >i >�g >�   �   �� >�v >�_ >C >\" >���=
��=���=,S�=�6�=0�=�B�=q�=^��=M >�N >0� >�� >Z;>G�>��>�5>�~>t�>3�>@>=+>�1>C(>�>��>Z�>�z>�6>_�>ȡ>W>�>�� >\� >}d >�? > ' >� >4 >� >�+ >V> >XS >"h >Gz >և >� >܎ >�   �   �� >w� >�� >1x >?V >�1 > >^��=:��=�z�=ji�=vp�=Z��=���=� >�K >�� >�� >�&>Uw> �>>X>��>��>k�>��>
 >R�>�>��>��>M>D>��>}>�6>�� >ɷ >!� >�Z >h< >* >Z# >2' >�3 >yG >�_ >Cy >/� >Ч >)� >� >� >�   �   ?� >�� >p� >E� >�� >�m >3F >�  >  >���=,��=
��=��=���=y >{H >̂ >F� >,>�W>��>��>�(>�`>L�>R�>��>��>N�>5�>�|>M>�>:�>��>uP>>�� >� >dp >�N >28 >�- >/ >�: >�N >7i >�� >�� >�� >�� >w� >�� >�>�   �   �D>�6>�>~ >� >�� >>� >
\ >�5 > >���=���=V��=� >� >�D >"v >9� >1� >g3>�v>��>��>�%>�N>�k>�{>V~>Vs>e[>�7>%
>��>[�>L[>5>�� >� >*~ >�Y >�@ >�3 >?2 >f< >�P >m >i� >մ >�� >�� >�>&4>]C>I>�   �   Ւ>��>Xn>N>�&>� >�� >�� >Ro >�H >?* > >� >/ >;# >n@ >ah >3� >�� >�>,H>w�>�>��>�
>+$>�1>�2>�&>!>��>�>F�>�V>�>� >v� >� >�\ >rA >�1 >�. >7 >�J >~h >ʍ >W� >L� >�>4;>�^>�z>$�>M�>�   �   !�>��>4�>̝>2t>�D>->�� >y� >�| >QV >c9 >�' >" >�( >�; >�Y >� >U� >P� >�>yJ>�y>͢>��>
�>��> �>��>0�>ɝ>.t>D>%>�� >w� >�| >LV >_9 >�' >" >�( >�; >�Y >� >W� >N� >>~J>�y>Ң> �>�>��>�   �   �2>�&>$>��>
�>J�>�V>�>� >{� >� >�\ >rA >�1 >�. >7 >�J >}h >ɍ >U� >H� >�>.;>�^>�z> �>L�>ђ>��>Un>N>�&>� >�� >�� >Qo >�H ><* > >� >1 >7# >o@ >ah >3� >�� >�>/H>{�>��>��>�
>.$>�1>�   �   Z~>Zs>f[>�7>*
>��>a�>O[>8>�� >� >.~ >�Y >�@ >�3 >?2 >h< >�P >m >f� >Դ >�� >�� >~>$4>YC>I>�D>�6>�>{ >� >�� >8� >\ >�5 >� >���=���=T��=� >� >�D > v >;� >2� >j3>�v>��>��>�%>�N>�k>�{>�   �   ��>Q�>5�>�|>M>�>=�>>zP>>�� >� >gp >�N >48 >�- >/ >�: >�N >4i >�� >�� >�� >�� >s� >�� >�>=� >�� >k� >B� >�� >�m >/F >�  >  >���=$��= ��=��=���=w >zH >̂ >F� >->�W>á>��>�(>�`>O�>T�>��>�   �    >U�> �>��>��>M>H>��>}>�6>�� >η >#� >�Z >j< >* >W# >0' >�3 >zG >�_ >>y >,� >Ч >$� >}� >� >� >s� >� >.x >>V >�1 >{ >V��=2��=�z�=di�=np�=T��=���=� >�K >�� >�� >�&>Yw>"�>>!X>��>��>n�>��>�   �   �1>D(>�>��>\�>�z>�6>b�>ɡ>W>�>�� >_� >|d >�? > ' >� >2 >� >�+ >T> >RS >#h >Fz >ԇ >�� >ێ >�� >�v >�_ >C >Y" >���=���=���=$S�=�6�=0�=�B�=q�=\��=M >�N >0� >�� >[;>I�>��>�5>�~>u�>3�>C>@+>�   �   QV>PM>�4>>��>ޜ>�V>C>�>*o>$>s� >m� >�k >rB >�$ >� >W >w >� >�% >7 >�H >?X >�c >i >�g >�^ >TN >`7 >. >���=r��=w�=0A�="�=��=`�=� �=VX�=4��=� >Q >� >7� >�J>��>y�>�O>&�>P�>!>�7>'O>�   �   �l>d>�K>�$>~�>��>|j>�>��>
~>�0>�� >ҧ >�p >D >?# >= > >c >:
 >~ >�% >F5 >+C >M >�Q >�O >F >k5 >e >m >���=n��=�K�=t�=T��=���=��=�=,I�=��=� >VR >N� >6� >4T>N�>X
>h_>��>V�>p%>1M>2e>�   �   my>�r>Z>�/>=�>˨>`O>H�>N|>6	>Д >�" >Zo�=t��=��=ރ�=0%�=��=���=���=�(�=J{�=��=v\�=~��=`�=���=( >�Y >�� >G� >�� >I� >�� >�� >�� >�� >�� >W� >8� >E� >�� >�>�G>m}>��>}�>�=>�>o�>5�>�.>�U>Lo>�   �   �q>Rk>gS>�)>�>v�>�K>��>�z>�>X� >�$ >�t�=2��=��=���=�2�=B��=���=��=~;�=���=���=>p�=��=Fs�=���=�0 >�a >� > � >v� >M� >�� >�� >�� >�� >�� >�� >�� >�� >�� >�>uA>+v>��>+�>+5>4x>y�>5�>�%>M>�f>�   �   \Z>�U>�?>>��>{�>�A>0�>Bv>K>�� >v) >
��=���=�.�=d��=[�=J*�=��=T9�=s�=8��=p2�=���=+�=���=� >hJ >�y >� >ۻ >�� >� >�� >�� >P� >� >�� >�� >� >�� >� >Q>H.>�`>`�>v�>|>�]>�>��>z>�3>jN>�   �   �4>�2>|>;�>��>V�>�0>��>�n>�>�� >K1 >d��=���=�]�=���=x��=�s�=�o�=��=<��=@%�=
��=�	�=|��=( >�> >�s >�� >�� >�� >�� >�� >�� >� >}� >�� >� >�� >ʴ >H� >�� >e� >2>>>�t>v�>��>$3>�r>��>��>

>�&>�   �   �>>��>W�>��>�e>�>�>id>/>� >�; >���=x"�=֜�=7�=V��=��=���=*�=�E�=С�=��=B��=� >�? >�x >�� >� >�� >�>�>�>�>>� >�� >� >� >C� >3� >Τ >�� >5� >]� >O>B>�{>��>��>Z8>Fs>{�>2�>��>�   �   ��>�>߾>��>�z>�B>��>a�>�W>�� >� >�H >���=�^�=���=ғ�=�_�=N�=f^�=ލ�=P��=�8�=^��=y >�M >� >+� >�� >H>,>H:>$=>w5>�$>h>�� >@� >h� >٠ >� >7� >� >Ԙ >� >� >�>�9>�t>�>��>�+>;a>̍>D�>�   �   |>t�>Ӂ>�m>K><>!�>Y�>�H>/� >v� >W >m >���=�A�=���=���=t��=���=8,�=~�=��=p* >�f >�� >�� >�>�8>qX>kl>bt>`p>a>'H>�'>[>J� >u� >͓ >y >Ug >` >�e >�v >O� >l� >�� >�%>�a>��>�>�>Q?>�c>�   �   .>�=>�>>�1>�>��>s�>�{>8>� >� >nf >�) >���=ؠ�= p�=t]�=�i�=��=���= >�L >� >� >�� >V4>�c>^�>��>��>��>�>��>�m>�C>X>�� >>� >�� >�_ >:C >2 >�- >w6 >ML >/n >k� >�� >�>�D>D�>1�>��>�>�   �   -�>�>��>��>*�>�>�>"`>�&>6� >Y� >:v >�D >1 >g >��=���=�  >1 >>C >�s >(� >E� >">z[>g�>�>5�>�>��>��>/�>
�>�>&`>�&>8� >Y� >8v >�D >1 >e >��=���=�  >/ >9C >�s >$� >>� >">r[>e�>�>�   �   X�>��>��>��>�>��>�m>�C>X>�� >>� >�� >�_ >;C >2 >�- >|6 >TL >0n >p� >�� >�>�D>J�>7�>��>�>.>�=>�>>�1>�>��>v�>�{>8>� >� >mf >�) >���=̠�=�o�=r]�=�i�=��=���= >�L >�� >� >�� >Q4>�c>�   �   �8>oX>fl>_t>^p>a>$H>�'>Z>G� >u� >Γ >y >Vg >�` >�e >�v >S� >n� >�� >�%>�a>��>�>�>T?>�c>|>y�>ց>�m>K>?>%�>\�>�H>0� >u� >W >n >���=�A�=���=���=f��=���=0,�=~�=���=k* >�f >�� >�� >}>�   �   �� >F>�+>E:>=>u5>�$>c>�� ><� >k� >ݠ >� >8� >�� >Ԙ >� >� >�>�9>�t>�>��> ,>Aa>э>I�>��>�>�>��>�z>�B>��>b�>�W>�� >!� >�H >���=�^�=���=Г�=�_�=�M�=d^�=ҍ�=J��=�8�=R��=u >�M >� >(� >�   �   � >
� >�� >�>�>�>�><� >�� >� >� >F� >3� >Ф >�� >6� >a� >R>B>�{>��>��>]8>Gs>��>7�> �>�>>��>W�>��>�e>�>�>id>0>	� >�; >���=x"�=Ԝ�=7�=X��=��=���= �=�E�=С�=~�=<��=� >�? >�x >�   �   �s >�� >�� >�� >�� >�� >�� >� >{� >�� >� >�� >ɴ >I� >�� >d� >5>>>�t>y�>��>&3>�r>��>��>

>�&>�4>�2>~>>�>��>Y�>�0>��>�n>�>�� >J1 >d��=���=�]�=���=x��=�s�=�o�=��=<��=:%�=���=�	�=p��=( >�> >�   �   gJ >�y >�� >ڻ >�� >� >�� >�� >P� >� >�� >�� >� >�� >� >O>M.>�`>_�>x�>}>�]>�>��>{>�3>mN>aZ>�U>�?>>��>{�>�A>0�>Bv>M>�� >u) >��=���=�.�=d��=[�=H*�=��=J9�=s�=8��=t2�=���=�*�=���=� >�   �   �0 >�a >�� >�� >v� >J� >�� >�� >�� >�� >�� >�� >�� >�� >�� >�>wA>,v>��>*�>-5>4x>z�>9�>�%>M> g>�q>Tk>cS>�)>�>w�>�K>��>�z>�>W� >�$ >�t�=6��=��=���=�2�=@��=���=��=�;�=���=���=:p�=��=@s�=���=�   �   ( >�Y >�� >G� >�� >I� >�� >�� >�� >�� >�� >Y� >7� >D� >�� >�>�G>n}>�>|�>�=>�>o�>6�>�.>�U>Oo>my>�r>Z>�/>:�>ɨ>`O>H�>L|>7	>ϔ >�" >Zo�=���=��=��=*%�=
��=���=���=�(�=J{�=��=p\�=|��=`�=���=�   �   �0 >�a >� >� >v� >O� >�� >�� >�� >�� >�� >�� >�� >�� >�� >�>wA>-v>��>*�>,5>4x>z�>6�>�%>M>g>�q>Tk>fS>�)>�>y�>�K>��>�z>�>X� >�$ >�t�=8��=��=���=�2�=F��=���=��=�;�=���=���=<p�=��=Fs�=���=�   �   hJ >�y > � >޻ >�� >� >�� >�� >O� >� >�� >�� >� >�� >	� >Q>N.>�`>`�>w�>~>�]>�>��>{>�3>nN>aZ>�U>�?>>��>{�>�A>2�>Cv>N>�� >w) >��=���=�.�=l��="[�=P*�=��=P9�=&s�=@��=x2�= ��=+�=���=� >�   �   �s >�� >�� >�� >�� >�� >�� >� >}� >�� > � >�� >ɴ >I� >�� >h� >;>>>�t>x�>��>(3>�r>��>��>
>�&>�4>�2>|>>�>��>Y�>�0>��>�n>�>�� >O1 >h��=���=�]�=���=���=�s�=�o�=��=F��=H%�=��=�	�=~��=+ >�> >�   �   �� >� >�� >�>�>�>�>?� >�� >� >� >K� >3� >Ҥ >�� >:� >c� >R>B>�{>��>��>^8>Js>��>6�>�>�>>��>Y�>��>�e>�>
�>nd>2>� >�; >���=~"�=��=7�=`��=$��=���=0�=F�=ޡ�=��=F��=� >�? >�x >�   �   �� >M>,>J:>&=>{5>�$>g>�� >E� >m� >� >� >9� >� >֘ >� >"� >�>�9>�t>�>��>�+>?a>ύ>I�>��>�>߾>��>�z>�B>��>d�>�W>�� >%� >�H >���=�^�=���=��=�_�=N�=n^�=ލ�=^��=�8�=f��=z >�M >� >.� >�   �   �8>vX>nl>et>ep> a>*H>�'>`>N� >{� >ғ >y >Yg >�` >�e >�v >U� >r� >�� >�%>�a>��>�>�>U?>�c>|>y�>ց>�m>K>@>$�>_�>�H>3� >{� >W >o >���=�A�=���=���=z��=��=B,�="~�=��=x* >�f >�� >�� >�>�   �   `�>��>��>��>�>��>�m>�C>^>�� >C� >�� >�_ >?C >2 >�- >�6 >SL >2n >p� >�� >�>�D>H�>7�>��>�>.>�=>�>>�1>�>��>v�>�{>8>� >� >sf >�) >���=��=p�=�]�=�i�="��=���= >M >	� >� >�� >Y4>�c>�   �   7�>�>��>��>2�>�>�>'`>�&><� >[� >Av >�D >4 >n >��=���=�  >4 >=C >�s >)� >E� >">y[>g�>�>3�>�>��>��>.�>
�>�>(`>�&>:� >[� >Av >�D >8 >n >*��=���=�  >8 >BC >�s >1� >J� >">|[>m�>�>�   �   .>�=>�>>�1>�>��>{�>�{>8>� >� >tf >�) >���=��=
p�=�]�=�i�= ��=���= >�L >� >� >�� >V4>�c>]�>��>��>��>�>��>�m>�C>\>�� >A� >�� >�_ >AC >2 >�- >�6 >WL >7n >v� >�� >�>�D>N�>;�>��>�>�   �   #|>}�>ف>�m>K>B>'�>`�>�H>5� >y� >W >n >���=�A�=���=���=n��= ��=8,�=~�=��=q* >�f >�� >�� >�>�8>rX>jl>ct>ap>a>'H>�'>`>L� >{� >ғ >y >\g >�` >�e >�v >Y� >s� >�� >�%>�a>��>�>�>X?>�c>�   �   ��>�>�>Ť>�z>�B>��>e�>�W>�� >#� >�H >���=�^�=���=ܓ�=�_�=N�=h^�=ލ�=T��=�8�=\��=v >�M >� >,� >�� >H>�+>G:>&=>x5>�$>i>�� >B� >n� >� >� >=� >�� >ۘ >
� >$� >�>�9>�t>�>��>,>Ba>ҍ>K�>�   �   �>> �>[�>��>�e>�>�>md>4>� >�; >���=|"�=ޜ�=
7�=\��=��=���=.�=�E�=С�=��=@��=� >�? >�x >�� >� >�� >�>�>�>�>?� >�� >� >� >H� >7� >դ >�� >?� >e� >W>B>�{>��>��>a8>Js>��>9�>�>�   �   �4>�2>>?�>��>[�>�0>��>�n>�>�� >O1 >b��=���=�]�=���=|��=�s�=�o�=��=>��=<%�=��=�	�=|��=( >�> >�s >�� >�� >�� >�� >�� >�� >� >�� >�� > � >�� >˴ >I� >�� >k� >9>	>>�t>{�>��>+3>�r>��>��>
>�&>�   �   _Z>�U>�?>>��>~�>�A>2�>Ev>O>�� >x) >��=���=�.�=h��=[�=L*�=��=P9�=s�=6��=p2�=��=+�=���=� >hJ >�y > � >ۻ >�� >� >�� >�� >R� >� >�� >�� >� >�� >� >T>N.>�`>c�>{�>�>�]>��>��>~>�3>nN>�   �   �q>Tk>hS>�)>�>y�>�K>��>�z>�>X� >�$ >�t�=4��=��=���=�2�=B��=���=��=�;�=���=���=6p�=��=Fs�=���=�0 >�a >� >� >y� >M� >�� >�� >�� >�� >�� >�� >�� >�� >�� >�>xA>-v>��>,�>.5>5x>~�>6�>�%>M>g>�   �   �>n�>�n>#=>��>�>�>��>�� >eY >`_�=V�=���=d��=���=���=�(�=���=0��=���=R'�=���=�|�=�c�=e�=Ls�=ȃ�=$��=�? >"� >�>lQ>��>(�>��>��>�>k�>%�>��>�>P�>,�>��>M�>��>Z*>�]> �>��>�>O:>Jd>��>�   �   9�>Ɓ>'h>+8>��>�>>��>& >�] >�j�=��=���=<��=��=0��=C�=f��=
��=��=�D�=��=���=��= �=�=��=��=sH >� >�>�U>ǋ>��>��>�>��>��>�>f�>E�>c�>4�>�>��>��> >�P>��>��>1�>�.>�Y>�w>�   �   ?l>)k>VU>])>L�>z�>>F�>�>�i >v��=2F�=@�=���=���=L&�=���=.7�=$�=?�=���=/�=���=T��=��=���=��=0��=Bb >"� >'>�b>p�>��>q�>�>P�>��>��>�>�>�>��>��>��>��>�>�(>ba>s�>��>B>�9>�Z>�   �   �A>�F>�6>5>��>�>�>��>�>d} >���=���=X_�=�L�=�]�=���=��=,��=>��=0��=�*�=Ի�=�w�=TU�=�H�=�G�=�F�=� >ҋ >4� >h;>'x>|�>h�>��>��>Ʋ>�>�>�n>y[>�O>M>�U>Sj>@�>��>��>!>^>�>��>S>%+>�   �   �>>�>�>�>�s>T>�>f#>g� >m >X��=���=8��=��=(9�="��=�n�=�_�=d��=���=Fx�=�/�=��=
��=���=���=�\ >_� >>*a>��>�>4�>��>͵>ĝ>>�]>J=>�!>�>K>4>>�3>G\>�>��>?	>�I>��>��>��>�   �   ��>J�>��>G�>�>�a><>.�>�5>`� >�0 >�T�=S�=g�=���=���=F��=RH�=�@�=,o�=���=l\�=�=.��=$��=���=;@ >:� >'>lS>��>��>��>��>0�>1�>��>LY>",>c >�� >_� >_� >� >5� >�� >{� >">(^>ɠ>	�>�)>�g>�>�   �   �q>J�><�>��>�}>�L>�>K�>J>�� >ba >���=��=��=Fa�=L��=,p�=�>�=�@�=�s�=���=�^�=�	�=��=���= : >#� >�� >YQ>ޒ>��>3�>�>��>W�>b�>$f>->�� >̹ >� >*^ >SB >�5 >n9 >�M >�q >1� >	� >%(>�r>I�>{>�@>�   �   �>VE>�_>Uf>�W>�4>�>е>�^>1� >� >�+ >2��=���=l6�=Լ�=�l�=I�=\T�=���=���=�u�=�=\��=<J >� >�>C\>ס>��>:�>�>��>/�>�>��>E>� >/� >�k >�+ >���=���=rt�=0n�=,��=t��=" >�Y >�� >� >,F>U�>��>�   �   �>)�>�>�/>a/>�>/�>k�>Ss>�!>�� >
p >� >\��=��=&��=~q�=�\�=�q�=���=��=���=� >o >�� >[!>�s>%�>-�>�>�/>f/>�>0�>m�>Rs>�!>�� >p >� >P��=��=��=pq�=�\�=�q�=���=��=���=� >�n >�� >U!>�s>�   �   <\>ҡ>��>7�>�>��>.�>�>��>	E>� >6� >�k >�+ >���=���=�t�=@n�=8��=���=) >�Y >ɣ >� >4F>\�>��>�>]E>�_>Yf>�W>�4>�>ҵ>�^>0� >� >�+ >&��=z��=Z6�=ʼ�=|l�=I�=PT�=���=���=zu�=��=R��=3J >� >�>�   �   �� >TQ>ڒ>��>.�>�>��>V�>b�>%f>�->�� >ѹ >� >/^ >WB >�5 >x9 >�M >�q >6� >� >,(>�r>Q�>�>�@>�q>N�>@�>��>�}>�L>�>J�>J>�� >_a >���=��=��=6a�=B��=p�=�>�=�@�=�s�=���=�^�=�	�=���=���=�9 >� >�   �   7� >%>iS>��>��>��>��>/�>.�>��>PY>(,>f >�� >c� >b� >� >=� >�� >�� >">.^>Ѡ>�>�)>�g>��>��>M�>��>K�>�>�a>>>/�>�5>_� >�0 >�T�=S�=�f�=r��=���=8��=@H�=�@�=o�=���=b\�=��=��=��=���=7@ >�   �   �\ >Z� >>'a>�>�>4�>��>̵>ŝ>>�]>M=>�!>�>P>:>>�3>M\>"�>��>F	>�I>ȇ>ž>��>�>>�>��>�>�s>T>�>c#>g� >l >R��=���=2��=
��=$9�=��=�n�=�_�=V��=���=<x�=�/�=��=���=t��=���=�   �   � >Ћ >/� >d;>!x>y�>g�>��>��>Ų>�>�>�n>}[>�O> M>�U>Zj>B�>��>��>!>^>�>�>X>(+>�A>�F>�6>8>��>�>�>��>�>a} >���=���=R_�=�L�=�]�=���=��= ��=.��=&��=�*�=ʻ�=�w�=LU�=�H�=�G�=�F�=�   �   *��=>b >"� >'>�b>o�>��>n�>�>O�>��>��>
�>�>�>��>��>��>��>��>�(>ga>v�>��>F>�9>�Z>Al>+k>[U>_)>O�>|�>>F�>�>�i >r��=,F�=<�=���=���=F&�=���=,7�="�=?�=���=/�=���=N��=��=���=��=�   �   ��=sH >|� >�>�U>Ƌ>��>��>�>��>��>��>g�>E�>c�>5�>�>��>��> >�P>��>��>7�>�.>�Y>�w><�>ʁ>(h>,8>��>�>>��>$ >�] >�j�=��=���=:��=��=0��=C�=`��=��=��=�D�=��=���=��=�=���=��=�   �   "��=�? >!� >�>jQ>�>&�>��>��>�>j�>%�>��>�>P�>)�>��>P�>��>Z*>�]> �>��>�>N:>Hd>ā>�>n�>�n>&=>��>�>�>��>�� >eY >\_�=T�=���=j��=���=���=)�=���=0��=���=V'�=���=�|�=�c�=e�=Fs�=ă�=�   �   ��=tH >|� >�>�U>ɋ>��>��>�>��>��>��>g�>F�>d�>3�>�>��>��> >�P>��>��>6�>�.>�Y>�w>:�>ǁ>(h>,8>��>�>>��>& >�] >�j�=��=���=<��=��=4��=$C�=h��=��=��=�D�=
��=���=��=�=���=��=�   �   2��=Db >$� >(>�b>q�>��>p�>�>P�>��>��>
�>�>�>��>��>��>��>��>�(>fa>u�>��>F>�9>�Z>@l>-k>\U>a)>P�>}�>>H�>�>�i >~��=4F�=D�=���=���=T&�=���=67�=.�=?�=���=
/�=���=V��=��=���=��=�   �   � >Ջ >4� >j;>&x>�>j�>��>��>ʲ>�>�>�n>~[>�O>#M>�U>Yj>D�>��>��>!>^>�>�>X>(+>�A>�F>�6>9>��>�>�>��>�>f} >���=�=\_�=�L�=�]�=���=��=6��=B��=2��=�*�=ܻ�=�w�=ZU�=�H�=�G�=�F�=�   �   �\ >`� >>0a>��>!�>8�>��>ε>ŝ>>�]>L=>�!>�>S>:>>�3>I\>#�>��>D	>�I>ć>¾>��>�>>�>��>"�>�s>V>!�>j#>k� >q >b��=���=B��=��=:9�=,��=�n�=�_�=l��=���=Rx�=�/�=��=
��=���=���=�   �   =� >->mS>��>��>��>��>4�>4�>�>TY>),>g >�� >f� >e� >
� >>� >�� >�� >">-^>Ҡ>�>�)>�g>��>��>O�>��>I�>�>�a>@>2�>�5>d� >�0 >U�= S�=g�=���=���=R��=^H�=�@�=8o�=���=�\�=�=4��=$��=���=>@ >�   �   �� >\Q>�>��>7�>�>��>\�>f�>(f>�->�� >й >� >0^ >ZB >�5 >w9 >�M >�q >7� >� >+(>�r>M�>>�@>�q>M�>B�>��>�}>�L>�>Q�>J>�� >ha >���=*��=��=Pa�=`��=>p�=?�=�@�=�s�=��=�^�=�	�=��=���=: >&� >�   �   F\>ܡ>��>=�>�>��>1�>�>��>E>� >7� >�k >�+ >���=���=�t�=>n�=:��=���=) >�Y >ƣ >� >0F>Z�>��>�>[E>�_>[f>�W>�4>�>ֵ>�^>7� >� >�+ >:��=���=x6�=��=�l�="I�=lT�=Ό�=��=�u�=$�=h��=?J >� >�>�   �   (�>4�>�>�/>l/>�>3�>p�>Vs>�!>�� >p >� >\��=��=*��=�q�=�\�=�q�=���=��=���=� >o >�� >X!>�s>"�>-�>�>�/>g/>�>0�>s�>Xs>�!>�� >p >� >n��=��=:��=�q�=�\�=�q�=���=��=���=� >o >�� >_!>�s>�   �   �>aE>�_>]f>�W>�4>	�>ӵ>�^>4� >� >�+ >0��=���=j6�=ڼ�=�l�=I�=`T�=���=���=�u�=�=\��=9J >� >�>C\>ء>��>;�>�>��>0�>�>��>E>"� >8� >�k >�+ >���=���=�t�=Nn�=H��=���=0 >�Y >ѣ >� >8F>_�>��>�   �   �q>S�>C�>��>�}>�L>�>N�>
J>�� >ca >���=��=��=Da�=T��=.p�=�>�=�@�=�s�=��=�^�=�	�=��=���=�9 >!� >�� >YQ>ޒ>��>4�>�>��>[�>g�>)f>�->�� >Թ >� >6^ >aB >�5 >~9 >�M >r >=� >� >3(>�r>V�>�>�@>�   �   ��>S�>��>N�>�>�a>B>3�>�5>c� >�0 > U�=S�=g�=���=���=H��=NH�=�@�=,o�=���=j\�= �=&��=��=���=<@ >:� >(>jS>��>��>��>��>6�>8�>�>TY>+,>k >� >k� >k� >� >B� >� >�� >">6^>٠>�>�)>�g>��>�   �   �>>�>��>!�>�s>X> �>h#>j� >o >\��=���=6��=��=.9�=&��=�n�=�_�=`��=���=Fx�=�/�=��=��=|��=���=�\ >^� >>,a>��>!�>6�>��>ӵ>ɝ>>�]>O=>�!>�>U>A>>�3>Q\>)�>��>N	>�I>ɇ>ʾ>��>�   �   �A>�F>�6>9>��>�>�>��>�>d} >���=���=Z_�=�L�=�]�=���=��=.��=<��=0��=�*�=ֻ�=�w�=TU�=�H�=�G�=�F�=� >ы >4� >i;>%x>{�>h�>��>��>ɲ>�>�>�n>�[>�O>(M>�U>\j>H�>��>��>!!>^>�>�>]>++>�   �   Bl>.k>[U>a)>R�>~�>>I�>�>�i >x��=2F�=:�=���=���=L&�=���=47�=$�=?�=���=/�=���=V��=��=���=��=0��=@b >#� >(>�b>p�>��>s�>�>P�>��>��>�>!�>�>��>��>��>��>��>�(>ja>z�>��>I>�9>�Z>�   �   :�>Ɓ>)h>/8> �>�>>��>' >�] >�j�=��=���=6��=��=0��=C�=b��=��=��=�D�=��=���=��=�=�=��=��=sH >~� >�>�U>Ƌ>��>��>�>��>��>��>j�>H�>f�>6�>�>��>��>#>�P>��>��>5�>�.>�Y>�w>�   �   �>��>�>ZR>}�>yu>��>�>�B >���=���=P��=��=4]�=H��=.��=P��=�#�=���=X!�=��=֓�=���=�3�=\��=̊�=tM�=��=���=E� >�1>��>X>7i>v�>­>��>L�>ω>xk>;L>�0>�>�>V>B(>7F>�o>ע>��>�>BO>�>d�>�   �   `�>2�>Z�>�M>0�>fu>6�>h>�I > ��=���=��=�0�=��=��=��=B��= O�=��=�M�=���=L��=^��=LZ�=
��=D��=6j�=��=D��=q� >�7>n�>� >ph>��>��>Ѩ>&�>�~>�^>�=>~ >K>>�>*>2>\>��>��>�>�?>�q>��>�   �   3�>��>�u>�@>h�>5u>��>�*>9^ >~��=�+�=�T�=l��=,��=q�= ?�=8[�= ��=h��=4��=�[�=�;�=*e�=���=X^�=Z�=���=2i�=N��=s� >dI>V�>%>#f>ԋ>��>��>�}>�]>�7>�>��>��>�>x�>��>=�>� >wV>@�>	�>>�G>\r>�   �   !X>	d>	V>�*>�>�t>$�>l@> >ZV�=��=j��=� �=(��=@$�=d��=0$�=Ξ�=�s�= ��=�,�=��=�'�=v��= 	�=|��=fI�=��=p- >P� >�e>��>�+>Ob>�}>�>�p>BQ>I'>B�>q�>�>�>6m>�i>�v>�>�>��>�9>�>��>P>M6>�   �   �>l+>�*>�>%�>=s>��>]>�� >j��=�*�=h��=$��=:g�=�=F��=�1�=���="��=���=�D�=��=�-�=8z�=���=�u�=B�=�~�=^o >S
>H�>�>�4>�\>j>�_>dA>>��>�>rf>~2>�	>�� >�� >�� >]>+<>�x>��>�>;\>��>`�>�   �   ��>J�>��>��>��>�p>>�~>�� >�+ >���=T�=���=�r�=9�=^7�=�y�=�=L��=�=��= c�=~k�=���=t�=�p�=���=# >� >�H>h�>�
>�>>�U>{Q>�5>3>��>�>o4>�� >�� >kw >%U >�F >�M >�i >�� >�� >�)>�>7�>�1>>�   �   �X>��>�>��>��>Ml>I>֣>�>)z >j��=�>�=��=���=��=ڙ�=v��=���=�o�=��=��=t��=���=X��=<�=���=���= � >f>7�>��>`)>�I>�L>~4>�>��>�n>�>�� >Y] >  >֜�=�D�=��=� �=dW�=,��=% >7| >�� >�E>ͫ>r	>�   �   .�>d9>2p>�>��>f>&>�>QU>#� >�7 >�9�=�=��=Z��=@�=,��=X*�=(�=pK�=r��=t�=Z�=�g�=���=
��=#t >�� >�w>��>� >�I>MT>�A>�>��>�s>�>3� >|+ >�=��=F)�=м�=��=���=x��=�!�=Z��= |�=;, >ޡ > >��>�   �   Uu>��>�%>�V>�i>^>�4>��>i�>�!>�� >� >1�=�5�=�W�=���=� �=,��=���=<�=8s�=`�=���=���=���=m| >�� >^u>��>�%>�V>�i>^>�4>��>h�>�!>� >� >
1�=�5�=�W�=���=� �=��=���=�=s�=H�=���=���=x��=d| >�� >�   �   �� >�w>��>� >�I>LT>�A>�>��>�s>�>:� >�+ >ր�=*��=\)�=��=:��=��=���=�!�=n��=|�=G, >� >>��>8�>l9>7p>�>��>f>&>�>OU>� >�7 >�9�=��=���=B��=0�=��=6*�=�=LK�=X��=t�=Z�=lg�=֍�=���=t >�   �   � >`>1�>��>\)>�I>�L>�4>�>��>�n>�>�� >b] >* >��=E�=��=� �=�W�=@��=% >A| >�� >F>ԫ>w	>�X>��>��>��>��>Ll>I>ԣ>�>%z >^��=�>�=���=���=��=ƙ�=b��=l��=�o�= ��=��=^��=l��=D��= <�=���=���=�   �    >޾ >�H>d�>�
>�>>�U>{Q>�5>4>��>�>w4>�� >� >rw >/U >�F >�M >�i >�� >�� >�)>&�>>�>�1>>��>N�>��>��>��>�p>>�~>�� >�+ >���=�S�=���=�r�=�8�=L7�=�y�=�=6��=��=Й�=c�=hk�=���=Z�=�p�=���=�   �   �~�=Yo >O
>F�>�>�4>�\>
j>�_>eA>>��>�>}f>�2>�	>�� >�� >�� >f>3<>�x>�>�>B\>��>g�>�>n+>�*>�>%�>@s>��>]>�� >`��=�*�=^��=��=.g�=��=:��=�1�=x��=��=��=�D�=t�=�-�=&z�=|��=�u�=:�=�   �   ���=m- >M� >�e>��>�+>Qb>�}>�>�p>EQ>P'>D�>x�>��>�>?m>�i>�v>�>#�>��>�9>�>��>U>S6>(X>
d>V>�*>�>�t>&�>k@> >XV�=��=`��=� �=��=4$�=X��=$�=���=�s�=��=�,�=��=�'�=h��=��=p��=`I�=�   �   ,i�=J��=p� >bI>T�>%>%f>ҋ>��>��>�}>�]>�7>�>��>��>�>�>��>B�>� >{V>E�>�>>�G>^r>7�>��>�u>�@>f�>4u>��>�*>7^ >~��=�+�=�T�=f��=&��=�p�=?�=4[�=��=Z��=(��=�[�=�;�="e�=���=F^�=L�=���=�   �   ��=@��=l� >�7>i�>� >nh>��>��>Ш>*�>�~>�^>�=>~ >N>>�>+>2>\>��>��>�>�?>�q>�>b�>4�>V�>�M>1�>ju>8�>f>�I > ��=���=��=�0�=��=��=��=<��=�N�=��=�M�=���=L��=V��=HZ�= ��=>��=0j�=�   �   ��=���=B� >�1>��>\>5i>s�>��>��>M�>ω>wk>:L>�0>�>�>X>B(>6F>�o>ע>��>�>@O>�>g�>�>��>�>[R>�>wu>��>�>�B >���=���=L��=��=8]�=F��=.��=L��=�#�=���=V!�=��=ғ�=���=�3�=X��=Ȋ�=vM�=�   �   ��=F��=o� >�7>n�>� >rh>��>��>Ө>(�>�~>�^>�=>~ >M>>�>+>2>\>��>��>�>�?>�q>�>b�>3�>[�>�M>1�>ju>8�>i>�I >��=���=��=�0�=��=��="��=N��=O�=��=�M�=���=P��=`��=NZ�=��=D��=4j�=�   �   4i�=V��=u� >dI>X�>%>(f>Ӌ>��>��>�}>�]>�7>�>��>��> �>~�>��>B�>� >yV>D�>�>>�G>^r>7�>��>�u>�@>h�>6u>��>�*>:^ >���=�+�=�T�=r��=2��=
q�=.?�=F[�=(��=p��=8��=�[�=�;�=2e�=���=V^�=X�=���=�   �   ��=u- >O� >�e>��>�+>Tb>�}>�>�p>FQ>S'>E�>w�>��>�>@m>�i>�v>�>"�>��>�9>�>��>Q>Q6>%X>d>V>�*>�>�t>'�>o@> >bV�=��=t��=� �=2��=N$�=r��=8$�=ڞ�=�s�=��=�,�=��=�'�=x��=	�=���=nI�=�   �   �~�=ao >V
>L�>�>�4>�\>j>�_>iA>>��>�>zf>�2>�	>�� >�� >�� >b>3<>�x> �>�>D\>��>f�>�>o+>�*>�>)�>Bs>��>
]>�� >r��=�*�=t��=.��=Fg�=�=V��=�1�=���=0��=��= E�=��=�-�=Bz�=���=�u�=L�=�   �   ( >� >�H>k�>�
>�>>�U>�Q>�5>6>��>�>t4>�� >� >sw >/U >�F >�M >�i >�� >�� >�)>#�>=�>�1>>��>N�>��>��>�>�p>%>�~>�� >�+ >���=T�=���=�r�="9�=t7�=�y�=,�=\��=�=���=4c�=�k�=���=x�=�p�=���=�   �   %� >l>:�>��>c)>�I>�L>�4>�>��>�n>�>�� >]] >* >��=E�=��=� �=zW�=>��=% >>| >�� >F>ӫ>w	>�X>��>��>��>��>Ql>M>ܣ>�>.z >v��=�>�=��=���=��=���=���=���=�o�=,��=��=���=���=f��="<�=���=���=�   �   �� >�w>��>� >�I>ST>�A>�>��>�s>�>:� >�+ >Ҁ�=*��=\)�=��=.��=
��=���=�!�=j��=|�=C, >� >>��>6�>l9>7p>"�>��>f>&>�>XU>*� >�7 >�9�=�="��=p��=Z�=F��=h*�=8�=�K�=���=4t�=4Z�=�g�=���=��=)t >�   �   cu>��>�%>�V>�i>^>�4>��>k�>�!>�� >� >1�=�5�=�W�=���=� �="��=���=2�=6s�=\�=���=���=���=k| >�� >^u>��>�%>�V>�i>^>�4>��>q�>�!>�� >� >.1�=6�=�W�=΢�=� �=<��=���=N�=Ps�=x�=���=���=���=s| >�� >�   �   =�>q9>:p>#�>��>f>&>�>TU>%� >�7 >�9�=��=��=`��=B�=,��=N*�= �=dK�=p��=t�=Z�=|g�=��=��=#t >�� >�w>��>� >�I>RT>�A>�>��>�s>>@� >�+ >��=<��=v)�=��=J��="��=���=�!�=���=.|�=M, >� >>��>�   �   �X>��>��>��>��>Ql>K>٣>�>*z >h��=�>�=��=���=���=ܙ�=|��=|��=�o�=��=��=r��=���=V��=<�=���=���=� >f>7�>��>b)>�I>�L>�4>�>��>�n>�>�� >j] >3 >���=$E�=��=� �=�W�=T��=% >J| >�� >F>٫>~	>�   �   ��>T�>��>��>�>�p>">�~>�� >�+ >���=
T�=���=�r�=9�=^7�=�y�=�=J��=�=ޙ�=c�=|k�=���=j�=�p�=���=" >� >�H>j�>�
>�>>�U>�Q>�5>;>��>�>~4>�� >
� >}w >8U >�F >�M >�i >�� >�� >�)>,�>C�>2>>�   �   �>s+>�*>�>+�>Bs>��>]>�� >n��=�*�=j��=$��=4g�=�=D��=�1�=���=��=���=�D�=��=�-�=4z�=���=�u�=B�=�~�=]o >S
>K�>�>�4>�\>j>�_>jA>>��>��>�f>�2>�	>�� >�� >�� >l>;<>�x>�>�>I\>��>h�>�   �   (X>d>V>�*>�>�t>'�>m@> >`V�=��=f��=� �="��=B$�=d��=,$�=Ȟ�=�s�=��=�,�=��=�'�=n��=��=v��=fI�=��=p- >Q� >�e>��>�+>Rb>�}>�>�p>IQ>V'>I�>~�>��>$�>Em>�i>w>"�>)�>��>�9>�>��>V>S6>�   �   8�>��>�u>�@>i�>6u>��>�*>9^ >���=�+�=�T�=h��=.��=q�="?�=8[�=��=`��=.��=�[�=�;�=,e�=���=X^�=X�=���=2i�=L��=t� >eI>Z�>%>&f>؋>��>��>�}>�]>�7>�>��>��>"�>��>��>G�>!>�V>I�>�>>�G>_r>�   �   f�>4�>[�>�M>4�>iu>5�>h>�I >��=���=��=�0�=��=��=��=@��=�N�=��=�M�=���=N��=X��=LZ�=��=B��=2j�=��=F��=q� >�7>n�>� >sh>��>è>Ѩ>&�>�~>�^>�=> >P>>�>,>2>	\>��>��>�>�?>�q>�>�   �   ��>��>�>Bj>�>�<>�`>�Z >�`�=.��=�+�=v{�=`��=\p�=L�=���= 5�=b�=�=�\�=P*�=�w�=�6�=�S�=<��=�J�=���=b��=h��=q >�>	�>@�>D >qK>~p>�u>Da>F:>O>p�>"�>Nj>�G>�5>6>�I>�n>�>��>g&>j>�>1�>�   �   *�>��>��>�e>��>?>9f>Hc >�x�=���=dP�=��=��=(��=���=|��="s�=���=�X�=.��=jh�=���=�o�=���=z��=�v�= �=��=��=c& >�>��>ˊ>��>�E>�g>.j>�R>�(>%�>��> �>0O>>+>>�>�+>sQ>��>��>'>?T>��>��>�   �   0�>~�>��>Y>��>:E>5v>�| >���=�N�=��=$�=��=A�=�+�=�s�=`*�=�]�=P�=X�= �=�d�=��=�'�=�{�=���=���=��=dc�=�C >�1>R�>-�>��>�4>AN>�G>�'>�>��>�t>F5>��>m�>a�>�>��>��>�3>Ky>��>>>�Y>\�>�   �   Xs>-�>0z>�C>U�>�N>o�>*� >�1�=���=tl�=V��=&��=4=�=<:�=��=�R�=\��=�H�=p��=�I�=ă�=P)�=�'�=�f�=v��=�<�=z��=2��=�s >R>Z>��>��>>�#>w>�>\�>T>�>&�>�{>wL>�1>\.>�B>�m>��>X�>�O>��>�>CB>�   �   �>�A>�G>�%>�>GZ>I�>e� >���=.��=V�=r��=��=B��=R��=�= ��=�$�=���=(!�=���=��=���=��=J��=j��=n3�=�q�=@��=5� >�|>�>̏>B�>^�>��>��>n}>�)>��>�m>V>�� >̑ >@q >!k >� >Ю >f� >L>]�>X>�{>|�>�   �   K�>k�>e>K�>�>�f>��>�>�> >��=�n�=ZE�=�$�=0%�="]�=���=Z��= �=���=6�=h��="��=RY�=� �=��=d;�=�]�=�m�='* >�� >=�>�6>>�>�>��>�\>a>��>�$>y� >�H >���=�X�=f	�=���="�=(��=� >�v >�� >d>K�>AL>�   �   %>�>I�>�>�>;s> >'d>�� >̌�=���=��=���=~��=O�=`��=���=�J�= �=�K�=R��=,��=0V�=���=���=
��=���=��=�� >�U>d�>S>�>*�>2�>�F>��>�r>�� >Sb >^��=��=��=�G�=���=���=
��=n�=x�=j�= >N� >�%>5�>�   �   ғ>�>�h>�>�>/~>�+>?�>�>�P >��=A�=���=���=�f�=x+�=�>�= ��=:}�=���=�H�=�:�=�{�=���=ȣ�=�`�=|�=s] >�>1�>�%>�o>Ռ>}>7C>z�>Zg>�� >�1 >��=��=��=h��=��=��=�r�=J��= �=��=���=��=2d�=�[ >�� >�   �   �� >�><>(b>�>ņ>�U>��>{>�� >|* >���=>R�=���=X��=~v�=v��=�"�=���=�+�= ��=0��=��=��=z��=��=�G >�� >�>C>,b>�>ņ>�U>��>{>�� >p* >���= R�=���=6��=Zv�=P��=|"�=���=�+�=ص�=��=���=��=Z��=��=�G >�   �   g] >�>*�>�%>�o>Ռ>}>:C>��>ag>�� >�1 >��=,��=,��=���=�=>��=�r�=t��=B �=8��=���=��=Pd�=\ >�� >ݓ>�>�h>�>��>0~>�+>;�>�>�P >���=�@�=օ�=���=�f�=X+�=�>�=֬�=}�=���=lH�=�:�=f{�=���=���=�`�=f�=�   �   ���=�� >�U>_�>
S>�>+�>4�>�F>��>�r>�� >cb >~��=:��="��=�G�=���=���=2��=2n�=��=��=# >]� >�%>@�>%>�>K�>�>�>;s>} >%d>�� >���=���=��=���=b��=�N�=D��=���=|J�=��=�K�=2��=��=V�=t��=���=��=l��=�   �   �m�=!* >�� >:�>�6>��>�>�>��>�\>m>��>�$>�� >�H >���=�X�=�	�=��=0"�=D��=� >�v >�� >(d>X�>LL>Q�>n�>h>M�>�>�f>��>�>�> >��=�n�=DE�=�$�=%�=]�=���=>��=��=h��=�=D��=��=2Y�=� �=��=N;�=�]�=�   �   �q�=0��=0� >�|>�>ʏ>C�>[�>��>��>v}>�)>��>�m>b>� >ؑ >Nq >.k >
� >ۮ >q� >L>g�>d>�{>��>�>�A>�G>�%>�>GZ>G�>c� >���=��=�U�=\��=س�=,��=6��=��=���=�$�=���=!�=���=n�=p��=��=,��=R��=b3�=�   �   p��=*��=�s >R>W>��>��>>�#>z>�>d�>T>�>/�>�{>L>�1>h.>�B>�m>��>_�>�O>��>�>MB>_s>1�>2z>�C>T�>�N>l�>'� >�1�=���=hl�=B��=��=$=�=.:�=Ԑ�=�R�=F��=�H�=T��=zI�=���=:)�=�'�=�f�=f��=�<�=�   �   ��=bc�=�C >�1>P�>*�>��>�4>@N>�G>�'>�>��>�t>M5>��>v�>l�>
�>��>��>�3>Ry>��>C>�Y>a�>5�>��>��>Y>��>7E>4v>�| >���=�N�=��=$�=ܜ�=A�=�+�=�s�=T*�=�]�=<�=X�=��=nd�=��=x'�=�{�=���=���=�   �   ��=��=_& >�>��>Ɋ>��>�E>�g>-j>�R>�(>%�>��>�>3O>C+>>�>�+>wQ>��>��>*>DT>��>��>.�>��>��>�e>��>?>9f>Hc >�x�=���=^P�=��=��=$��=���=p��=s�=���=�X�="��=bh�=���=zo�=x��=l��=�v�=��=�   �   Z��=j��=o >�>�>@�>E >qK>zp>�u>Ca>G:>O>n�>"�>Lj>�G>�5>6>�I>�n>
�>��>i&>j>�>3�>��>��>�>Bj>�>�<>�`>�Z >�`�=.��=�+�=t{�=`��=\p�=L�=��=5�=b�=�=�\�=T*�=�w�=�6�=�S�=6��=�J�=���=�   �   ��=��=b& >�>��>ˊ>��>�E>�g>.j>�R>�(>$�>��>�>1O>C+>>�>�+>vQ>��>��>*>BT>��>��>-�>��>��>�e>��>
?>;f>Jc >�x�=���=fP�=��=��=,��=���=���=,s�=���=Y�=.��=jh�=���=�o�=���=z��=�v�=��=�   �   ��=nc�=�C >�1>U�>,�>��>�4>?N>�G>�'>�>��>�t>M5>��>w�>i�>	�>��>��>�3>Ry>��>B>�Y>`�>7�>��>��>Y>��>;E>7v>�| >���=�N�=��=$�=��=A�=�+�=�s�=l*�=�]�=\�=&X�= �=�d�=��=�'�=�{�=���=���=�   �   ���=<��=�s >
R>]> �>��>>�#>}>�>a�>T>�>0�>�{>�L>�1>e.>�B>�m>��>^�>�O>��>�>IB>cs>2�>1z>�C>Z�>�N>p�>-� >�1�=��=�l�=`��=4��=F=�=P:�=���=S�=j��=�H�=|��=�I�=؃�=\)�=�'�=�f�=|��=�<�=�   �   �q�=H��=9� >�|>�>Ϗ>D�>_�>��>��>s}>�)>��>�m>c>� >֑ >Kq >+k >� >ۮ >q� >L>f�>d>�{>��>�>�A>�G>�%>�>MZ>M�>k� >���=8��=V�=���=���=R��=b��= �=��=�$�=��=6!�=��=��=���=��=P��=r��=z3�=�   �   �m�=.* >�� >@�>�6>Ȑ>�>$�>��>�\>k>��>�$>�� >�H >���=�X�=�	�=���=."�=@��=� >�v >�� >&d>U�>KL>T�>p�>i>Q�>�>�f>��>�>�> > ��=�n�=nE�=�$�=D%�=:]�=���=r��=�=���=L�=|��=8��=fY�=� �=��=l;�=�]�=�   �   ��=�� >�U>i�>S>�>/�>:�>�F>��>�r>�� >^b >t��=8��="��=�G�=���=���=$��=,n�=��=��= >X� >�%>?�>%>�>P�>�>�>Bs>� >0d>ģ >ڌ�=���=��=���=���=O�=���=���=�J�=6�=�K�=l��=H��=LV�=���=���=��=���=�   �   y] >�>5�>�%>�o>ی>}>:C>��>bg>�� >�1 >��="��=&��=���=�=.��=�r�=l��=8 �=.��=���=��=Fd�=\ >�� >ܓ>�>�h>�>��>7~>�+>H�>�>�P >��= A�=
��=���=�f�=�+�=�>�=��=P}�=̱�=�H�=�:�=�{�=���=֣�=�`�=��=�   �   �� >�>H>1b> �>̆>�U>��>{>�� >{* >���=4R�=���=V��=~v�=r��=�"�=���=�+�=���=&��=��=��=p��=��=�G >�� >�>D>0b>�>̆>�U>��> {>�� >�* >���=PR�=���=v��=�v�=���=�"�=��=�+�=��=N��=2��=�=���=��=�G >�   �   �>�>�h>�>��>5~>�+>@�>�>�P >��=A�=��=���=�f�=x+�=�>�=��=0}�=���=�H�=�:�=~{�=���=���=�`�=|�=r] >�>3�>�%>�o>ی>}>BC>��>ig>�� >�1 >��=D��=F��=���=4�=T��=s�=���=^ �=T��=���=��=^d�=\ >�� >�   �   #%>��>Q�>�>�>@s>� >,d>�� >̌�=���= ��=���=v��=�N�=`��=���=�J�=�=�K�=N��=$��=(V�=���=���=��=~��=
��=�� >�U>h�>S>�>3�>>�>�F>��>�r>�� >ib >���=T��=@��=H�=���=��=J��=Ln�=��=��=, >c� >�%>G�>�   �   Z�>v�>k>S�>�>�f>��>�>�> >��=�n�=XE�=�$�=*%�="]�=���=V��=��=���=0�=^��=��=JY�=� �=��=^;�=�]�=�m�=(* >�� >B�>�6>ǐ>�>)�>��>�\>t>��>�$>�� >�H >���=�X�=�	�=��=J"�=`��=� >�v >�� >.d>]�>QL>�   �   �>�A>�G>�%>�>KZ>K�>h� >���=0��=V�=n��=��=:��=L��=�=���=�$�=���=!�=���=��=���=��=>��=b��=n3�=�q�=>��=6� >�|>�>Џ>H�>b�>��>��>{}>�)>��>�m>l>� >� >Yq >8k >� >� >~� >L>p�>j>�{>��>�   �   ds>6�>6z>�C>X�>�N>n�>)� >�1�=���=tl�=R��="��=,=�=<:�=��=�R�=V��=�H�=l��=�I�=���=J)�=�'�=�f�=t��=�<�=|��=2��=�s >R>]>��>��>>�#>�>�>g�>T>�>8�>�{>�L>�1>p.>�B>�m>
�>h�>�O>��>�>NB>�   �   6�>��>��>Y>��>;E>3v>�| >���=�N�=��=$�=��=A�=�+�=�s�=^*�=�]�=P�=X�=  �=xd�=��=�'�=�{�=���=���=��=fc�=�C >�1>X�>.�>��>�4>CN>�G>�'>�>�>�t>R5>��>|�>m�>�>��>��>�3>Xy> �>H>�Y>f�>�   �   -�>��>��>�e>��>?>:f>Hc >�x�=���=bP�=��=��="��=���=x��=s�=���=�X�=,��=lh�=���=�o�=���=x��=�v�=��=��=��=d& >�>��>ˊ>��>�E>�g>.j>�R>�(>)�>��>�>6O>F+>>�>�+>xQ>��>��>+>ET>��>��>�   �   �,>&%>��>�z>��>G�>�� >�|�=�A�=���=��=�G�=���=�1�=�%�=��=���=z��=�=`z�=��=���=R�=�=x��=�7�=���=,��=�9�=0t�=Ԥ >t�>]�>�s>��>X>�(>�>��>��>>1>��>��>eQ>s)>�>e'>�M>��>W�>`,>A�>��>p>�   �   �>�>��>�v>��>��>�� >
��=Lf�=��=�<�=���=���=D~�=x�=���=��=���=�u�=F��=���=0��=&_�=f�=P��=�s�=/�=��=�\�=���=�� >��>b�>�o>k�>y>q>��>Q�>h>�>j�>�f>�'>u�>{�>5�>h#>Oa>]�>p	>�c>��>��>�   �   ��>%�>��> i>��>��>n� >~��=���=�n�=���=�<�=Բ�=�`�=�k�=(��=P�=T��=���=d��=2�=���=^N�=�C�=��=�%�=B��=X_�=���=t��=b� >t�>Y�>�b>��>��>A�>��>=j>>4�>`H>.�>'�>c>o>�|>�>�>c@>��>�>f>K�>�   �   �>��>k�>�Q>Z�>D >�� >i�=�}�=�E�=r��=�c�=���=4��= ��=���=>��=���=�D�=���=:��=�t�=��=̩�=���=�E�=,��=�0�=Tl�=�Y�=�� >��>��>�L>?�>��>Ό>CI>��>�{>�>�>h2>H� >�� >� >� >N� >�(>�>��>�q>�>�D>�   �   >>�M>�[>;0>��>M>I/>�	 >�b�=
d�=�2�=��=j��=^��= �=(��=��=���=t��=v��=���=���=��=8��=^��=b��=X�=*I�=�L�=]  >{'>�>��>->�Z>�O>w>F�>R=>��>�)>z� >�1 >��=�:�=��=*1�=Ĝ�=C% >� >�>T�>v1>��>�   �   �w>��>�
>�>e�>|7>�p>$o >Ru�=���=���=���=��="�=`|�=�_�=��=&��=g�=H��=l��=�4�=�J�=���=О�=��=���=���=T[�=�d >�h>�1>��>�>\>��>��>��>�f>H� >� >@��=d��=�=���=Xe�=j��=�=v��=���=� >w� >�V>�>�   �   5�>�N>��>J�>�>XU>P�>� >
��=l@�=��=t��=�,�=��=H�=:V�=���=z��=<��=|��=~��=�'�=��=N`�=���=��=Xu�=L�=&��=X� >��>ZP>��>=�>I�>.W>��>�+>4n >.M�=���=�U�=��=�+�=8��=\W�=���=�=���=�(�=(��="�=�Y >>�   �   �>P�>�<>y�>J�>�q>o>NW>3x >~��=Z��=h$�=L��=b�=PH�=���=n*�=�O�=V��=r=�=z�=lS�=*�=&'�="|�=���=e�=���=Qj >5M>��>6n>�>��>lC>,�>�>�@ >f��=���=&�=�m�=��=��=C�=z�=z2�=b��=R��=�:�=���=f��=N��=�, >�   �   1 >�>��>�F>D�>�>�K>��>t>OB >��=�r�=�N�=L?�=h_�=��=��=���=n��=���=�o�=*��=^(�=,�=~�=�?�=�b�="1 >�>��>�F>F�>�>�K>��>j>EB >΍�=tr�=�N�=?�=2_�=���=ޑ�=h��=6��=j��=�o�=���=*(�=��=N�=l?�=�b�=�   �   x��=Fj >,M>��>2n>�>��>rC>8�>�>�@ >���=��=R�=n�=�=:��=>C�=��=�2�=���=���=�:�=���=���=r��=�, >�>]�>�<>~�>M�>�q>j>HW>)x >h��=8��=B$�= ��=�a�=H�=L��=6*�=�O�="��=4=�=D�=<S�=��=�&�=�{�=f��=�d�=�   �   2�=��=N� >��>XP>��>?�>M�>7W>��>�+>En >RM�=���=V�=.�=
,�=n��=�W�=Ђ�=B�=���=)�=X��=N�=�Y >>C�>�N>��>L�>�>TU>L�>�� >���=P@�=��=P��=d,�=���=�G�=
V�=���=B��=��=F��=H��=X'�=��="`�=���=Ĳ�=8u�=�   �   h��=B[�=�d >�h>�1>��>�>_>��>��>��>�f>Z� >� >j��=���=>�=���=�e�=���=4�=���=���=� >�� >�V>�>�w>��>�
>�>d�>{7>�p>o ><u�=j��=���=`��=���=� �=.|�=�_�=���=���=�f�=��=<��=�4�=�J�=���=���=Н�=l��=�   �   I�=�L�=X  >t'>�>��>->�Z>�O>�>R�>`=>��>�)>�� >�1 >6��=�:�=��=P1�=��=T% >� >�>e�>�1>��>F>�M>�[>?0>��>L>D/>�	 >�b�=�c�=�2�=���=H��=:��=��=��=t�=R��=J��=D��=t��=X��=���=��=8��=D��=B�=�   �   �0�=Jl�=�Y�=�� >��>��>�L>?�>��>Ԍ>MI>��>�{>�>�>s2>X� >ͱ >� >'� >[� >�(>�>��>�q>�>�D>�>��>n�>�Q>[�>D >�� >
i�=�}�=�E�=^��=�c�=���=��=���=���=��=ʪ�=�D�=ڝ�=��=�t�=���=���=���=�E�=��=�   �   L_�=z��=l��=_� >q�>U�>�b>��>��>G�>��>Dj>>;�>hH>5�>0�>p>o>�|>��>�>j@>��>�>&f>Q�>��>(�>��>i>��>��>m� >r��=v��=zn�=���=�<�=Ʋ�=�`�=�k�=��=>�=<��=z��=L��=�=���=FN�=�C�=���=�%�=6��=�   �   ��=�\�=���=�� >��>c�>�o>k�>w>s>��>U�>h>�>o�>�f>�'>z�>��><�>n#>Ta>c�>x	>�c>��>��>�>�>��>�v>��>��>�� >��=Ff�=��=�<�=���=���=:~�=x�=���=��=���=�u�=<��=v��=.��=_�=�e�=D��=�s�=�.�=�   �   (��=�9�=,t�=Ҥ >r�>]�>�s>��>S>�(>�>��>��><1>��>��>eQ>t)>�>f'>�M>��>W�>_,>@�>��>q>�,>&%>��>�z>��>H�>�� >�|�=�A�=���=��=~G�=���=�1�=�%�=��=���=r��=�=Xz�=��=���=J�=�=j��=�7�=���=�   �   ��=�\�=���=�� >��>d�>�o>k�>w>t>��>U�>h>�>m�>�f>�'>y�>~�>:�>m#>Ta>d�>w	>�c>��>��>�>�>��>�v>��>��>�� >��=Pf�=��=�<�=���=���=L~�= x�=���=�=���=�u�=N��=���=>��=,_�=
f�=T��=�s�=/�=�   �   \_�=���=x��=c� >w�>Z�>c>��>��>C�>��>Bj>>:�>hH>4�>2�>m>o>�|>��>�>j@>��>�>!f>O�>��>)�>��>i>��>��>s� >���=���=�n�=���=�<�=��=�`�=�k�=>��=d�=b��=���=t��=@�=���=tN�=�C�=��=�%�=J��=�   �   �0�=bl�=�Y�=�� >��>��> M>@�>��>Ռ>KI>��>�{>�> �>s2>X� >ɱ >� >#� >X� >�(>�>��>�q>
�>�D>�>��>p�>�Q>`�>K >�� >i�=�}�=�E�=���=�c�=���=F��=��=Д�=T��=��=�D�=��=H��=�t�=��=ܩ�=���=�E�=:��=�   �   8I�=�L�=d  >'>�>��>->�Z>�O>�>P�>`=>��>�)>�� >�1 >0��=�:�=��=D1�=ޜ�=Q% >� >�>a�>1>��>E>N>�[>B0>��>T>M/>�	 >�b�=d�=�2�="��=���=x��=<�=J��=��=���=���=���=���=���="��=H��=n��=p��=h�=�   �   ���=j[�=�d >�h>�1>��>�>b>��>��>��>�f>T� >� >`��=���=6�=���=ze�=���=*�=���=���=� >�� >�V>�>�w>��>�
>�>l�>�7>�p>-o >hu�=���=��=���=:��=:�=z|�=�_�=8��=L��=8g�=n��=���=5�=K�=���=��= ��=���=�   �   `�=<��=^� >��>aP>��>C�>O�>8W>��>�+>Cn >JM�=���=V�=&�=,�=b��=�W�=�=6�=���=)�=N��=>�=�Y >>A�> O>�>R�>�>^U>X�>� >"��=�@�=&��=���=�,�=��=@H�=`V�=���=���=^��=���=���=�'�=�=f`�=��= ��=lu�=�   �   ���=]j >;M>��>;n>�>��>vC>6�>�>�@ >���=��=D�=�m�=��=0��=.C�=��=�2�=���=v��=�:�=���=���=l��=�, >�>^�>�<>��>T�>�q>x>ZW>?x >���=r��=�$�=h��=Bb�=vH�=���=�*�=P�=|��=�=�=��=�S�=R�=D'�=8|�=���="e�=�   �   ,1 >�>��>�F>O�>�>�K>��>t>PB >��=�r�=�N�=<?�=b_�=��=��=���=b��=���=�o�=��=T(�=�=n�=�?�=�b�= 1 >�>��>�F>O�>�>�K>��>�>[B >��=�r�=O�=n?�=�_�=D��=F��=���=���=ʺ�= p�=X��=�(�=H�=��=�?�=�b�=�   �   �>f�>�<>��>T�>�q>t>OW>4x >���=T��=b$�=<��=b�=HH�=v��=f*�=�O�=N��=\=�=p�=`S�=�='�=|�=���=e�=���=Rj >8M>��><n>�>��>~C>B�>�>�@ >���=<��=t�=,n�=,�=d��=fC�=��=�2�=���=���=�:�=��=���=���=�, >�   �   J�>O>	�>T�>�>\U>U�>� >��=h@�=��=t��=x,�=��=H�=2V�=���=h��=0��=r��=t��=�'�=��=F`�=���=��=Ru�=H�=(��=X� >��>aP>��>G�>V�>CW>��>�+>Qn >pM�=��=@V�=V�=0,�=���=�W�=��=h�=��=0)�=r��=d�=�Y >$>�   �   �w>��>�
>�>l�>�7>�p>&o >Ru�=~��=���=z��=��=�=V|�=�_�=��=��=
g�=B��=\��=�4�=�J�=���=Ğ�=��=���=���=X[�=�d >�h>�1>��>�>l>��>��>��>
g>d� >� >���=���=b�=ؗ�=�e�=���=V�=���=��= >�� >�V>�>�   �   P>N>�[>C0>��>Q>K/>�	 >�b�=d�=�2�=
��=b��=T��=�=&��=��=r��=f��=l��=���=v��=���=.��=P��=X��=R�=*I�=�L�=^  >|'>�>��>->�Z>�O>�>Z�>j=>��> *>�� >�1 >R��= ;�=��=n1�=��=b% >� >�>m�>�1>��>�   �   �>��>q�>�Q>_�>J >�� >i�=�}�=�E�=r��=�c�=���=,��=���=���=:��=��=�D�=���=.��=�t�=��=���=���=�E�=,��=�0�=Vl�=�Y�=�� >��>��>�L>F�>��>܌>RI>��>�{>�>�>�2>d� >ױ >-� >0� >h� >)>&�>��>�q>�>�D>�   �   ��>*�>��>i>��>��>o� >���=���=�n�=���=�<�=в�=�`�=�k�=.��=P�=N��=���=d��=*�=���=XN�=�C�=��=�%�=B��=T_�=���=t��=e� >x�>^�>c>��>��>I�>��>Jj>>C�>qH>>�>8�>v>o>�|>�>%�>t@>��>�>+f>T�>�   �   �>�>��>�v>��>��>�� >��=Lf�=��=�<�=���=���=D~�=x�=���=��=���=�u�=J��=���=6��=$_�=f�=R��=�s�= /�=��=�\�=���=�� >��>e�>�o>q�>}>t>��>U�>h>>t�>�f>�'>~�>��>@�>r#>Wa>j�>x	>�c>��>��>�   �   �r>�f>V>w>t�>>5>N"�=p:�=��=���=���=ވ�=�Y�=6r�=�
�=.Z�=X��='��=Z2�=<��=�w�=�<�=��=>\�=pP�=:��=n��=��=
�=L��=��=�n>c�>վ>Wd>+�>.�>;�>�N>;�>�f>�>wz>�>��>-�>��>��>�B>��>	>3�>��>�G>�   �   %Y> T>y
>�q>��>�<>�=�=b�=���=�-�=`�=>��=ҽ�=,��=j��=6��=��=�W�=λ�=J�=���=���=xc�=���=~��=B��=f,�=nW�=�9�=h��=��=�t>��>ݸ>�W>��>;�>�>m(>��>?6>��>�B>?�>��>��>��>)�>�
>�p>x�>~_>N�>�'>�   �   *>�>��>�a>��>/R>L��=V��=ȕ�=���=���=F��=x��=�(�=��=�S�=D��=���=vQ�=���=^��=4-�=��=��=d��=��=j�=��=X��=D�=���=��>k�>R�>2>�m>Uc>�!>��>�4>%�>>
�>17>�� >B� >�� >�>�d>��>�V>{�>�^>��>�   �   N�>��>�>eE>��>�s>� >���=h��=�=�c�=\��=���=�8�=l#�=>��=��=�t�=��=v`�=,��=���=���= �=ʖ�=o�=�Y�=�&�=��=2��=�* >�>�>��>r�>�>��>��>� >d>�>�> � > >���=�_�=�x�=J��=�V >u� >�m>E>է>�.>�   �   ��>�@>jU>X>4�>��>�Z >0��=���=���=hH�=���=�<�=H��=�=���=^e�=���=�E�=ּ�=�6�=ƞ�=���=���=��=҈�=�&�=���=���=ة�=qu >i�>x�>�U>��>�>�:>��>�	>�J>U� >4��=M�=LH�=z��=xP�=�o�=���=���=��=�4 >�� >u�>^>�   �   >��>��>t�>T�>d�>� >���=D^�=��=h��=a�=@8�="C�=���=f��=�[�=���=t[�=���=�"�=�\�=*U�=���=���=��=xT�=2u�=dN�=���=�� >2�>��>>�&>��>9f>=�>,� >���=��=�Y�=���=���=���=6��=P��=,\�=e�=��=m�=7�=T� >W]>�   �   O%>4�>[i>��>�{>=�>�(>���=��=���="�=xY�=���=t��=x��=���=���=�q�=���=�N�=$��=6��=~D�=|��=� �=���=��=|��=���=���=�,>>G�>d�>P�>�&>�m>8� >���=���=���=x��=���=��=ر�=�U�=���=�>�=�s�=��=�=� �=
O�=�4 >�   �   � >]>��>,L>qj>$.>��>f� >��=��=���=���=�#�=���=V��=br�=���=^I�=���=2"�=\;�=b�=^x�=�`�=t��=z�=�r�=���="��=i� >��>R3>�|>Mk>>qN> Z ><o�=P��=a�=l��=���=,��=��= �=t��=���=z��=j&�=F�=D�=���=xT�=��=�   �   ���=J9 >|:>��>R>�X>�>M[>Mf >�h�=x��=6��=���=���=�L�=��=$W�=�9�=��=��=�=H��=���=�X�=4�=x2�=�+�=���=Y9 >�:>��>R>�X>�>B[>>f >�h�=H��=���=���=>��=�L�=��=�V�=d9�=���=z�=��= ��=X��=XX�=�3�=F2�=�+�=�   �   ~��= ��=_� >��>N3>�|>Tk>�>�N>1Z >jo�=���=Va�=���=��=p��=:�=p�=į�=*��=���=�&�=��=LD�=���=�T�=<��=� >m>�>3L>uj>$.>��>[� >���=��=V��=j��=�#�=���=��=r�=\��=I�=���=�!�=;�=�=x�=�`�=8��=H�=xr�=�   �   V��=���=���=�,>>G�>i�>X�>�&>n>O� >���=���=ܢ�=���=���=\��=&��=6V�=L��=�>�=�s�=��=L�=� �=:O�=�4 >b%>A�>bi>�>�{>:�>�(>���=��=���=�!�=DY�=���=4��=0��=n��=^��=�q�=r��=�N�=؉�=���=:D�=<��=� �=���=���=�   �   u�=LN�=l��=�� >/�>��>>�&>�>If>R�>F� >��=��=�Y�=
��=:��=��=v��=���=l\�=Ve�=@��=>m�=J7�=j� >j]>>��>��>y�>V�>b�>�� >���=$^�=��=@��=�`�=8�=�B�=p��="��=�[�=���=,[�=���=�"�=d\�=�T�=���=N��=`�=RT�=�   �   ���=���=ȩ�=lu >f�>z�>�U>��>&�>�:>��>�	>�J>i� >l��=6M�=�H�=���=�P�=p�=���=��=��=�4 >�� >��>%^>��>�@>qU>[>4�>��>{Z >��=j��=���=BH�=���=�<�=��=��=���=e�=���=bE�=���=V6�=���=���=P��=���=���=x&�=�   �   �&�=��="��=�* >�>�>��>r�>�>��>��>� >/d>��>�>2� >% >Ƣ�=�_�=y�=t��=�V >�� >�m>U>�>�.>Z�>��>�>fE>��>�s>� >���=T��=�=�c�=6��=���=�8�=@#�=��=f�=Xt�=���=D`�=���=h��=j��=��=���=�n�=�Y�=�   �   r�=N��=:�=���=��>h�>S�>2>�m>Zc>�!>��>�4>0�>+>�>B7>� >P� >�� >�>�d>��>�V>��>�^>��>2>�>��>�a>��>/R>L��=L��=���=���=���=*��=b��=�(�=���=�S�="��=���=XQ�=���=<��=-�= ��=~�=D��=���=X�=�   �   dW�=�9�=^��=��=�t>��>ܸ>�W>��>>�>��>v(>��>B6>��>�B>G�>��>��>��>2�>�
>�p>��>�_>V�>�'>+Y>T>{
>�q>��>�<>�=�=b�=���=�-�=R�=0��=Ľ�=��=Z��="��=��=�W�=���=�I�=���=~��=hc�=z��=f��=6��=X,�=�   �   ��=
�=N��=���=�n>a�>Ӿ>Vd>)�>/�><�>�N>9�>�f>�>wz>�>��>-�>��>��>�B>��>
>4�>��>�G>�r>�f>Z>w>s�><5>R"�=p:�=��=���=���=ڈ�=�Y�=8r�=�
�=.Z�=S��='��=X2�=7��=�w�=�<�=��=:\�=hP�=6��=n��=�   �   pW�=�9�=h��="��=�t>��>�>�W>��>=�>�>p(>��>F6>��>�B>F�>��>��>��>/�>�
>�p>�>�_>T�>�'>*Y>T>}
>�q>��>�<>�=�= b�=��=�-�=f�=B��=ֽ�=6��=t��=>��=��=�W�=ֻ�=J�=���=���=�c�=���=���=J��=j,�=�   �   ��=d��=H�=���=��>l�>U�>2>�m>\c>�!>��>�4>,�>(>�>A7>� >O� >�� >�>�d>��>�V>��>�^>��>1>�>��>�a>��>6R>Z��=b��=ҕ�=���=���=R��=���=�(�=��= T�=`��=��=�Q�=���=t��=J-�=2��=��=p��=��=v�=�   �   �&�=(��=>��= + >�> �>��>s�>�>��>��>� >+d>��>�>.� ># >���=�_�=y�=n��=�V >�� >�m>S>�>�.>Z�>��> �>lE>��>�s>� >���=|��=.�=�c�=p��=��=�8�=�#�=\��=��=�t�=$��=�`�=F��=���=���=6�=ܖ�=(o�=�Y�=�   �   Υ�=���=��=xu >o�>��>�U>��>&�>�:>��>�	>�J>d� >`��=0M�=xH�=���=�P�=p�=���=��=��=�4 >�� >��>$^>��>�@>uU>`>?�>��>�Z >H��=���=²�=�H�=ܼ�=�<�=r��=4�=*��=�e�=���=�E�=���=�6�=��=��=���=*��=��=�&�=�   �   Hu�=|N�=���= � >8�>ƭ>>�&>�>Ff>Q�>A� >��=��=�Y�=��=.��=��=h��=���=\\�=Je�=6��=,m�=>7�=e� >i]>>��>��>�>]�>q�>� >���=\^�=.��=���=6a�=f8�=JC�=ޯ�=���= \�=,��=�[�=��=#�=�\�=TU�=���=���=��=�T�=�   �   ���=���=���=�,>>N�>p�>\�>�&>n>K� >���=���=΢�=���=���=P��=��=&V�=:��=�>�=�s�=��=>�=� �=4O�=�4 >a%>C�>hi>�>|>I�>�(>���=��=���=6"�=�Y�=���=���=���=���=���=r�=���=O�=Z��=j��=�D�=���=� �=���=(��=�   �   ���=@��=s� >��>\3>�|>Yk>�>�N>/Z >bo�=z��=Da�=���=ғ�=d��=,�=^�=���=��=���=�&�=|�=<D�=��=�T�=8��=� >p>�>:L>�j>2.>��>v� >:��=��=���=ʄ�=$�=��=���=�r�=��=�I�=$��=l"�=�;�=��=�x�=*a�=���=��=�r�=�   �   ��=f9 >�:>��>R>�X>�>N[>Kf >�h�=n��=,��=���=p��=�L�=��=W�=�9�=���=��=��=<��=���=�X�=4�=l2�=�+�=���=Y9 >�:>��>R>�X>�>][>^f >i�=���=`��=���=���=M�=�=hW�=�9�=>��=�=>�=���=���=�X�=B4�=�2�=,�=�   �   � >{>�><L>�j>/.>��>g� >��=��=|��=���=�#�=���=L��=Xr�=���=FI�=���="�=J;�=X�=Nx�=�`�=d��=n�=�r�=���=&��=l� >��>\3>�|>bk>�>�N>BZ >�o�=���=�a�=���=��=���=v�=��=���=`��=���=�&�=��=vD�=��=�T�=\��=�   �   o%>O�>oi>�>|>E�>�(>���=��=���="�=tY�=���=d��=h��=���=���=�q�=���=�N�=��=(��=lD�=l��=� �=���=��=x��=���=���=�,>>R�>u�>f�>�&>n>c� >��=���=
��=��=��=���=Z��=jV�=~��=$?�=2t�=�=t�=� �=XO�=�4 >�   �   )>��>��>��>_�>k�>� >���=D^�=��=\��=a�=28�=C�=���=V��=�[�=���=b[�=���=�"�=�\�=U�=���=v��=��=pT�=0u�=hN�=���=�� >:�>ŭ>>�&>�>Yf>c�>S� >D��=��=Z�=:��=r��=J��=���=¾�=�\�=�e�=r��=`m�=f7�=w� >y]>�   �   ��>�@>yU>b>;�>��>�Z >6��=���=���=^H�=���=�<�=<��=�=���=Pe�=���=�E�=ļ�=�6�=���=���=x��=��=ƈ�=�&�=���=���=ܩ�=vu >p�>��>�U>�>2�>�:>��>�	>�J>}� >���=bM�=�H�=��=�P�=8p�="��=@��=�=�4 >�� >��>.^>�   �   b�>��>'�>lE>��>�s>� >���=l��=�=�c�=P��=���=�8�=b#�=2��=��=~t�=���=l`�=��=���=���=�=�=o�=�Y�=�&�=��=8��=�* >�>"�>��>|�>�>��>��>� ><d>�>�>C� >6 >��=`�=.y�=���=�V >�� >�m>a>�>�.>�   �   3>�>��>�a>��>2R>R��=Z��=ƕ�=���=���=@��=p��=�(�=��=�S�=@��=���=vQ�=���=X��=0-�=��=��=\��=���=f�=��=X��=H�=���=��>o�>Y�>"2>�m>ac>�!>��>5>=�>5>!�>K7>� >^� >�� >�>�d>��>�V>��>�^>��>�   �   +Y>T>}
>�q>��>�<>�=�=b�=���=�-�=\�=<��=ʽ�=*��=j��=2��=��=�W�=Ȼ�= J�=���=���=vc�=���=x��=>��=`,�=pW�=�9�=l��="��=�t>��>�>�W>��>A�>�>x(>��>I6>��>�B>L�>ã>��>��>5�>�
>�p>��>�_>X�>�'>�   �   ��>З>�'>!K>L�>
/ ><��=N��=�h�=���=Dj�=���=�x�=#Y�=���=�p�=K�=���=Ƹ=K��=U,�=L�=��=�D�=z�=(�=P��=��=Z��=*�=l��=�� >�w>��>w�>�7>aO>>>��>D
>�_>��>z>��>@>�>�>�S>��>�8>�>;m>��>xo>�   �    �>i}>�>�C>��>m: > �=���=���=�=���=pn�=�
�=6��=ږ�=�/�=�=�|�=���=�i�=t�=��=p�=���=v�=��=��=�Z�=.�=D\�=v��=b� >�w>j�>�>�>�*>N�>�n>v�>M>�l>��>�H>�� >�� >v� >�>�h>��>Ӎ>�1>:�>=C>�   �   �>M/>��>�->\>�Z >�z�=xd�=���=J�=��=���=���=��=���=�a�=@_�=�ؼ=���=���=�5�=�,�=�m�=��=ޟ�=:��==�=�S�=h��=��=�'�=]� >)w>ı>�t>��>y�> e>h�>�>NX>�>�� >�[ >���=ښ�=���=A >�� >�>��>��>K/>b�>�   �   r>�>ޑ>>�>y� >�2�=zn�=
��=(��=�!�=�D�=\k�=(��=���=Q��=�=���=$ſ=P��=���=���=K��=^��=5�=�'�=�#�=���=f1�=N��=\��=.� >�r>��>�>�C>B>i�>��>3�>�>�; >"��=P��=F��=�|�=
��=r(�=�'�=t~�=
� >�`>d3>��>�   �   �>�>a>��>Y>�� >�!�=`��=D��=���= ��=�i�=L �=���=�J�=��=���=ڦ�=���=���=e��=64�=]��=�u�=��=8%�=��=*��=���=$�=ґ�=�>@h>s>>}�>I�>�>�g>E|>u >���=���=�=:��=Ȳ�=�G�=j�=��=TC�=���=���=D��=� >��>�   �   `n>R+>��>�>9	>�>&8�=�m�=p��=��=f�=�,�=�H�=���=�}�=S�=���=��=���=�s�=Co�=��=���=$�=��=>��=`��=�=���=�=��=�G>�T>�>��>ũ>��>b >گ�=�0�=4��=�V�=jJ�=��=H��=z"�=zP�=| �=���=�a�=��=l	�=���=�m >�   �   Y$ >/>�>w+>��>�V>�3 >�;�=�G�=P��=x��=b`�=��=^��=�E�=L�=�<�=�E�=ʇ�=��=X��=���=2��=XA�=c�=��=>(�=�R�=��=,�=A >dy>�6>4w>�@>��>0� >���=z��=���=t��=P4�=���=b��=̹�=�5�=r�=k�=��=bE�=Z��=@��=��=���=�   �   @o�=� >�>��>C�>�>�� >��=T��=,��=�}�=h��=��=,��=._�=(��=P�=<G�=
��=�
�=D��=�/�=t��=<��=bJ�=$�=v��=�V�=Ll�=���=�� >�>%>��>�j>t >�K�=�,�=`��=$5�=��=���=���=���=�?�=��=<��="�=��=^��=��=�,�=���=�7�=�   �   *j�=j��=�K >�F>��>��>h>� >�g�=�!�=t`�=�V�=x7�=B7�=z��=Xd�=���=�[�=d��=�=�t�=v��="��=�M�=�G�=�n�=V��=bj�=���=�K >G>��>��>h>�� >�g�=�!�=0`�=PV�="7�=�6�=��=�c�=J��=N[�=��=��=jt�=��=���=PM�=�G�=~n�=��=�   �   fV�=$l�=���=�� >�>%>��>�j>*t >�K�=-�=���=r5�=@��=��=���= ��=(@�=~��=���=�"�=:�=���=r��= -�=Ⱥ�=�7�=po�= >�>��>G�>�>{� >��=*��=���=Z}�=��=f�=֊�=�^�=���=��=�F�=���=`
�=Ԛ�=6/�=��=��=J�=��=<��=�   �   �R�=��=�+�=A >`y>�6><w>�@>ɞ>I� >.��=���=<��=���=�4�=R��=���=8��=6�=pr�=zk�=,�=�E�=���=���=F��=���=q$ >&/>"�>+>��>�V>�3 >�;�=�G�=��=:��=`�=T�= ��=,E�=�K�=J<�=wE�=Z��=�=���=`��=Р�= A�=�b�=���=(�=�   �   �~�=���=���=��=�G>�T>�>��>ԩ>�>} >��=1�=���=�V�=�J�=<��=���=�"�=�P�=� �=��="b�=P��=�	�=ȃ�=�m >tn>`+>��>�>8	>�>8�=�m�=F��=��=.�=�,�=@H�=���=x}�=��=z��=���=H��=ws�=�n�=���=x��=��=���=���=*��=�   �    ��=|��=�=���=>?h>z>>��>S�>�>�g>a|>)u >���=���=^�=���=��=�G�=Zj�=��=�C�=��=<��=���=$� >��>�>�>g>��>Y>�� >�!�=H��=$��=���=���=Xi�=
 �=8��=�J�=���=i��=p��=p��=b��=��=�3�=��=Pu�=ؤ�=�$�=���=�   �   ���=P1�=:��=N��='� >�r>��>�>�C>N>{�>��>H�>�>�; >V��=���=���=�|�=N��=�(�=�'�=�~�=$� >�`>w3>��>"r>�>�>>�>w� >�2�=hn�=���=��=�!�=�D�=$k�=���=l��=��=��=W��=�Ŀ=��=���=l��=
��=!��=�4�=�'�=�#�=�   �   �S�=X��=���=�'�=[� >&w>Ʊ>�t>��>��>(e>u�>�>]X>�>� >�[ >���=��=(��=W >�� >�>�>��>Z/>k�>�>V/>��> .>X>�Z >�z�=nd�=x��=4�=t�=���=f��=���=���=fa�=_�=pؼ=���=`��=^5�=�,�=�m�=ů�=���=��=�<�=�   �   �Z�=.�=<\�=p��=_� >�w>m�>�>�>�*>T�>�n>|�>U>�l>��>�H>� >�� >�� >�>�h>��>ۍ>�1>B�>GC>)�>o}>�>�C>��>m: >��=���=��=�=���=\n�=�
�=��=���=�/�=��=�|�=���=�i�=T�=��=�o�=g��=^�=Ԅ�=��=�   �   |�=\��=�)�=h��=�� >�w>��>w�>�7>bO>=>��>D
>�_>��>z>��>@>�>�>�S>��>�8>�>:m>��>{o>��>ӗ>�'>!K>M�>	/ >@��=L��=�h�=���=@j�=���=�x�=#Y�=���=�p�=K�=���=Ƹ=G��=T,�=L�=��=�D�=z�= �=T��=�   �   �Z�=.�=D\�=z��=b� >�w>m�>�>�>�*>T�>�n>|�>T>�l>��>�H>� >�� >� >�>�h>��>ڍ>�1>B�>EC>(�>o}>�>�C>��>q: >�=���=���= �=���=xn�=
�=E��=��=�/�=�=�|�=���=�i�=|�=�=p�=���=z�=��=��=�   �   �S�=x��=��=�'�=c� >,w>ɱ>�t>��>�>)e>u�>�>XX>�>� >�[ >���=���= ��=U >�� >�>�>��>V/>n�>>W/>��>.>`>�Z >�z�=�d�=���=Z�=��=��=���=-��=ң�=�a�=h_�=�ؼ=���=���=�5�=-�=n�=��=��=H��==�=�   �   ���=�1�=\��=l��=6� >�r>��>�>�C>M>y�>��>F�>�>�; >N��=���=|��=�|�=@��=�(�=�'�=�~�=� >�`>v3>��>#r>�>�>!>�>�� >�2�=�n�= ��=@��=�!�=
E�=�k�=V��=���=���=H�=ޢ�=Vſ=���=��=��=x��=~��=,5�=�'�=$�=�   �   H��=���=<�=��=�>Kh>~>>��>W�>�>�g>\|>%u >���=���=T�=x��=
��=�G�=Hj�=��=�C�=��=6��=t��=� >��>�>�>m>��>g>�� >�!�=~��=f��=���=$��=�i�=| �=���=K�="��=��=��=��=���=���=w4�=���=�u�=F��=X%�=��=�   �    �= ��=܌�=��=�G>�T>�>��>ש>�>y >��=1�=n��=�V�=�J�=.��=���=�"�=�P�=� �=���=b�=@��=�	�=���=�m >un>e+>��>�>H	>�>F8�=n�=���=<��=��=-�=�H�=6��=~�=��=(��=`��=��=+t�=�o�=&��=��=^�=H��=d��=���=�   �   �R�=��=8,�=A >py>�6>Fw>�@>ɞ>I� >&��=���=(��=���=�4�=B��=���="��=�5�=Vr�=fk�=�=�E�=���=~��=>��=���=q$ >)/>+�>�+>�>�V>�3 >�;�=�G�=z��=���=�`�=��=���=�E�=lL�==�==F�=��=��=���=��=z��=�A�=Pc�=.��=h(�=�   �   �V�=tl�=��=�� > �>4>�>�j>)t >�K�=-�=���=^5�=0��=��=���=��=@�=h��=���=h"�=$�=���=Z��=-�=���=�7�=po�= >>ɿ>V�> �>�� >��=���=^��=�}�=���=��=x��=�_�=~��=��=�G�=d��=*�=���=�/�=���=z��=�J�=V�=���=�   �   �j�=���=�K >G>��>��>h>� >�g�=�!�=j`�=�V�=d7�=07�=h��=Dd�=���=�[�=N��=��=�t�=`��=��=�M�=�G�=�n�=H��=\j�=���=�K >G>��>��>h>� >h�= "�=�`�=�V�=�7�=�7�=ʊ�=�d�=��=\�=���=h�=.u�=ȴ�=p��=�M�=H�=�n�=���=�   �   �o�=" >>Ϳ>V�>�>�� >��=T��=*��=�}�=\��=��=��=_�=��=<�= G�=���=�
�=.��=�/�=\��=&��=NJ�=�=t��=�V�=Rl�=���=�� > �>7>�>�j>@t >�K�=B-�=��=�5�=���=P��=@��=r��=z@�=Э�= ��=�"�=��=
��=���=T-�=���=�7�=�   �   �$ >8/>4�>�+>�>�V>�3 >�;�=�G�=J��=p��=X`�=��=H��=�E�=L�=�<�=�E�=���=x�=B��=���=��=BA�=c�=���=4(�=�R�=��=$,�=A >oy>�6>Nw>�@>ޞ>^� >^��=���=t��=��=�4�=���=��=���=P6�=�r�=�k�=x�=�E�=���=���=r��=��=�   �   �n>r+>��>�>G	>�>28�=�m�=p��=��=Z�=�,�=xH�=��=�}�=?�=���=���=���=�s�=)o�=˪�=���=�=��=.��=V��=�~�= ��=Č�=��=�G>�T>"�>��>�>#�>� >H��=P1�=���=<W�=�J�=���=��=#�=Q�=!�=J��=bb�=���=�	�=���=�m >�   �   ,�>�>u>��>g>�� >�!�=d��=F��=���=���=�i�=< �=r��=�J�=Ԑ�=���=���=���=���=S��=&4�=O��=�u�=
��=(%�=ܬ�=$��=���=*�=ޑ�=�>Lh>�>>��>e�>�>�g>v|>Au >���=��=��=���=V��=8H�=�j�=(�=�C�=\��=l��=���=3� >�>�   �   -r>'�>�>#>�>� >�2�=~n�=��=&��=�!�=�D�=Pk�=��=���=G��=�=���=ſ=>��=���=���=7��=P��=�4�=�'�=�#�=���=h1�=R��=f��=6� >�r>��>>�C>[>��>��>[�>�>�; >���=���=���=
}�=v��=�(�=�'�=�~�=4� >�`>�3>��>�   �   >]/>��>.>`>�Z >�z�=~d�=���=H�=��=���=~��=
��=���=�a�=6_�=�ؼ=���=���=�5�=�,�=�m�=��=֟�=4��=�<�=�S�=d��=��=�'�=d� >0w>α>�t>��>��>4e>��>�>iX>-�>� >�[ >���=(��=F��=f >�� >�>�>��>c/>u�>�   �   *�>q}>�>�C>��>n: > �=���=���=�=���=ln�=�
�=.��=Ԗ�=�/�=��=�|�=���=�i�=j�=��=p�=u��=p�=���=��=�Z�=.�=F\�=z��=f� >�w>o�>��>�>�*>Z�>�n>��>_>�l>��>�H>
� >�� >�� >�>�h>��>�>�1>C�>IC>�   �   G�>�>H>��>O>�D�=� �=l��=L8�=���=k[�=6��=S��=�>�=���=0��=�P�=6d�=��=�M�=�)�=?^�=n��=Q/�=/Ƚ=���=���=>I�= �=$��=bF�=|��=��>��>2�> �>V�>x]>F�>��>>� >uN>� >y, >���= ��=�A >u� >cp>p;>�>l�>9l>�   �   V�>�{>��>F�>�>>d�=TY�=p�=��=*1�=^��=M�=*��=o0�=���=$��=�="��=�>�=q��=�S�=w�=���=��=딾=6~�=xZ�=d��=�c�=
�=Lv�=���=��>��>2�>�`>�v>� >z>��>e�>��>C� >97 >b{�=\�=P�=`��=�Z >)>��>+�>�>�0>�   �   �>�>z�>ձ>�>���=���=���=���=���=���=�r�=��=���=tǭ=���=x��=x-�=�ך=|�=ƿ�=���=���=�ö=T��=T��=|�=�'�=�}�=���=��=���=Y�>�q>E{>R�>��>�l>��>��>��>�� >fk�=���=���=�q�=���=�+�=Q�=���=� >��>��>�>�   �   �>d>9>s}>#>:G�=0��=x�=|��=T"�=���=���=0��=�i�=0��=~;�=���=��=噠=��=�9�=�ڪ=�F�=��=9��=���=~��=�f�=xB�=(#�=���=>S�=y�>�.>��>�8>Z�>qF>�M>|(>&��=��=Ɔ�=��=T��=B;�=�Y�= �=@j�=3�=P�=�J >�g>�_>�   �   �>�x>�>3>)>D��=�J�=�d�=�Z�=8X�=B��=�p�=@2�=iG�= �=�+�=.Ҭ=�i�=�-�=05�=$p�=r��=쎸=���=ո�=��=�p�=�`�=���=���=���=���=��>~�>�Q>?>�>��>�{ >b.�=T�=\��=�;�=�V�=��=�|�=Χ�=���=0�=�;�=H��=�z�=,7�=�� >�   �   ,X >�U>I�>C�>,(>���=B��=T��=�d�=6*�=8�=���=f�=3<�=���=�`�=Vu�=(O�=7%�=��=���=Q��=��=�x�=���=.B�=���=��=2`�=���=8�=i+ ><�>7X>]z>]
>,>��=L�=0�=��=^z�=ح�=�w�= ��=�Y�=���=Į�=B��=��=�!�=�q�=���=���=�   �   7�=S >�� >X> >�; >j�=#�=���=�d�=U�=���=�B�=���=�/�=�m�=d��=Z�=H�=Tл=�h�=D��= F�=��=R�=V �=L��=���=�s�=.�=4��=�n >�l>��>{>� >���=�8�=�T�=�6�="�= U�=��=�q�=p��=��=fT�=���=<��=���=X��=���=���=��=�   �   _�=��=Z��=v� >>ՙ >��=ȵ�=�=�=���=���=%�=�u�=b��=9�=^��=���=]�=_�=*�=;H�=���=���=��=�N�=��=(��=J�=���=�`�= ��=� >_5>a>�Z >��=���=�U�=ƚ�=
��=l��=�`�=��=��=$��=��=� �=ؿ�=�v�=�=�o�=�5�=&'�=���=�   �   :F�=l��=���=8) >� >o� >W >�C�=D��=�H�=t�=*z�=���=��=r��=T_�=���=f��=��=�A�=�/�=
c�=ƨ�=���=:\�=�1�=v��=�F�=���=���=B) >� >k� >�V >�C�=��=�H�=�=�y�=~��=(�=���=�^�=��=���=b��=
A�=�.�=rb�=:��=���=�[�=1�=��=�   �   �=Į�=�`�=��=� >a5>m>�Z >��=���=V�=.��=x��=���=Pa�=���=t��=ȅ�=���=�!�=p��=|w�=��=p�=H6�=�'�=@��=N_�=�=|��=�� >>Й >��=���=�=�=���=8��=�$�=Bu�=���=� �=���=��=p\�=d^�=z�=�G�=���=K��=���=ZN�=>�=���=�   �   ���=�s�=�=��=�n >�l>��>{>� >ҝ�=9�=FU�=T7�=�"�=�U�=<	�=zr�=��= �=�T�=��=���=j��=΢�=���=���=.��=N7�=j >�� >X>>�; >�i�=�"�=���=�d�=�T�=X��=xB�=��=Y/�=	m�=���=��=��=�ϻ=(h�=���=uE�=���=�Q�=���=���=�   �   ���=�_�=���=�7�=b+ ><�>AX>lz>p
>F>L��=��=��=p��=�z�=H��=bx�=���= Z�=v��=>��=���=�=&"�=r�="��=���=GX >�U>X�>H�>)(>���=*��=,��=Ld�=�)�=�7�=���=�e�=�;�=j��=V`�=�t�=�N�=�$�=P�=<��=ú�=�=ex�=��=�A�=8��=�   �   t`�=���=���=���=���=��>��>�Q>(?>3�>ϸ>�{ >�.�=`T�=���=P<�=W�=�="}�=:��=&��=��="<�=���=�z�=p7�=�� >0�>�x>��>3>)>6��=�J�=td�=ZZ�=�W�=���=kp�=�1�=�F�=��=+�=�Ѭ=Fi�=6-�=�4�=�o�=�={��=��=v��=s�=�p�=�   �   Rf�=RB�=
#�=���=6S�=v�>/>��>�8>j�>�F>N>�(>`��=b��=��=R��=���=�;�=Z�=N�=�j�=b3�=LP�=�J >�g>�_>�>d>9>v}>#>4G�= ��=�w�=Z��=$"�=n��=���=���=`i�=Ь�=;�=N��=E�=r��=���=�9�=rڪ=#F�=��=��=���=L��=�   �   �'�=�}�=���=��=���=V�>�q>I{>X�>��>�l>��>��>��>ٟ >�k�=���=���=�q�=܇�=,�=HQ�=���=/� >�>��>�>�>�>}�>ر>�>���=v��=���=���=���=���=Zr�=Q�=���=)ǭ=f��=/��=-�=�ך=$�=y��=P��=p��=�ö=��=#��=X�=�   �   T��=�c�=�=Dv�=��=��>��>4�>�`>�v>� >!z>��>q�>��>O� >F7 >�{�=~�=p�=|��=[ >5>��>8�>��>�0>`�>�{>��>G�>�><d�=PY�=d�=Ρ�=1�=B��=�L�=��=M0�=x��=���=�~�==�>�=F��=�S�=�v�=���=��=˔�=~�=hZ�=�   �   :I�= �= ��=^F�=x��=��>��>0�>��>S�>x]>G�>��>>� >tN>� >{, >���=��=�A >x� >dp>t;>�>o�><l>J�>�>G>��>N>�D�=� �=l��=F8�=���=d[�=,��=Q��=�>�=v��=!��=�P�=0d�=��=�M�=�)�=6^�=m��=Q/�='Ƚ=���=���=�   �   p��=�c�=�=Tv�= ��=��>��>5�>�`>�v>� >!z>��>n�>��>N� >E7 >|{�=v�=j�=z��=[ >3>��>4�>��>�0>a�>�{>��>O�>�>Fd�=bY�=|�=��=61�=j��=M�=<��=�0�=���=:��=(�=7��=�>�=���=�S�=w�=ċ�=��=���=F~�=�Z�=�   �   �'�=�}�=���=��=���=^�>�q>N{>Z�>��>�l>��>��>��>؟ >�k�=���=���=�q�=҇�=,�=BQ�=���=)� >�>��>�>�>�>��>�>�>ƽ�=���=��=���=Դ�=��=�r�=��=��=�ǭ=���=���=�-�=ؚ=��=���=ɰ�=ރ�=Ķ=r��=j��=��=�   �   �f�=�B�=<#�=��=VS�=��>/>��>�8>l�>�F>N>�(>V��=T��=��=J��=���=�;�=�Y�=B�=�j�=V3�=BP�=�J >�g>�_>�>d>!9>�}>#>VG�=L��= x�=���=z"�=ػ�=-��=j��=�i�={��=�;�=��=�=7��=T��=B:�=$۪=�F�=�=l��=���=���=�   �   �`�=Ҙ�=���=��=���=�>��>�Q>/?>.�>ɸ>�{ >�.�=LT�=���=F<�=�V�=��=}�=$��=��=��=<�=���=�z�=d7�=�� >2�>�x>�> 3>)>d��=K�=�d�=�Z�=dX�=z��=q�=�2�=�G�=n �=�+�=�Ҭ=<j�=%.�=�5�=�p�=ѩ�=A��=ι�=��=��= q�=�   �   B��=^`�=���="8�=y+ >M�>LX>rz>v
>G>B��=��=x�=\��=�z�=6��=Nx�=l��=Z�=`��=(��=���=��="�=r�=��=���=GX >V>]�>V�>@(>��=l��=���=�d�=l*�=J8�=4��=`f�=�<�=X��=Xa�=�u�=�O�=�%�=b�=?��=���=��=2y�=Ӱ�=lB�=���=�   �   4��=t�=X�=Z��=�n >�l>�> {>� >Н�=
9�=8U�=>7�=t"�=hU�=&	�=dr�=��=�=�T�= ��=���=T��=���=ޢ�=��=$��=J7�=n >�� >$X>>�; >@j�=@#�=.��=*e�=ZU�=��=LC�=���=W0�=n�=���=��=��=�л=:i�=���=oF�=e��=RR�=� �=���=�   �   ��=4��=a�=J��=� >v5>w>�Z >��=ؗ�=V�= ��=`��=���=<a�=p��=V��=���=n��=p!�=P��=^w�=n�= p�=46�=z'�=<��=L_�=�=���=�� >>� >��=���=$>�=��=޴�=`%�=v�=���=��=���=D��=�]�=�_�=��=�H�= �=P��=p��=&O�=��=n��=�   �   �F�=���=��=W) >)� >�� >W >�C�=J��=�H�=d�=z�=��=��=Z��=8_�=���=F��=��=�A�=o/�=�b�=���=h��=\�=l1�=j��=~F�=���=Ĭ�=P) >&� >�� >#W >D�=���= I�=��=�z�=T��=�=���=�_�=*��=��=���=/B�=0�=�c�=:��=��=�\�=�1�=���=�   �   �_�=B�=���=�� >>� >��=е�=�=�=���=���=�$�=�u�=J��=�=D��=���=�\�=�^�=�=H�=i��=���=���=�N�=��= ��=D�= ��=�`�=4��= � >y5>�>�Z >.�=��=dV�=~��=ԯ�=N��=�a�=���=���=>��=��="�=���=�w�=��=tp�=�6�=�'�=���=�   �   �7�=� >�� >*X>>�; >(j�=#�=���=�d�=U�=���=�B�=p��=�/�=�m�=H��=<�=&�=2л=�h�=(��=�E�=���=�Q�=B �=@��=���=�s�=8�=J��=�n >�l>�>2{> � >
��=V9�=�U�=�7�=�"�=�U�=�	�=�r�=p��=��=hU�=���=,��=���= ��=D��=<��=l��=�   �   `X >V>j�>\�>>(>ֲ�=L��=X��=�d�=4*�=�7�=���=�e�=<�=���=�`�=?u�=O�=%�=��=���=3��=n�=�x�=m��=B�=t��=��=0`�=���=8�=y+ >P�>UX>�z>�
>b>���=��=��=���=&{�=���=�x�=���=�Z�=Ԗ�=���=��=`�=v"�=`r�=`��=,��=�   �   F�>�x>
�>!3>)>R��=�J�=�d�=�Z�=2X�=8��=�p�=-2�=QG�= �=x+�=Ҭ=�i�=�-�=5�=p�=Z��=Ԏ�=n��=���=��=�p�=�`�=���=���=��=���=
�>��>�Q>C?>F�>�>| >�.�=�T�=��=�<�=fW�=X�=t}�=���=x��=��=l<�=޿�={�=�7�=�� >�   �   
>'d>,9>�}>#>LG�=8��=x�=���=N"�=���=���="��=�i�=!��=n;�=���=��=͙�=�=�9�=�ڪ=lF�=��=*��=���=x��=zf�=vB�=,#�=���=TS�=��>/>��>�8>~�>�F>+N>�(>���=���=P��=���=���=�;�=DZ�=��=�j�=�3�=xP�=K >�g>�_>�   �    �>�>��>�>�>���=���=���=���=���=���=�r�=��=���=fǭ=���=p��=d-�=�ך=j�=���=���=���=�ö=H��=J��=v�=�'�=�}�=���=��=���=b�>�q>X{>g�>��>�l>ͦ>��>ʤ>� >�k�=��= ��=r�=��=D,�=rQ�=��==� >#�>��>�>�   �   f�>�{>��>M�>�>Bd�=ZY�=n�=��=,1�=\��=M�=$��=k0�=���=��=�=��=�>�=o��=�S�=�v�=���=��=䔾=4~�=tZ�=f��=�c�=�=Pv�=���=��>��>:�>�`>�v>� >+z>��>z�>��>\� >R7 >�{�=��=��=���=[ >A>��>>�> �>�0>�   �   d�>�b>v�>_>�D�=���=�B�=\��=��=�Z�=��=}Э= ��=�_�=��=��g=p�T=�H=��D="�H=V�T=�Pg=��=�[�=�=u7�=�&�=�B�=>�=�\�=���=�{�=� >�>y�>o�>��>�^>&�>?|>SF>N>d��=�6�=^��=~h�=F{�=�5�=l��=�) >~8>�S>VY>�!>�   �   �F>F3>Tw>��>�I�=P��=��=dn�=P��=��=�g�=��=n�=�ȏ=r��=�k=<zX=2�L=�H=�mL=�X=��j=$x�=$��=�;�=L;�=���=s��=���=���=*�=��=� >�>��>4a>	>{>�2>�>��>ߑ >���=��=~��=�@�=�U�=�=�t�=0Q�=,� >��>n�>Y�>�   �   F�>p�>T>��>Y�=�R�=�u�=���=�K�=�K�=��=��="Ƣ=��=
B�=�u=�c=��W=�S=�AW=zub=dt=��=���=8��=M7�=�}�=���=�<�=���=���=���=n� >u�>�.>��>��>�>�>��>�n >�&�=z��=p��=do�=���=b��=��=bB�=FP�=���=�� > �>*�>�   �   �S>J�>��>��>&m�=�=��=���=��=���=�T�=9�=`��=�=���=|�=<�s=X�h=de=�h=$s=Z��=��=h�={O�=8��=�|�=�:�=���=@��=��=�{�=� >r>�>S�>�|>��>�Q>.��=Z�==�=0{�=BF�=���=*�=<�=�:�=`��=za�=Z8�=�E�=C >�g>�   �   ˰ >0�>�>!>,}�=2��=>��=��=���=l�=���=���=9H�=�7�=V0�=*��=�=��=@�{==Ha�=�-�=�k�=zz�=`��=�L�=	��=���=F�=�3�=*��=L&�=�s >��>H�>�>��>� >���=<�=P(�=8z�=>�=���=d��=�)�=�c�=Λ�=x��=���= �=���=�l�=Ŀ�=�   �   �Y�=v��=h� >$� >�}�=H�=���=F��=��=8��=��=���=�S�=�o�=|�=~�=cё=F(�=�p�=�̌=�&�=&1�=�v�=2f�=G`�=���=N�=���=��=6�=(U�=@��=�P >WR>=�>g� >�i�=���=��=��=Df�=���=�"�=��=��=R/�=Ă�=��=��=��=�K�=,��=@t�=���=�   �   v��=�s�=���=D��=,c�=��=d��=�#�=���=���=|��=\,�=�C�=���=�ۮ=3s�=�=켛=�(�=Q�=�#�=W^�=혭=jR�=��=n	�=J��=�,�=�T�=��=3�="��=' >Վ >G. ><�=��=���="��=���=�B�=���=�]�=���=_�=\^�=x��=T��=���=|#�=�7�=���=}�=���=�   �   �u�=ā�=�D�=&��=�%�=�
�=`2�=.��=|��=:	�=�q�=�&�=ޛ�=gL�=o��=�O�=v��=�٪=k�=n`�=�=4�=x<�=���=�	�=4��=,�=D�=���=�9�=�=<�=���=�V�=�_�=���=��=4@�=D��=���=���=���=2:�=^��=�*�=��=���=���=���=f��=��=��=T��=�i�=�   �   p��=�>�=�S�=���=J��=���=nY�=��=�S�= 3�=d�=4�=��=��=Vx�=��=��=Lع=���=�T�=��=���=U��=��=D�=\�=�l�=���=6?�=�S�=���=T��=���=NY�=��=VS�=�2�=� �=��=d��=`��=�w�=��=��=X׹=���=�S�=��=��=���=��=��=�[�=l�=�   �   ��=���=�9�= �=�;�=���=�V�=�_�=���=*�=�@�=ү�=J��=���=h��=;�=>��=�+�=h�=���=`��=���=)��=��=���=޷�=j�=v�=
��=E�=<��=�%�=�
�=>2�=���=*��=��=pq�=&�=.��=�K�=���=�N�=|��=�ت=j�=t_�=��=T�=�;�=ַ�=	�=���=�+�=�   �   �,�=�T�=f�=�2�=��=( >� >^. >��=\��=H��=���=t��=HC�=z��=�^�=T��=�_�=,_�=L��=��=���=.$�=�8�=j��=�}�=&��=ʬ�=�s�=���=\��=.c�=��=@��=�#�=T��=0��=���=�+�=C�=ä�=�ڮ=Mr�=�=�=�'�=&P�=#�=v]�=��=�Q�=���=��=���=�   �   ���=N�=�=
U�=2��=�P >cR>O�>�� >.j�=0��=V��=�=�f�=R��=6#�=��=��=0�=v��=z�=���=� �=4L�=���=�t�=��=Z�=���=z� >.� >�}�=6�=v��=��=l�=���=s��=��=ES�=o�=G{�=��=~Б=V'�=�o�=̌=�%�=Q0�=�u�=�e�=�_�=��=��=�   �   8��=
�=�3�=��=@&�=�s >��>V�>(�>��>-� >H��=��=�(�=�z�=�>�=P��=���=*�=zd�=^��= ��=��=v�=��=m�=��=� >G�>&�>%!>&}�="��=��=��=z��=�k�=���=x��=�G�=�6�=�/�=dߌ=B�=L�=��{=t=�`�=�,�=k�=�y�=ة�=HL�=���=�   �   �:�=���=��=��=�{�=� >!r>��>e�>}>�>�Q>|��=lZ�=d=�=�{�=�F�=j��=��=�<�=L;�=���=�a�=�8�=2F�=f >�g>
T>\�>��>��>$m�=�=���=`��=��=w��=�T�=��=眨=k��=��=p{�=��s=��h=e=��h=�
s=���=^�=��=O�=���=Z|�=�   �   ���=�<�=h��=���=���=k� >|�>�.>��>�>�>�>��>o >('�=���=���=�o�=���=���=,��=�B�=�P�=о�=�� >8�>=�>W�>}�>]>��>Y�=�R�=�u�=���=�K�=�K�=x�=.�=�Ţ=&�=�A�=�u=�c=�W=�S=�@W=�tb=@ct=a�=H��=븢=
7�=~}�=�   �   ^��=r��=���=�=��=� >�>��>8a>>�>�2>�>��>� >���=��=���=�@�=�U�=<�=u�=VQ�=A� >��>{�>g�>�F>L3>Tw>��>�I�=L��=��=Rn�=2��=��=�g�=R�=>�=�ȏ=2��=Tk=�yX=��L=��H=,mL=VX=<�j=�w�==�;�=&;�=���=�   �   �B�=:�=�\�=���=�{�=� >>y�>m�>��>�^>'�>@|>SF>O>f��=�6�=`��=�h�=L{�=�5�=p��=�) >�8>�S>VY>�!>c�>�b>x�>^>�D�=���=�B�=T��=��=�Z�=��=sЭ=�ߝ=�_�=��=��g=X�T=��H=��D=�H=L�T=�Pg=��=�[�=�=q7�=�&�=�   �   ���=���=���=,�="��=�� >�>��>:a>>�>�2>�>��>� >���=��=���=�@�=�U�=4�=u�=RQ�==� >��>z�>f�>�F>P3>Zw>��>J�=^��=(��=rn�=\��=��=�g�=��=��=ɏ=���=$k=�zX=��L=l�H=nL=&X=��j=Lx�=<��=�;�=`;�=���=�   �   ���=�<�=���=��=���=w� >��>�.>��>�>�>�>��>o >'�=���=���=�o�=���=���="��=�B�=zP�=Ⱦ�=�� >5�>?�>Y�>��>d>��>&Y�=�R�=v�=��=L�=L�=��=��=[Ƣ=��=PB�=Tu=�	c=��W=��S=�BW= vb=�dt=�=޴�=q��=y7�=�}�=�   �   ;�=��=b��=��=�{�=� >,r>��>k�>}>�>�Q>t��=\Z�=Z=�=�{�=�F�=V��=��=~<�=8;�=���=�a�=�8�=&F�=a >�g>	T>b�>��>ʅ>Fm�=:�=@��=���= �=���=2U�=��=���=V��=��=�|�=:�s=\�h=de=�h=s=���=R�=��=�O�=~��=�|�=�   �   ʃ�=z�=�3�=T��=t&�=�s >��>^�>0�>��>*� >:��=��=�(�=�z�=t>�=>��=���=*�=`d�=H��=��=���=f�=��=m�=
��=� >K�>0�>6!>T}�=^��=n��=L��=���=Bl�=D��=X��=�H�=�7�=�0�=���=��=4�=��{=P=�a�=*.�=6l�=�z�=ƪ�=M�=V��=�   �   D��=��=n�=TU�=r��=�P >rR>Y�>�� >.j�=*��=F��=��=�f�=>��= #�=��=l�=�/�=X��=`�=n��=j �=L�=���=�t�=��=$Z�=���=�� >@� >�}�=~�=Խ�=���= �=���=L��=��=bT�=]p�=�|�="�=ґ=�(�=�q�=�͌=M'�=�1�=8w�=�f�=�`�=���=��=�   �   <-�=U�=��=N3�=T��=? >� >g. >��=\��=:��=���=X��=0C�=\��=d^�=8��=�_�=
_�=$��=���=z��=$�=n8�=R��=|}�=��=Ȭ�= t�=���=���=fc�=�=���= $�=��=���=���=�,�=7D�=��=vܮ=�s�=��=���=O)�=�Q�=�$�=_�=���=�R�=���=�	�=���=�   �   ��=F��=0:�=T�=F<�=���= W�=`�=���=$�=�@�=���=0��=���=N��=�:�=��=�+�=B�=`��=8��=���=��=x�=���=ķ�=�i�=v�=��=.E�=h��=6&�=�
�=�2�=x��=Ή�=�	�=Zr�=4'�=e��=M�=��=HP�=8��=�ڪ=�k�=4a�=���=��=$=�=$��=(
�=���=t,�=�   �   $��=�?�=0T�=��=���=���=�Y�=�=�S�=3�=R�="�=���=��=9x�=x�=��="ع=���=�T�=��=͵�=2��=j�=(�=�[�=�l�=���=>?�=T�=���=���=���=�Y�=D�=�S�=z3�=��=��=���=���=�x�=R�=��=ٹ=v��=jU�=h�=���=���=�=��=~\�=�l�=�   �   Rv�=T��=ZE�=z��=8&�=�
�=~2�=>��=���=4	�=�q�=�&�=���=HL�=R��=jO�=L��=�٪=�j�=B`�=Ū�=�=S<�=l��=�	�=��=,�=<�=���= :�=:�=@<�=̦�="W�=<`�=.��=��=A�=D��=���=.��=��=�;�=���=v,�=	�=<��=��=P��=���=$�=��=D��=fj�=�   �   ��=:t�=���=���=hc�=
�=|��=�#�=���=���=n��=M,�=�C�=e��=�ۮ=s�=��=¼�=`(�=�P�=�#�=-^�=Ƙ�=ER�=Y��=P	�=8��=�,�=�T�=��=23�=N��=F >� >�. >��=���=���=��=���=�C�=
��= _�=���=t`�=�_�=���=���=0��=�$�=9�=���=�}�=z��=�   �   hZ�=���=�� >G� >�}�=l�=���=P��=��=2��=ܑ�=���=�S�=�o�=�{�=X�=?ё=(�=�p�=�̌=x&�=�0�=zv�=f�='`�=���==�=��=��=B�=@U�=l��=�P >�R>o�>�� >xj�=���=���=p�=Dg�=���=�#�=@�=�=�0�=��=�=��=!�=�L�=��=�t�=:��=�   �   � >`�>;�>:!>V}�=N��=N��=��=���=�k�=���=總=$H�=f7�=:0�=��=��=��=��{=�="a�=u-�=�k�=Wz�=C��=�L�=���=���=D�=�3�=>��=l&�=�s >��>q�>I�>��>P� >���=��=$)�="{�=�>�=ʬ�=p��=�*�=�d�=М�=j��=v��=��=l��=Vm�=P��=�   �   !T>p�>��>ͅ>Jm�=2�=$��=���=��=���=�T�=)�=O��=ۊ�=���=�{�= �s=�h=$e=ځh=�s=@��=��=M�=hO�=*��=�|�=�:�=���=F��=��=�{�=� >4r>�>|�>'}>0�>�Q>�=�Z�=�=�=�{�=G�=���=��=�<�=�;�=��=*b�=�8�=pF�=� > h>�   �   e�>��>k>��>&Y�=�R�=�u�=���=�K�=�K�=��=v�=Ƣ=|�=�A�=�u=�c=��W=��S=�AW=Lub=�ct=��=���=,��=D7�=�}�=���=�<�=���=
��=���=z� >��>/>��>�>�>>�>$o >Z'�=���=���=�o�=*��=���=f��=�B�=�P�=���=�� >J�>N�>�   �   �F>U3>]w>��> J�=X��="��=fn�=N��=��=�g�=y�=k�=�ȏ=i��=�k=(zX=$�L=��H=�mL=�X=��j=x�=��=�;�=B;�=���=t��=���=���=0�=$��=�� >�>��>Da>>�>�2>
>��>�� >���=�=���=�@�=�U�=X�=(u�=pQ�=J� >��>��>p�>�   �   2�>�>�>Ħ >2��=D��=.X�=J��=���=�t�=���=��=*_=�0=�
=@�<��<�xH<�/<p]G<�ć<�<��=(1=��_=���=8�=0´=	��=���=�|�=vW�=�v�=�>�%>�B>�~>� >O�>�>r� >d��=\��=R��=�"�=f`�=dy�=�k�=@$�=��=~G�=�>�k>p>�   �   ��>��>j�>� >$��=�2�=���=:��=���=���=&M�=���=L�b=�*5=g�
=>c�<p��<�X_<�3F<�^<Ĥ�<�?�<�a
=\"5=Jc=B4�=1�=�ĵ=�Q�=�l�=��=��=�q�=��>��>r>)>ޗ>�{>g>�_ >4~�=���=n8�=ę�=���=��=0��=D��=,)�=>�=W� >��>8>�   �   ֦>��>�>q[ >|�=���=��=�w�=�L�=��=�3�=VM�=��m=��A=f�=���<P��<�%�<<�<�J�<<}�<���<&�=�A=�m=Н�=�٣=���=(��=&�=8��=��=c�=��>�r>�>>|+>%a>>�a >��=ȁ�=RL�=\��=��=� �=�G�=df�=jg�=�#�=�`�=���=U� >9�>�   �   h>�>�I>���=$�=��=���=Dj�=�I�=�м=�k�=��=��~=|ZU=��.=�g=�(�<�3�<�|�<��<��<=X]-=(7T=�F~=���=���=�q�=:C�=��=��=��=hE�=�+>ؕ>��>�>c>Rf�=�Z�=	�=��=$$�=/�=0-�=8A�=�y�=(��=�3�=p�=�F�=�_�=�S�=4��=�   �   d��=z��=�6 >4��=D=�="$�=�{�=.;�=�x�=4q�=���=�j�=KɊ=o=\sK=��,=��=�=� =p�=Tb=��*=JfI=:-m=J��=�=�^�=���=��=�=ִ�=��=`�=� >Xg>rK>�R >@J�=,��=���=V��=���=~%�=`��=�J�="?�=���=r@�=�*�=L�=���=���=��=O�=�   �   Zj�=���=���=ʘ�=�D�=��=�`�=���=܄�=3�=��=�̩=��=��=m=5Q=p�;=D�-=��(=��,= �9=,�N=�Bj=?�=�Ɩ=~ɨ=4h�=f��=F��=h�=�*�=2��=x��=�d�=���=�V�=��=�c�=���=�T�=>��=���=�o�=<�=	p�=�;�=ɳ�=��=�n�=tN�=h�=�f�=ֵ�=&��=�   �   �=3�=���=@��=�(�=Z�=�r�=�m�=��=N��={��=�9�=qz�=��=9=��x=�e=�VY=<�T=�.X=�c=��u=��=4E�=�Ƥ=X��=;O�=L��=ƞ�=�]�=.��=���=f;�=�f�=�`�=�S�=�~�=z6�=���=��=��=P��=J;�=�,�=���=�r�=b�=��=B<�=r>�=:b�=�-�=^�=,��=�   �   r��=$��=���=4�=���=R_�=J��=@H�=`��=W�=�A�=e�=ig�=)��=���=(А=Nu�=B�=���=8g�=�:�=� �="��=~ݥ=�N�=�!�=���=��=���=<��=.^�=��=F��=��=�f�=
��=��=v��=���=)�=`��=b��=^�=�ӱ=Zݭ=XC�=�"�=�n�=~�=�E�=���=T�=:�=��=�   �   x&�=F�=���=��=LY�=ƌ�=�k�=6��=6i�=(��=x��=V��=�%�=���=��=�ߤ=��=�=%8�=NZ�=Ma�=^�=�ܫ=�M�=���=�s�=���=�&�=��=��=.��=\Y�=���=dk�=���=�h�=���=���=���=
%�=���=��=�ޤ=���=��=�6�=�X�=�_�=�=�۫=�L�=ɹ�=4s�=X��=�   �   <�=���=���=^�=��=R��=��=�f�=p��=B�=��=x��=�)�=^��=x��=��=ձ=�ޭ=�D�=H$�=>p�=��=G�=���=.��=�:�=���=���=���=���=V�=���=@_�=��=�G�=���=rV�=<A�=��=nf�=��=^��=�ΐ=�s�=��=[��=�e�=M9�=t�=�=fܥ=�M�=� �=��=�   �   ���=^��=T]�=��=���=n;�="g�=�`�=HT�=@�=7�=L��=F�=d�=N��=Z<�=�-�=���=�s�=��=(��=K=�=f?�= c�=�.�=
�=���=��=`3�=*��=Z��=�(�=@�=�r�=�m�=^�=���=ā�=�8�={y�=��=���=(�x=@�e=�SY=X�T=,X=Z�c=P�u=��=(D�=�Ť=���=�N�=�   �   ���=��=$�=�*�=��=|��=�d�=���=W�=0�=2d�=X��=�U�=��=���=�p�= =�=
q�=�<�=ȴ�=���=�o�=DO�=.�=Fg�=n��=���=�j�=8��=���=���=�D�=��=�`�=P��=l��=|2�=&�=�˩=�=��=�m=~2Q=Ț;=x�-=̨(=2�,=d�9=��N=�@j=>�= Ɩ=�Ȩ=�g�=�   �   8��=6�=��=���=ڬ�=`�=+� >kg>�K>�R >�J�=���=��=���=H��=8&�=*��=�K�=�?�=`��=6A�=x+�=��=H��=v��=|��=xO�=���=���=�6 >J��=B=�=
$�=�{�=�:�=jx�=�p�==�i�=vȊ="o=:qK=4�,=c�=m�=] =�=`=l�*=TdI=|+m=���=r�=E^�=�   �   pq�=�B�=���=Ə�=���=dE�=�+>�>��>�>>c>�f�=�Z�=�	�=���=�$�=�/�=�-�=�A�=�z�=���=x4�=�p�=:G�=4`�=�S�=���=�>�>�I>���=�#�=��=\��=j�={I�=gм=Fk�=f��=(�~=�XU=��.=f=�$�<�/�<�x�<���<� �<L=�[-=�5T=\E~=p��=O��=�   �   R��=���=�=$��=���=c�=ģ>�r>�>>�+>@a>2>�a >��= ��=�L�=¹�=l��=Z!�=H�=�f�=�g�=&$�=$a�=B��=x� >R�>�>�>�>u[ >z�=���=��=�w�=�L�=���=73�=�L�=��m=��A=�=���<���<�"�<D�<�G�<hz�<<��<�=�A=4�m=p��=�٣=�   �   �ĵ=zQ�=�l�=��=��=�q�=��>��>}>&)>�>�{>x>�_ >\~�=Ȓ�=�8�=���=���=V��=d��=x��=Z)�=l�=k� >��>F>��>��>n�>� >&��=�2�=���=��=_��=ʋ�=�L�=b��=��b=�)5=��
=�a�<ಓ<XU_<�0F<�^<X��<v>�<ga
=�!5=�Ic=4�=�0�=�   �   .´=��=���=�|�=rW�=�v�=�>�%>�B>�~>� >M�>�>n� >d��=\��=R��=�"�=l`�=fy�=�k�=@$�=��=�G�=�>�k>p>2�>��>�>Ħ >0��=B��=,X�=D��=���=�t�=���=��=_=��0=l
=�<ଈ<hxH<H/<0]G<�ć< �<��=01=��_=���=;�=�   �   �ĵ=�Q�=�l�=*��=���=�q�=��>��>}>')>�>�{>x>�_ >Z~�=ƒ�=�8�=��=���=J��=\��=n��=V)�=h�=j� >��>H>��>��>p�>� >4��=�2�=���=L��=���=��=>M�=���=��b=�*5=��
=d�<���<�Z_<�5F<^<䥒<�@�<�b
=�"5=dJc=h4�=+1�=�   �   ƺ�=W��=P�=X��=$��="c�=̣>�r>�>>�+>=a>3>�a >��=��=�L�=���=^��=J!�=H�=�f�=�g�=$�=a�=<��=p� >T�>�>�>�>�[ >��=���=��=�w�=M�=8��=�3�=�M�=>�m=��A=G�=z��<���<�'�<|�<�L�<T�<���<�=X A=ȱm=��=ڣ=�   �   r�=|C�=��=��=4��=�E�=�+>�>��>�>;c>�f�=�Z�=�	�=���=�$�=�/�=�-�=�A�=lz�=���=b4�=~p�=*G�=&`�=�S�=���=�>�>�I>���=4$�=F��=���=|j�=J�=Ѽ='l�=p��=��~=�[U=�.=Li=�+�<�6�<$��<��<��<~=�^-=L8T=�G~=b��=��=�   �   	��=��=\�=��= ��=��=<� >vg>�K>�R >�J�=���=��=ޖ�=4��=&�=��=�K�=�?�=@��=A�=Z+�=��=4��=d��=j��=tO�=���=���= 7 >t��=�=�=`$�=|�=v;�=!y�=�q�=��=/k�=�Ɋ=�o=�tK=H�,=��=��=� =\�=Dd=\�*=�gI=�.m=���=��=;_�=�   �   ���=���=��= +�=r��=���=�d�=���="W�=,�=0d�=F��=~U�=���=���=`p�=�<�=�p�=�<�=���=���=�o�=$O�=�=.g�=Z��=���=�j�=L��=п�=��=E�=h��=6a�=���=@��=|3�=^�=;ͩ=��=⢆=�m=7Q=��;=|�-=ȭ(=�,=�9=*�N=�Dj=�?�=�ǖ=ʨ=�h�=�   �   ���=(��=�]�=x��=��=�;�=Jg�=�`�=PT�=@�=7�=8��=,�=H�=1��=5<�=�-�=���=�s�=`�=���=(=�==?�=�b�=`.�=��=���=��=p3�=N��=���=�(�=��=@s�=Hn�=@�=ʤ�=��=H:�=={�=��=7È=��x=R�e=2YY=��T=41X=N�c=��u=��=F�=�Ǥ=���=�O�=�   �   @�=l��=���=~^�=h��=���=��=g�=z��=>�=��=d��=�)�=<��=V��=h�=�Ա=sޭ=vD�=$�=
p�={�=�F�=���=��=�:�=x��=���=���=��=��=0��=�_�=���=�H�=���=�W�=�B�=�=2h�=��=���=?ѐ=vv�=n�=��=_h�=�;�=�!�=!��=Wޥ=\O�=4"�=7��=�   �   t'�=�=n��=���=�Y�=
��=�k�=R��=:i�=$��=h��=B��=�%�=���=��=�ߤ=浝=��=�7�=Z�=a�=+�=�ܫ=�M�=���=�s�=���=�&�=��=0��=\��=�Y�=��=�k�=���=�i�=���=��=��=�&�=���=��=�=4��=;�=J9�=j[�=fb�=g	�=�ݫ=�N�=p��=�t�=���=�   �   b��=���=F��=��=8��=�_�=r��=TH�=d��=W�=�A�=N�=Cg�=��=n��=�ϐ=u�=�=���=�f�=w:�=� �=�=Jݥ=nN�=n!�=���=��=��=R��=Z^�=^��=���=�=\g�=ܥ�=��=���=��=�*�=1��=d��=��=$ֱ=�߭=�E�=W%�=Bq�=��=�G�=���=݀�=b;�=
��=�   �   ��=�3�=���=���=�(�=��=s�=�m�=��=F��=i��=�9�=Pz�=��==t�x=��e=lVY=̶T=n.X=��c=t�u=��=E�=�Ƥ=3��="O�==��=Ȟ�=�]�=T��=��=�;�=jg�=a�=�T�=��=�7�=���=��=&�="��=>=�=�.�=���=�t�=��=��=,>�=2@�=�c�= /�=��=6��=�   �   k�=���=���=&��=E�=L��=a�=���=���= 3�=��=�̩=��=졆=�m=�4Q=�;=��-=�(=��,=��9=��N=`Bj=�>�=�Ɩ=\ɨ=h�=Y��=H��=t�=�*�=h��=Ľ�=�d�=4��=pW�=��=�d�=Ԫ�=(V�=���=d��=Fq�=�=�=�q�=�=�=���=���=hp�=�O�=��=�g�=��=��=�   �    ��= ��=7 >���=~=�=J$�=�{�=8;�=�x�=(q�={��=�j�=0Ɋ=�o=sK=6�,=q�=��=w =�=b=<�*=�eI=�,m='��=��=�^�=���=��=(�=��=��=��=H� >�g>�K>�R >K�=��=���=~��=ސ�=�&�=Ц�=tL�=�@�=��=�A�=,�=��=���=���=���=�O�=�   �   �>7�>J>��=2$�=8��=���=Hj�=�I�=�м=�k�==d�~=JZU=��.=�g=(�<3�<P|�<��<�<�=]-=�6T=^F~=ڨ�=���=�q�=7C�=��=���=*��=�E�=�+>�>��>(�>cc>g�=V[�=�	�=��=(%�=20�=N.�=VB�={�=:��=�4�=�p�=�G�=�`�=8T�=ʷ�=�   �   �>%�>�>�[ >��=���=��=�w�=�L�= ��=�3�=MM�=l�m=��A=5�=*��<���<,%�<��<dJ�<�|�<P��<��=dA=�m=���=�٣=���=&��=,�=J��=��=(c�=գ>�r>�>>�+>Ya>Q>b >>�=j��=M�=��=���=�!�=fH�=g�=h�=p$�=`a�=~��=�� >k�>�   �   ��>��>y�>� >:��=�2�=���=>��=���=���=M�=���=<�b=�*5=S�
=c�<@��<HX_< 3F<�^<���<~?�<�a
=@"5=�Ic=74�=�0�=�ĵ=�Q�=�l�=��=���=�q�=��>��>�>/)>��>�{>�>�_ >�~�=��=�8�= ��= ��=|��=���=���=|)�=��=y� >�>S>�   �   P�>�>y?>p�=�r�=E�=t6�=��=���=��=p�a=��=Е�<�;P�1��ɼ����,���6��"-��K�\�ʼ �2�P�;�Ѵ<�� =N�d=)�=i/�=5��=��=�L�=̬�=R: >i>Ov>��>�">��>:>��=Z��=�Q�= a�=\�= d�=J��=���=��=�=­�=�i�=*� >r7>�   �   �q>�M>">l��="��=J��=���=
�=�7�=���=:�e=}�#=@��<=�;H�Pǹ��@�L�#�ؘ-�|V$����@��Ȑ�@�;�n�<�O%=�wh=!f�=O�=�n�=ڃ�=���=��=� >=�>�">�U>�>o1>3O >�e�=-�=�_�=�Q�=D9�=�9�=lc�=���=��=.C�=�	�=\��=IJ >��>�   �   �1>�^>o >\T�=p��=�~�=���=��=�Ͱ=TN�= Mq=>W1=��<�q5<�s��$l����޼�
��u�"�
�<�� ���@ꈻP�3<l��<�`2=�7s=J��=��=���=���=H;�=���=j��=�">=*>�>�>yS >�J�=��=���=���=��=���=���=h��=6q�=��=���=��=̘�=���=�  >�   �   �A�=��=��=�f�=R��= ��=�C�=d��=dy�=g��=H��=�(G=r�=��<`"�;`r�,�����¼`wԼ�Kļ�l��Є��4v;��<��=�)G=}'�=�=�̷=s}�=�V�=nQ�=���=T\�=�	>��>�� >���=�d�=��=|B�= ��=N��=���=x�=���=��=4��=@2�=���=���=:F�=Z��=��=�   �   և�=Bm�=��=$�=��=���=���=_#�=�ѽ=��=�z�=L�c=�*=��<q<�+c;����x�2��T��@7�d��`�:;X;f<\��<4(=�Fb=�K�=$a�=̏�=�P�=�_�=��=�c�=*��=\	�=(��=��=v��=x��=t��=���=$��=��=��=���=n�=0��=\>�=hD�=���=�$�=�	�=���=���=�   �    F�=��=��=�_�=V6�=���=��=�W�=�X�=�!�=.2�=�L�=^�P=A�=h��<X�<@<��; �;�Tl;pM	<To�<�B�<�B=|�M=�=�T�=۽�=Vq�=X��=l��=f6�=V�=���=l/�=B�=���=�<�=l�=���=���=�k�=	�=M8�=�[�=���=�g�=�a�=cq�=?�=pN�=� �=���=��=�   �   j��=8��=�O�=�;�=�$�=���=`�=���=[��=��=��=6�=��z=0N=�H$=e =0w�<���<8g�<�ן<���<f�<��=eI=n�v=�D�=|��=� �=��=���=\��=���=�}�=��=D��=�U�=X��=
�=���=*�=��=��=.��=Xy�=�̣=�ߡ=�Ԣ=Ĝ�=���=�r�=�~�=fc�=N[�=N��=�   �   
��=�W�=�h�=P��=���=p��=X[�=���=��=H�=pF�=ƒ�=�	�=�f=�Z[=\<=վ#=��=b�=�7=�o =��7=�V=��y=tH�=�=� �=Җ�=t��=��=2.�=�
�=��=���=�1�=ؚ�=z�=�B�=׉�=}�=�y�=�ˡ=̖=01�=V��=~O�=J��=�X�=N:�=��=�=Ċ�=@/�=�,�=�   �   ��=�I�=���=���=r�=�V�=�X�=2�=n�=�;�=�1�=���=="�=^͗=���=2�v=�b=��T=�hO=\�R=p�^=�q=t��=a��=K��=���=���=���=HJ�=���=���=~�=�V�=�X�=�1�=��= ;�=�0�=���=� �=�˗=֌�=x�v=�
b=x�T=�dO=D�R=�|^=x�q=С�=䤔=���=���=���=�   �   ��=��=j�=�-�=n
�=(��=���=R2�=d��=�z�=zC�=��=��={�=i͡=�͖=�2�=6��=^Q�=(��=�Z�=�;�=���=��=���=H0�={-�=���=4X�=Ni�=���=���=V��=[�="��=v��=AG�=rE�=���=-�=�c=W[=v<=��#==�=�=�3=�k =��7=N
V=��y=!G�=��=��=�   �   ���=���="��= ��=���=�}�=��=���=DV�=���=��=���=B�=�=f��=���=�z�=_Σ=+�=8֢=Z��=H��=�s�=��=zd�=8\�=��=���=���=P�=�;�=�$�=���=�=l��=���=��=��=�4�=�z=�N=EE$=u  =�n�<��<�^�<ϟ<`��<��<��=bI=Ąv=�C�=���=�   �   /��=�p�=���=2��=N6�=\�=֞�=�/�=��=D��=Z=�=�l�=���=���=m�=E
�=�9�=D]�=鸹=`i�=Vc�=�r�=:@�=�O�=��=���=���=�F�=
�=\��=�_�=R6�=���=���=jW�=3X�=� �=41�=ZK�=��P=�=h��<���<0<���;�x;@l;�=	<(h�<�;�<@=��M=���=�S�=�   �   �`�=V��=hP�=�_�=���=�c�=J��=�	�=x��=j�=��=��=4��=d��=��=��=��=���=@o�=V��=p?�=jE�=t��=t%�=T
�=���=��=<��=�m�=��=<�=��=���=z��=�"�=ѽ=��=�y�=$�c= *=p��<p
q<@�b;�έ��3��!T��O7�p����w:;�/f<8��<�(=Eb=
K�=�   �   v��=~̷=.}�=jV�=XQ�=���=p\�=�	>֐>�� >d��=e�=d�="C�=���=��=���=T�=���=��=��=3�=p��=j��=�F�=ڌ�=^�=.B�=^��=8��=g�=P��=���=�C�=��=�x�=ʜ�=���='G=a�= �<��;�}�0����¼�}Լ�Qļhr������v;��<��=`(G=�&�=�   �   �=���=���=���=4;�=���=|��=�">N*>�>�>�S >TK�=��=p��= ��=R�=���=���=���=�q�=P �=h��=J�=.��=,��=�  >�1>�^>o >hT�=f��=�~�=l��=���=NͰ=�M�=Lq=�U1=��<�j5<����Xp���޼�
��w�\�
�d�༸���������3<܁�<�_2=�6s=�   �   �e�=�N�=�n�=ȃ�=���=
��=� >B�>�">V>��>�1>JO >�e�=>-�=`�=�Q�=�9�=:�=�c�=��=�=jC�=(
�=���=^J >��>�q>�M>'>n��="��=B��=���=��=�7�=I��=��e=��#=|��<5�;���ɹ�"B���#��-��W$����<����0y�;�m�<�N%=fwh=�   �   /�=m/�=9��=��=�L�=Ь�=R: >h>Nv>��>�">��><>��=X��=�Q�=a�=
\�=$d�=N��=���=��=�=ĭ�=�i�=)� >p7>S�>�>y?>l�=�r�=E�=n6�=��=���=p�=D�a=��=x��<�
�;(�1��ɼ���2�,���6��"-��K�X�ʼإ2���;�Ѵ<�� =^�d=�   �   Qf�=6O�=�n�=���=���=��=� >H�>�">V>��>�1>IO >�e�=8-�=`�=�Q�=�9�=:�=�c�=ޱ�=�=`C�=&
�=���=YJ >��>�q>�M>->���=:��=`��=���=�=8�=���=|�e=ԗ#=0��<�A�;�
��Ź�@�p�#���-��U$�������������;p�<�O%=@xh=�   �   ���=d��=��=��=r;�= ��=���=�">V*>�>�>�S >NK�=��=d��=��=D�=z��=|��=���=�q�=< �=X��=<�=(��=$��=�  >�1>�^> o >�T�=���=�=ȇ�=��=�Ͱ=�N�=�Mq=X1=��<�v5<�h��$i��P�޼�
��s�f�
���༸����ވ�h�3<���<�a2=t8s=�   �   h��=>ͷ=�}�=�V�=�Q�=ڑ�=�\�=�	>ސ>�� >^��=e�=Z�=C�=���=���=|��=<�=���=x�=���=�2�=Z��=P��=�F�=Ҍ�=V�=2B�=j��=X��=<g�=���=>��="D�=���=�y�=֝�=ҵ�="*G= �=t�<�2�;�i�P�����¼DrԼ�Fļ�g���{��Uv;��<D�=(+G=
(�=�   �   �a�=C��=Q�=<`�=V��=(d�=t��=�	�=���=l�= ��=��="��=N��=���=���=��=���=o�=,��=L?�=LE�=V��=`%�=:
�=���=��=F��=�m�=��=x�=N�=��=��=�#�=ҽ=>�=�{�=�c=�*=���<!q<@Xc;����H�2�T��47��L����:;�Ef<ġ�<(=|Hb=xL�=�   �   z��=�q�=���=���=�6�=��=
��=�/�=��=D��=P=�=�l�=|��=���=�l�=$
�=|9�=]�=���=5i�='c�=}r�=@�=_O�=��=t��=���=�F�=&�=���=�_�=�6�=��=x��=NX�=`Y�=/"�=�2�=xM�=��P=��= ��<��<�M<���;��;��l;�Z	<�u�< H�<bE=��M=��=qU�=�   �   J�=���= ��=Ɗ�=���=~�="�=���=TV�=���=��=n��=#�=��=D��=���=�z�=.Σ=��= ֢=%��=��=�s�=��=Sd�= \�=���= ��=���=2P�=�;�=X%�=��=��=`��=��=x�=��=7�=D{=� N=�K$=� =4~�<��<�n�<�ޟ<h��<��<�=�gI=��v=�E�=N��=�   �   ���=��=L�=�.�=�
�=���=��=x2�=p��=�z�=hC�=ъ�=��=�z�=?͡=�͖=�2�=���=$Q�=蚇=LZ�=�;�=f��=��=΋�='0�=m-�=���=JX�=xi�=���=��=��=�[�=��=���=�H�=LG�=Γ�=�
�=�i=�][=�!<=V�#=�=�=�;=4s =ț7=�V=V�y=�I�=��=n!�=�   �   v��=�J�=t��=&��=��=
W�=Y�=22�=z�=�;�=�1�=���="�=3͗=`��=Ȱv=fb=�T=2hO=��R=�^=��q=:��=(��=��=|��=u��=���=XJ�=��=��=��="W�=NY�=�2�=�=x<�=�2�=���=b#�=�Η=���=Z�v=0b=�T=8lO=��R=��^=2�q=礅=���=b��=���=\��=�   �   X��=�X�=�i�=��= ��=���=�[�=���=��=H�=_F�=���=n	�=�f=LZ[=�<=^�#=��=��=c7=,o = �7=@V=D�y=BH�=��=� �=ǖ�=���=��=l.�=�
�=���=8��=�2�=���=n{�=BD�=ԋ�=��=9|�=�Ρ=Eϖ=�4�=ʓ�=�R�=���=\�=h=�=�=�=���=%1�=C.�=�   �   ���=0��=zP�=<�=Z%�=���=��=���=e��=��=��=�5�=��z=�N=�H$=� =Hv�<���<$f�<\֟<h��<B�<s�=�dI= �v=�D�=`��=� �=#��=���=���=��=~�=P�=��=�V�=���=��=R��=5�=)�=���=���=P|�=�ϣ=��=�ע=���=���=
u�=���=de�= ]�=���=�   �   "G�=��=�=
`�=�6�=���=6��=�W�=�X�=!�=2�=jL�=�P=��=���<t�<h><�݀;�; Ll;0K	<Pn�<�A�<xB=�M=� �=�T�=ɽ�=Vq�=l��=���=�6�=��=,��=0�= �=ʠ�=�=�=�m�=h��=���=n�=^�=�:�=q^�=��=�j�=xd�=�s�=@A�=fP�=��=8��=Z��=�   �   ���=�m�=.�=��=N�=���=���=o#�=�ѽ=��=�z�=�c=T*=���<�q<`&c;ഭ�h�2��T��B7� h�� �:;�9f<���<�(=�Fb=�K�=a�=ȏ�=�P�=`�=:��=4d�=���=�	�=޳�=��=���=���=���=&��=���= ��=�	�=���=7p�=H��=]@�=JF�=J��=0&�=�
�=$��=���=�   �   ~B�=���=���=Tg�=���=*��=�C�=m��=gy�=^��=7��=�(G=F�=h�<` �;�s�܏��d�¼(xԼpLļ�m�����`.v;8�<g�=�)G=b'�=ނ�=�̷=~}�=�V�=�Q�=ޑ�=�\�=�	>��>�� >���=ze�=��=�C�=T��=���=D��=
�=r��=L�=���=�3�=
��=���=DG�=<��=��=�   �   �1>�^>+o >�T�=���=�=���=��=�Ͱ=LN�= Mq=$W1=D�<8q5< u���l��(�޼�
��u�v�
���༈����숻 �3<��<�`2=|7s=:��=��=���=���=f;�=&��=���=�">k*>>�>�S >�K�=j��=���=���=��=���=��=n��=0r�=� �=���=��=���=p��=! >�   �   �q>�M>6>���=<��=Z��=���=�=�7�=���=$�e=c�#=��<�<�;���ǹ�A�l�#� �-��V$�������X��0~�;�n�<dO%=�wh=f�=O�=�n�=���=���="��=� >N�>�">V>�>�1>aO >�e�=p-�=@`�=R�=�9�=L:�=�c�=��=L�=�C�=R
�=���=oJ >��>�   �   b*>�� >B�=R��=./�=��=s�=jt�=ns�=E==r�< �r9̼̂�M�R��ný���s�����;����G�/`ý����M���ȼ )v:�k�<|BB=Ba�=$��=z�=[�=�&�=p��=�->l>�n>�>� >Ls�=LS�=�'�=\u�=���=P�=4��=4�=���=��=���=^E�=��=�f�=xY >�   �   ;� >�q >���=x��=dK�=>�=�G�=���= /�=��A=x��<���:4ﻼ'D��}������`޽8��<��:����޽N`������>�C�����g';�.�<6F=��= ݬ=Z��=���=L/�=H��=_� >�>�>��>�* >��=��=6��=���=���="�=@��=�= ��=���=��=�=:�=���=4W�=�   �   J�=:��=��=L��=��=*V�=���=Y`�=8A�=�O=�!�< ��;؎����'�Gn��<4���2˽��߽���4ཚ�˽嫽����X[(�쀊� ~�;���<8�R={��=N*�=C��=���=�A�=���=� >�j>nD>���=�^�=®�=�l�=�6�=X��=)�=~!�=��=��=��=���=���="?�=B.�=Һ�=�:�=�   �   h��=n��=��=J��=0�=�a�=���=�0�=�E�=��c=��=��p<��������UR��9��H���@��`
ǽ����F���a��x�T�Xm�����p�q<o2=|wf=)	�=�i�=>)�=�[�=P�=2{�=Bk�=&��=��=x��=t��=`��=�1�=���=��=���=�$�=W��=�	�=*��=���=���=���=@�=K�=�N�=�   �   ���=`��=d��="H�=�r�=���={y�=/��=袟=� =�5=PS�< T�;v��Z���V�	r��T藽�*��?����ć���Y�������`yr;V�<�s5=��==[9�=@v�=d�=6F�=^��=$��=���=2N�=4+�=(�=@��=�W�=��=d��=hW�=��=�"�=^ٶ=��=���=�!�=���=�H�=�n�=x��=�   �   45�=���=pH�=��=���=��=�!�=a�=柫=�%�=�]=�=�F�< �&����X�J>4��MS�^��U�̙7�z�`薼�ɞ�D׌<�S=�Z=α�=�ǫ=P�=�g�=���=B�=��= ��=�|�=bT�=��=���=��=F�=�C�=
�=��=���=Nw�=�{�=��=2¦=�<�=Ve�=#]�=�;�=��=�   �   xl�=X�=��=�G�=H��=���=��=ޡ�=L}�=���=���=:%I=��=�4�<`�;�I0��ϫ� ��<���0�$�����E� <Q:pȀ<|�=�)D=^��= ��=tͷ=7��=��=L��=vq�=�z�=�R�=�i�=�;�=,W�=n�=�W�=r�=e��=�֋=��=Ȱv=�\q=�/t=��~=�y�=r�=��=��=���=��=�   �   ��=�=���=���=|^�= x�=���=N��=���=��=5�=N�}=��E=�E=H!�<�k2<�B;��`� ���"��@%�: [<�<��=$�>=�w=|{�=o��=}�=��=��="��=P\�=�W�=j�=$��=�>�=
��=��=� �=��=6fp="+Q=�8=ܴ(=1^"=.&=��3=DwJ=�^h=���=ή�=���=6ҽ=�   �   1�=.��=�O�=R��=Vd�=ز�=,x�=��=�'�=Զ�=h!�=�9�=�
�=$�S=�
(=�=h��<P��<��<��<�?�<:,�<Zb =�tK=�y=f�=��=.�=���=0P�=���=ld�=���=�w�=t��=�&�=Ƶ�= �=�7�=��=��S=�(=z
=��<\�<���<���<�4�<�!�<�] =�pK=t�y=�d�=ҿ�=�   �   h��=��=.�=���= ��=f\�=$X�=��=���=�?�=J��=6�=�"�=� �=�jp=0Q=�8=<�(=�c"=n3&=��3=|J=,ch=x��=���=jë=`ӽ=���=��= ��=&��=�^�=�w�=.��=���=���=��=�3�=܄}=~�E=&A=��<�T2< �;�9a�0M��@U��@f�:E<�<M�=V�>=�w=3z�=�   �   ���=�̷=���=ʞ�=.��=�q�= {�=,S�=Rj�=�<�=FX�=To�=7Y�=2	�=X��=�؋=�=x�v=�aq=\4t=�~=|�=t�=ɉ�=���=���=��=Dm�=��=|��= H�=F��=j��=j�=;��=a|�=���=��=�!I=��=+�<�,;�`0� ܫ� ��8����(�0ɳ�ЫE���O:���<��=�&D=��=�   �   װ�=Dǫ=��=�g�=ҥ�=D�=:��=\��=^}�=U�=ԗ�=���=�=��=fE�=��=��=|��=Hy�=�}�=鮟=�æ=>>�=�f�=h^�=�<�=r�=�5�=��=�H�= �=���=���=P!�={`�=��=�$�=]=��=�>�< �8��&���ZD4��SS��^��#U���7��� 򖼀R���ό<�P=��Z=�   �   @�=J��=�8�=�u�=�c�=4F�=���=h��=��=�N�=�+�=�(�=P��=�X�=&�=���=�X�=d�=Z$�=�ڶ=,�=a��=�"�=*��=�I�=�o�=2��=D��=���=���=>H�=�r�=v��=y�=���=��=��~=x�5=M�<7�;|~���^�,�V��t��0뗽p-�����PǇ���Y�J������@Er;�P�<�q5=�   �   vf=��=]i�=)�=�[�=P�=V{�=xk�=v��=��=��=��=&��=v2�=���=��=η�=�%�=���=�
�=H��=���=���=���=�@�=�K�=�O�=Қ�=���=:��=X��=�=pa�=Q��=T0�=.E�=�c=��= �p<�������YR� <�����QC���ǽ����|
���c�� �T��s��@����q<�0=�   �   H�R=$��=*�=��=��=�A�=���=� >�j>�D>���=V_�=<��=Dm�=.7�=��=�)�=F"�=Ƚ�=��=P�=>��=>��=�?�=�.�=H��=;�=��=l��=�=^��= ��=V�=A��=�_�=�@�=dO=��<pq�;t���x�'��o���5��s4˽t�߽�����.�˽�櫽6����](������q�;(��<�   �   �~F=���=ݬ=G��=��=F/�=L��=h� >+�> �>��>�* >X��=��=���=���=��=��=���=v�=~��=��= �=f�=|�=Ծ�=dW�=N� >�q >��=~��=VK�=&�=lG�=Ǵ�=�.�=��A=t��<���:�񻼐(D��~������a޽6��=������޽a��(���Z�C�|���[';�-�<�   �   �BB=Ha�=.��=~�=[�=�&�=r��=�->l>�n>�>� >Rs�=JS�=�'�=^u�=���=X�=4��=<�=���=��=���=dE�=��=�f�=xY >c*>�� >@�=L��=$/�=���=�r�=Zt�=Vs�=�D==�q�< �r9P�̼^�M�z���ý�低�����B����G�)`ý����M�L�ȼ�1v:l�<�   �   �F=I��=Nݬ=~��=��=d/�=`��=o� >/�>"�>��>�* >V��=��=~��=���=��=��=���=n�=v��=��=�=b�=t�=ξ�=dW�=R� >�q >��=���=~K�=Z�=�G�= ��=</�=�A=4��<���:��4&D�7}��=���_޽����;��x���޽�_��䣒�"�C�� ��`t';@0�<�   �   0�R=䣏=�*�=���=6��=�A�=���=� >�j>�D>���=R_�=:��=8m�="7�=���=�)�=0"�=���=��=@�=.��=.��=�?�=�.�=>��= ;�=��=���=.�=���=B��=bV�=���=�`�=�A�=�O=�#�<���;������'�7m��	3��k1˽J�߽b����6�˽�㫽����NY(�\}�����;��<�   �   �xf=�	�=+j�=�)�=N\�=^P�=�{�=�k�=���=�=
��=��=��=d2�=���=��=���=�%�=l��=�
�=)��=���=n��=���=�@�=�K�=�O�=ؚ�=ҋ�=^��=���=��=�a�=��=@1�=^F�=�c=@�=H�p<��������QR�8��b���>��Vǽ����[��)`��.�T��g�� ����q<4=�   �   ��=���=�9�=�v�=~d�=�F�=ʀ�=���=&��=�N�=�+�=�(�=:��=�X�=�=���=�X�=?�=2$�=�ڶ=�=:��=�"�=��=�I�=�o�=(��=N��=���=���=�H�=,s�=��=�y�=���=���=x=�5=,X�<`k�;Lo��8V���V��o���嗽(��ҟ��X�P�Y���,��r;�Z�<�u5=�   �   ���=�ȫ=��=rh�=r��=��=���=���=x}�= U�=ԗ�=���=��=��=BE�=��=��=J��=y�=W}�=���=�æ=>�=�f�=L^�=�<�=n�=�5�=8��=�H�=V�=`��=���=F"�=�a�=���=�&�=4]=̞=8M�< X�����	�*94�LHS�Z�^�zU���7�bu��ߖ��Q���݌<wV=L�Z=�   �   ���=Jη=��=���=���=�q�=h{�=`S�=hj�=�<�=>X�=>o�=Y�=	�=1��=�؋=��=�v=6aq=�3t=��~=�{�=�s�=���=f��=���=��=Hm�=�=���=VH�=���=(��=l�=���=~�=���=Ȳ�=$(I=F�=�<�<��;�50��ī�������漐�����E� \R:@Ѐ<��=�,D=���=�   �   j��=R�=d�=���=���=�\�=rX�=�=���=�?�=:��=�=^"�=� �=Njp=�/Q=��8=��(=c"=�2&=4�3=�{J=�bh=:��=J��=@ë=Jӽ=���=��=X��=z��=_�=�x�=*��=��=x��=��=96�=@�}=�E=�I=L*�<P2<`�;�|`���p����͓:�n<'�<��=��>=�w=�|�=�   �   &�=���=�P�=2��=�d�=J��=zx�=.��=�'�=Ѷ�=V!�=e9�=z
�=īS=x
(=a=`��<$��<��<l�<�>�<�*�<�a =8tK=��y=�e�=���=#�=���=dP�=��=�d�=j��=�x�=���=v(�=ҷ�=�"�=�:�=N�=��S=*(=�=t��<��<d�<�<�I�<r5�<�f =zxK=P�y=vg�==ª=�   �   ���=��=���=���=_�=�x�=���=v��=���=��=�4�=�}=:�E=jE=l �<�i2<@9;��`�����(��@�:xX<��<,�=��>=rw=]{�=c��=��=��=h��=���=�\�=�X�=��=���=�@�=c��=��=
$�=l"�=�np=H4Q=��8=�(=Zh"=8&=H�3=D�J=gh=+=���=�ī=yԽ=�   �   n�=��="��=�H�=���=���=�=��=X}�=���=w��= %I={�=�3�<�z;�K0��Ы�p�ἤ����演���H�E��Q:Dǀ<��=l)D=<��=즞=|ͷ=Z��=X��=���=r�=�{�=�S�=k�=z=�=DY�=p�=�Z�=�
�=��=�ڋ=�=��v=�eq=h8t=  =�}�=�u�=L��=嵱=���=��=�   �   �6�=���=FI�=~�=`��=n��=�!�=6a�==�%�=�]=ɛ=�E�< (�x�����>4�FNS�t�^��U�z�7��z��閼�ݞ�(֌<TS=��Z=���=�ǫ=e�=h�=L��=��=���=��= ~�=�U�=���=���=0�=�=�F�=b�=��=4��= {�=@�=���=�Ŧ=�?�=h�=�_�=�=�=N �=�   �   ���=R��=��=�H�=,s�=���=�y�=G��==� =��5=�R�<�Q�;�v���Z�n�V�Lr���藽�*�������ć�D�Y��������qr;HU�<�s5=��=硠=m9�=hv�=Xd�=�F�=���=ދ�=���=^O�=�,�=�)�=6��=�Y�=J�=��=EZ�=��=�%�=Nܶ=��=���=$�=4��=�J�=np�=���=�   �   H��="��=���=���=|�=�a�=ŉ�=�0�=�E�=��c=��=��p<����$���^UR�:�����)A���
ǽ�������1b���T�Tn��x�� �q<)2=Fwf=&	�=�i�=c)�=.\�=bP�=�{�=�k�=޼�=t�=���=���=���=:3�=���=��=Ƹ�=�&�=���=��=E��=���=`��=Z��=�A�=PL�=P�=�   �   ��=���=P�=���=B��=PV�=���=d`�=:A�=�O=�!�<��;@����'�gn��d4���2˽ܹ߽��g���˽M嫽%����[(�����|�;��<�R=x��=T*�=]��=��=�A�=���=� >k>�D>8��=�_�=���=�m�=�7�=���=p*�=�"�=x��=p�=��=ܳ�=А�=8@�=6/�=���=t;�=�   �   e� >�q >*��=���=~K�=N�=�G�=��=/�=��A=H��<���:xﻼ'D��}������`޽T��<��V����޽i`������t�C���� e';�.�<,F=��=&ݬ=e��=
��=h/�=l��=y� ><�>3�>��>�* >���=�=̬�=2��=t��=��=���=��=���=d��=h�=��=��=��=�W�=�   �   �=6��=���=��=lW�='��=�p�=R��=� &=�ES<�����\�� ���h�}�)�2�J���d���u�l\{�j�u�Z�d���J���)�`�������X�`����9n<��-=4܆=��=�b�=��=P��=���= � >�e>2i >���=6��=:`�=���=��=���=ʑ�=R�=\�=ֈ�=d�=���=���=*��=�>�=zo�=�   �   L�=L��=*�=���=B��=k�=��=m�=|�*= 3m<<����R�ʹ�:� �y%�y�E��_�</p���u�Wp���_�P1F�.�%��� �������N�0�~�0?�<412=bs�=Z�=e��=�2�=l��=�$�=�_ >B� >��=�g�=�A�=pV�=�_�=:�=��=�t�=��=t:�=f��=l��=`�=�y�=��=J �=���=�   �   ���=V��=M�=H�=�=N�=��=t��=�+9=hg�<��2�ڸ4�*���2콪:��Q8�-�P�!�`�d1f���`��BQ�i�8�;���U콃>���E2�#����<�d?=�=��=�v�=`u�=��=�%�=��=B-�=��=\��=�W�=T7�=F%�=v��=��=�=<N�=���=׌�=�U�=���=�7�=P��=2?�=�'�=�   �   $��=.l�=d�=$��=���=0>�=�_�= ��=ظO=���<��ֺ����e��.�ʽQ���"�ݱ9�f_H���M�ͻH�T:���#����m�˽�؆��;����4��<,OT=�}�=��=���=���=<'�=���=�_�=J��=Zl�=���=��=���=F�=�%�=��=�Y�=OG�=P �=�w�=�n�=�k�=+��=��=r��=���=�   �   ���=��=��=x��=4��=*��=�A�=�%�=��l=XM=P/(<Tޒ�PD���O۽��p(��k)��).���)�~�H��oݽ���1G�pe���''<,�=�go=Z�=��=n��=�=r��=���=���=&��=�`�=���=#:�=�J�=�Ȳ=��=R�=��=��=R��=|�=�ã=���=t�=\��=���=���=�   �   Pr�=Ԃ�=�^�=Z2�=�G�=D�=!!�=�1�=)�=px>=HU�<��E�l)^��$��]�н����9�u
�����\��o�ӽ�a���kd��� ��$�<dl==�c�=��=F��= 6�=���=�y�=v8�=0��=�g�=st�=���=�ϳ=t7�=�P�=+L�=�wt=F�e=|�_=�b= �n=�,�=�K�=���=l�=�5�=
�=�   �   -y�=@��=��=�v�=�o�=$-�=dg�=K�=@�=ڱm=8=X��<�m��غ�B�O�7U��tN���^½(�ɽ9�ý)���������W�����pC����}<�D=�pj=;�=��=)�=R~�=�h�=��=��=���=��=Ľ=t��=�=�ƀ=�JY= �5=;=2�=�� =2�=J=ff-=��N=�>v=2 �=�=Ñ�=�   �   ��=��=ؘ�=���=~��=T��=���=%��=8�=b��=�Z=(8=�l�<��e�싳�(����O���q��D~��t���U���#�x�ż����0 `<^=f�S=h�=�L�=d��=@D�=2]�=��=���=�<�=m��=�=���=�"�=(�e=h�0=0q�<��<�K=< 0�;�|;`�;@[$<�͒<$��<�z%=�Z=Ї=�Π=�   �   �?�=͹=q4�=���=B��=>��=&�=��=�y�=��=8��=��W=��=XV�<�η;���P���`Y̼ �ἀ�Ҽ,����� _P;�'�<�a=
JN=T�=�@�=ι=5�=���=X��=��=��=	�=ix�=���=T��=�W=F�=�I�<���;PP�������j̼��ἴ�Ҽ���P�� �O;p�<�\=�EN=NR�=�   �   �=�K�=���=�C�=
]�=��=N��=�=�=p��=m�=R��=%�=�e=�0=�}�<�!�<8i=<�m�;`�|;�C�;px$<�ے<l��<,�%=��Z=҇=lР=��=��=t��=��=���=��=��=N��=�=б�=�Z=B3=(a�<�Zf�4��������O��q��M~��t�\�U���#���ż�Ŀ��
`<�=��S=�   �   nj=:�=*�=��=$~�=�h�=D�=D�=���=��=�Ž=F��=$�=�Ȁ=DPY= �5=�$=��=P� =г=�=Pl-=(O=xCv=A"�=��=)��=Ez�=
��=���=w�=�o�=�,�=�f�=f�=�=��m==\}�<��������O��Y��S���c½�ɽ��ý����$咽:X����� o��x�}<�@=�   �   �i==�b�=,�=ۯ�=�5�=���=�y�=�8�=���=�h�=�u�=.��=�ѳ=�9�=8S�=�N�=$}t=��e=�_=��b=`�n='/�=�M�=���=&�=7�=8�=6s�=|��=R_�=�2�=�G�=��=� �= 1�=�'�=Du>=@M�< ����P�60^��(����н$���;�lw
� ��Pa��u�ӽxe�� rd�$!� =�D�<�   �   ȅ=�eo=��=���=F��=�=���=���=:��=��=�a�=ؕ�=�;�=�L�=Yʲ=��=n�=,�=8��=~��=� �=tţ=L��=�=Ƌ�=���=~��=`��=D�=��=���= ��=���=A�=�$�=��l=fJ=� (<\璼�D�=���۽���*�n)��+.���)�����Lrݽ����5G�$m���'<�   �   h��<�MT=|}�=���=���=���=^'�=���=�_�=���=m�=���=��=���=��=0'�=�=E[�=�H�=��=Py�=8p�=�l�=a��=*��=V��=���=���=�l�=��=4��=���=�=�=>_�=q��=�O=���<�%׺����g����ʽ����"���9�=aH�h�M���H��U:��#�0����˽�چ��>� d���   �   ��<�c?=��=��=pv�=Xu�=���=�%�=0��=�-�=d��=��=PX�= 8�=(&�=h��=��=�=RO�=���=ۍ�=�V�=���=�8�= ��=�?�=d(�=���=���=(M�=T�=�=�M�=��==z*9=�c�<H�2���4�����4��;�S8�w�P�x�`��2f��`��CQ�|�8�(��`W��?��H2��!#��   �   >�<�02=>s�=B�=R��=�2�=v��=%�=` >W� >��=h�= B�=�V�=f`�=��=���=u�=���=;�=��=��=��=�y�=:�=� �=��=v�=l��=*�=���=0��=�j�=̛�=�l�=��*=�.m<�����R�δ�ο ��y%�+�E�ԫ_��/p���u��Wp�P�_��1F���%��� �������N�H�~��   �   p:n< �-=@܆=��=�b�=��=V��=���=�� >�e>6i >���=<��=8`�=���=��=���=Α�=V�=\�=ֈ�=
d�=���=���=,��=�>�=|o�=�=4��=���=��=\W�=��=�p�=7��=E &=xDS<����\�� ���h���)�L�J��d���u�t\{�m�u�V�d���J�ҝ)�R�ݜ��X�X������   �   �@�<�12=�s�=��=���=�2�=���=(%�=` >\� >��=�g�=B�=�V�=^`�=��=���=u�=���=�:�=܋�=ܡ�=��=�y�=0�=� �=��=��=t��=**�=���=^��=/k�=(��=(m�=��*=�4m<����R�̴�� ��x%��E���_��.p�A�u�hVp��_��0F���%� � �1�����N�Д~��   �   ���<�e?=��=�=�v�=�u�=(��=&�=N��=�-�=f��=��=HX�=8�=&�=V��=��= �=<O�=���=ȍ�=�V�=���=�8�=���=�?�=j(�=���=���=NM�=��=Z�=hN�=8�=Ր�=�,9=�i�<��2��4�󾢽�0��9��P8��P� �`�<0f���`��AQ�`�8�L��'T�$=���C2��#��   �   @��<�PT=�~�=���=(��=���=�'�=(��=`�=���=m�=���=��=���=��='�=��=![�=�H�=��=/y�=p�=�l�=D��=��=H��=���=���=�l�=��=���=��=�>�=2`�=���=P�O=<��<�wֺ����c���ʽ�|�"�]�9��]H��M�4�H��R:�"�#����7�˽�ֆ��8� Ŗ��   �   ��=vio=!�=���= ��=��=��=��=^��=���=�a�=̕�=v;�=mL�=6ʲ=屧=B�= �=
��=P��=b �=Hţ=%��=��=���=���=|��=p��=l�=J��=��=���=���=<B�=V&�=��l=�O=�:(<(ג��	D����[۽t���&��i)��'.���)��
����lݽ���,G�^���3'<�   �   o==e�=��=��=�6�=Z��=Xz�=69�=��=�h�=�u�="��=�ѳ=^9�=S�=|N�=�|t=V�e=��_=�b=�n=�.�=�M�=���=�=�6�=2�=Ds�=���=�_�=�2�=�H�=��=�!�=�2�=/*�={>=�[�<�q��\;ἴ#^�p!����н���~7��r
�����X����ӽ�^��
fd���`���!�<�   �   �sj=B<�=��=��=�=pi�=��=��=���=��=�Ž=1��= �=�Ȁ=�OY=��5=0$=L�=ȍ =6�==�k-=�O=�Bv="�=��=��=Nz�=2��=��=�w�=�p�=�-�=2h�=:�=f�=��m=�"=���< E����x�O�qQ��WJ���Z½վɽ��ý�3ݒ���W��������P�}<H=�   �   ��=)N�=\��=E�=�]�=��=���=�=�=���=r�=L��=�$�=��e=��0=}�<� �<g=<�h�;��|;`>�;�u$<Hڒ<@��<�%=@�Z=�ч=XР=��=��=���=P��=0��=��=p��=!��=a�=Ҵ�=��Z=h<=�v�<��e��~�������O�l�q�<~���t���U�h�#��ż c��04`<�=��S=�   �   ZB�=?Ϲ=6�=���=��=���=��=�=�y�=��=*��=n�W=]�=�U�<pʷ;��������Z̼����Ҽ������ TP;,&�<6a=�IN=�S�=�@�=6ι=X5�=T��=���= ��=��=��=�z�=|��=扊=��W=��=pa�<� �;����x����I̼x��(�Ҽh堼�����P;x2�<|f=NN=�U�=�   �   �=� �=Z��=���=H��=���=���=[��=N�=e��=�Z=�7=l�< �e����������O�z�q�TE~���t�h�U���#���żp����`<�= �S=\�=M�=���=�D�=�]�=��=��=d>�=���=��=ឥ=�&�=`�e=�0=4��<.�<Ѓ=<��; �|;�z�;�$<�<���<"�%= �Z=�Ӈ=�Ѡ=�   �   i{�=��=p��=�w�=�p�=�-�=�g�=v�=P�=ұm==䆋< q��Ȼ���O��U���N��W_½��ɽ��ý����mᒽ��W�0����H��`�}<?D=�pj=";�=
�=x�=�~�=�i�=��=�=���=��=�ƽ=䮪=�='ˀ=$UY=X�5=X*=��=R� =��=Q=�q-=O=�Gv=#$�=d�=���=�   �   2t�=X��=`�=23�=�H�=��=f!�=$2�=))�=^x>=�T�<�����E��)^��$����н����9�?u
����Y]����ӽFb���ld��켠 �`�<.l==�c�=��=���=�6�=X��=�z�=�9�=���=�i�=�v�=���=@ӳ=V;�==U�=�P�=�t=��e=�_=|�b= �n=a1�=�O�=���=��=r8�=b�=�   �   0��=��=���=*��=���=���=�A�=�%�=��l=HM=x.(<�ޒ��D�N���۽@���(�l)��).��)���z��poݽ���1G�xf��8&'<�=vgo=s�=L��=���=��=.��=~��=���=���=�b�=���=�<�=�M�=�˲=γ�=O�=�=4��=r��=u"�=8ǣ=���=��=	��=���=r��=�   �   N��=m�=�=���=��=z>�=�_�=6��=�O=d��< �ֺ���e��X�ʽk���"� �9��_H���M���H�@T:���#�����˽�؆��;�� ��̮�<(OT=~�=1��=���=���=�'�=j��=z`�=t��=�m�=���=��=���=��=�(�=r�=�\�=jJ�=`�=�z�=�q�=
n�=t��=��=$��=\��=�   �   B��=��=|M�=��=V�=NN�=�=���=�+9=8g�<p�2��4�E���42콽:��Q8�D�P�<�`��1f���`��BQ���8�Y���U콴>��@F2�#�D��<�d?=!�=��=�v�=�u�=<��=0&�=���=.�=؜�=���=�X�=�8�=�&�=F��=��=�=JP�=���=ǎ�=�W�=���=f9�=���=T@�=�(�=�   �   ��=���=B*�=���=b��=$k�=��=
m�=x�*=�2m<`����R�ʹ�A� �y%���E�*�_�K/p���u�Wp���_�`1F�<�%��� �����N���~�?�<012=ls�=k�=v��=�2�=���=>%�=$` >p� > 	�=Dh�=jB�=(W�=�`�=&�=��=�u�=
��=v;�=^��=V��=< �=Vz�=��=� �=0��=�   �   F��=J��=F:�=�*�=|"�=��=u�=JP =���;^S��a������<�J�v����x|���BľU�оpiվѾB[ľ�����g��"Fv�o�;�J������(�����<��*=�݊={1�=<��=���=���=���=�=҂�=�#�=p��=̕�=@6�=ʎ�=�W�=8�=`3�=L��=H��=��=,S�=��=���=$��=]�=�   �   �(�=�q�=6|�=���=t�=���=>�="8%=��	<�=���f��![ �-8��^q��Q��,ꬾ1b����̾�HѾ�;�������K����p�h87�_��kᕽ�t� U/<�E/=8Q�=���=���=��=/�=RP�=64�=��=0,�=hR�=�=��=6��=���=��=��=��= .�=��=J��=.��=�F�=���=���=�   �   ���=��=�/�=8�=�Z�=�O�= Ջ=�3=��Y<Ȟ��N��,��F�*��ea�V��a���g ��Q��HKžwB��b���΢��>��ea��C*���FX�������y<�[<=���=V@�=`|�=Ό�=��= [�=P��=���=B@�=L��=6/�=���=(\�=<ɹ=n��=q�=�.�=�ܶ=�1�=ٝ�=�X�=�t�=���=���=�   �   "(�=F��='�=���=8��=��=RH�=:J= ��<�X��Y�I�Ƚ���>mH��Dy�oY��򋣾���0����㮾����ؒ�j,z�SI�$���Ƚ�V�X�F�Я�<�Q=L5�=ʺ=^F�=���=2x�=j��=�8�=���=�?�=���=���=��=�٧=É�=�R�=��=䵖=�j�=�k�=��=�`�=(S�=L��=L`�=�   �   T��=�4�=�3�=���=!�=���=�ќ=��f=���< X�\��hΜ�Z�����(���T�B�{�4��<0��𿚾�����͍��}��V�8�)�2���+՝�n�� ��9��=�k=�=�5�=���=4��=�)�=(��=ζ�='j�=��=u�=v4�=F��=���=ܲo=`=��Y=��\=T�h=��}=��=%��=��=[9�=���=�   �   %5�=<��=./�=t�=}�=�=4��=��=X-=�Iw<l5����U�c#������*�S�L�O�g��Hy�J���z�2[i�n�N�f-����_�����Z���� �r<|�-=�>�=���=�=�8�=���=���=��=�	�=Uͼ=�*�=Zf�=X�y=N�N=�(=�\
=��<@��<`_�<` =�p=�wB=`Ul=<i�=�T�=�b�=�   �   N��=���=��=��=%`�=/*�=��=z��=nw^=�H�<@P�;,�ؼ0r��+���t��� ���2���A��EG�`�B��4�,{�@���n½N�{����`�&;�_�<�|\=��=Mɳ=���=��=
/�=���=
��=u:�=��=/�=j%U=�.=��<@JK< �B;��R� ����r�����:�� <ح<�5=v�F= �=���=�   �   ��=rh�=b��=��=���=r8�=P�=�C�=��=d�A=��< EF�XE��
d�/?���+ؽ	���T�N��6]�#� ��cݽ�<���`p�؛����U��@�<I;=�؅=%�=(ƽ=���=9�=���=���=�p�=���=r#�=0== ��<��*<�޻4ǳ�v�
���*�&f7�H(/�&����ɼ4#����;��<��/=�t=�   �   �x=���=ҡ�=���=W��=xB�=�2�=kܷ=���=�t�=n�5=�v�< E�:|��V<.�|�����-ǰ�:d���沽jĠ����
;�\Ǽ�ں�<D�+=Ćx=ۅ�=���=��=t��=<B�=�1�=\۷=6��=�r�=@�5=�i�<�P�:\&��zF.�D|��ǜ�wͰ��j���첽Rʠ������;�|!Ǽ��ں4s�<~�+=�   �   :E;=Pׅ=-�=�Ž=���=f�="��=���=r�=���=�%�=�	==��<�*< �ݻ������
���*�[7�T/������ɼ0#����;�"�< �/=X�t=ɒ�=�i�=1��=��=���=8�=��=aB�=�=�A=d
�<��G��U�ld��D���1ؽ���bX�����`�[� ��iݽB��jp�@����,V��6�<�   �   �W�<�y\=��=�ȳ=p��=��=|/�=���=6��=	<�=���=��=8+U=J5=4��<�kK<�YC;@R��r�� (��@ܐ:�� <��<v<=�F=X"�=���=ļ�=���=Q�=��=`�=�)�=��=B��=�s^=�?�< "�;d�ؼ�r��0���z��$�: 3���A�GIG���B�]�4�:~����fs½.�{�Ш��N&;�   �   8sr<��-=�=�=��=��=�8�=���=���=Զ�=�
�=�μ=�,�=�h�=��y=��N=��(=�c
=h��<���<�n�<�'=�w=�}B=�Zl=�k�=�V�=!d�=V6�=��=�/�=��=e�=�~�=j��=X�=� -=@8w<�@����U��'�����o�*���L���g�~Ly����!z�|^i�l�N�-�Ύ�.�����Z�Д���   �    ��92�=d�k=`=�5�=���=v��="*�=��=ط�=wk�=���=�v�=�6�=���=Y��=��o=`=��Y=�\=�h=@�}=���=P��=洭=�:�=���=L��=�5�=84�=ā�=�=���=�М=x�f=���< ������ќ�K����(�M�T�5�{��5���1������<���ύ��}�V�K�)������ם�����   �    �F����<jQ=�4�=�ɺ=XF�=��=�x�=��=f9�=���=*A�=���=1��=���=�ۧ=苞=U�=M��=��=�l�=�m�=��=Ub�=�T�=t��=>a�=�(�=���=\'�=���=��=h�=�G�=R
J=��<�X���Y��Ƚl��;oH�Gy��Z��H���䦮������䮾����(ْ�l.z�I�����Ƚl�V��   �   h�����y<�Z<=P��=1@�=\|�=���= ��=z[�=ʨ�= ��=A�=@��=H0�=���=r]�=�ʹ=豴=�r�=&0�=B޶=%3�=��=�Y�=nu�=H��=P��=��=:��=�/�=&8�=�Z�=wO�=�ԋ=t�3=��Y<�����K�꽊�*�!ga�,��O���c!��V��LLžpC���b��zϢ��?��Jfa��D*���sY���   �   4v弰R/<�E/=Q�=���=���=���=$/�=�P�=t4�=��=�,�=�R�=��=���=݇�=o��=���=̉�=��=�.�=���=��=���=HG�=4��=���=�(�=r�=H|�=���=�s�=̞�=��=:7%=x�	<A���g���[ ��8�m_q�zR���ꬾ�b���̾/IѾy;2������rK���p��87����ᕽ�   �   ������<��*=�݊=�1�=<��=���=���=���=�=؂�=�#�=v��=ȕ�=F6�=̎�=�W�=?�=d3�=R��=I��=��=,S�=��=���=&��=]�=<��=H��=@:�=�*�=l"�=�=u�=P =p��;�S��a��	 �ù<�t�v�#����|���Bľ_�оtiվѾ<[ľ�����g��Fv�S�;�.��k����   �   r�Y/<�F/=�Q�=3��=���=��=>/�=�P�=x4�=��=�,�=�R�=��=v��=ԇ�=e��=���=���=}�=�.�=���=֩�=���=@G�=,��=���= )�=0r�=b|�=���=;t�=+��=j�=�8%=��	<h<��if���Z ��8�^q��Q���鬾�a���̾/HѾ~;D������J����p��77�b�������   �   h���0�y<]<="��=�@�=�|�=8��=P��=�[�=Ԩ�=&��=
A�=4��=40�=���=b]�=�ʹ=ұ�=�r�=0�=*޶=3�=���=�Y�=`u�=<��=R��=��=V��=�/�=x8�=&[�=!P�=�Ջ=�3=�Y<P���3�����^�*��da�����������p��bJž�A��-a���͢�@>���ca��B*�J��V���   �   x�F�|��<�Q=6�=�ʺ=�F�=~��=�x�=��=r9�=���=$A�=���=��=s��=jۧ=ɋ�=�T�=(��=�=�l�=om�=b�=:b�=yT�=l��=@a�=�(�=���=�'�=N��=���=X��=�H�=�J=<��<��X���Y�'�Ƚn���kH��By�`X��ʊ��E�������F⮾�����֒�r*z��I����GȽ,�V��   �    _�9p�=H�k=�ß=�6�=H��=���=r*�= ��=��=|k�=���=�v�=�6�=���=4��=>�o=�`=<�Y=��\=��h=��}=S��=(��=̴�=�:�=���=^��=�5�=�4�=P��=��=���=dҜ=�g=�< ���,���˜������(�`�T���{��2���.��n���#���̍�\}�OV�4�)�����gҝ�����   �   ��r<��-=�?�=���=��=d9�=r��=���=��=�
�=ϼ=�,�=�h�=��y=D�N=z�(=zc
=l��<���<�m�<'=(w=�}B=lZl=sk�=�V�=d�=n6�=N��=0�=D�=E�=��=.��=��=L-=�Xw<�+����U�������*���L�E�g��Ey���Kz�"Xi���N�� -�Y��������Z�T����   �   �g�<�\=d��=aʳ=���=ȭ�=0�=��=_��=<�=���=��= +U=�4=h��<�iK< QC; R��w���-���Ɛ:� <��<�;=��F=7"�=x��=ռ�=���=��=��=�`�=+�=��=���=�z^=�P�<�w�;�ؼ�r�^'���o�����2���A�YBG��B��4�Lx����Fj½Ν{����`�&;�   �   M;=\څ=r�=Cǽ=���=8�=���=<��=Hr�=���=�%�=�	==�<��*<��ݻ����~�
�P�*��[7�/�����ɼ #����;�!�<��/=0�t=В�=�i�=���=��=���=g9�=e�=�D�=N�=\�A=d�< �D��6�0d�C:��&&ؽ���Q���Z�&� �X^ݽ�7��JXp�4��� gU��J�<�   �   ��x=n��=���=8��=x��=EC�=3�=�ܷ=㷟=�t�=T�5=Lv�<�9�:h���<.��|������ǰ��d��粽�Ġ������
;��Ǽ�*ں ~�<��+=��x=���=��=���=L��=tC�=�3�=�ݷ=J��=yv�=�5=��<��:���:3.��|�
���x���i^���ಽ򾠽~��� ;�` Ǽ�<ٺ|��< �+=�   �   ���=k�=f��=���=���=*9�=��=�C�=��=p�A=P�< TF�8F�Bd�y?���+ؽn	��,U����s]�d� �WdݽQ=���ap�D��� �U��?�<�H;=�؅=e�=�ƽ=t��=X�=%��=��=�s�=L��=�'�===��<�+<@�ݻ����<�
���*��P7�D/�����ɼ��"���;/�<B�/=��t=�   �   Z��=��=q�=��=a�=�*�=�=���=�w^=�H�< O�;��ؼ�r�,��Hu��!���2�&�A��EG���B�L�4�n{�~��+o½�{�4�� �&;,_�<�|\=G��=�ɳ=S��=ԭ�=h0�=���=|��=�=�=v��=��=�0U=p;=��<P�K<`�C;�~Q� -�� 䈻@�:H� <���<�B=lG=�$�=n��=�   �   �7�=:��=�0�=��=F�=��=���=��=|-=�Iw<�5���U��#��*����*���L���g�*Iy�����z�u[i���N��-��Ė��>�Z�����r<|�-=�>�==��=X9�=���=���=��=�=�м=�.�=�j�= �y=H�N=,�(=�j
=`�<���<�|�<f.=~=ʃB=�_l=�m�=�X�=�e�=�   �   ^��=�6�=5�=���=��=j��=�ќ= g= �< ������Μ����� (�ǇT�n�{�.4��X0����������͍�8}��V�p�)�����x՝���� |�9��=R�k=*ß=86�=<��=$��=�*�=г�=��=�l�=$��=�x�=�8�=��=Ь�=�o=�`=:�Y=n�\=`i=4�}=ʸ�=V��=���=t<�=,��=�   �   �)�=z��=�'�=v��=���=��=�H�=rJ=L��<`�X�:�Y�n�ȽԻ�YmH��Dy��Y���������I����㮾����ؒ��,z��I�K���ȽZ�V�h�F����<�Q=~5�=Xʺ=�F�=���=y�=���=*:�=~��=FB�=K��=���=2��=^ݧ=ٍ�=W�=Z��=��=�n�=ho�=4�=�c�=�U�=���=6b�=�   �   ���=���=40�=�8�=&[�=�O�=FՋ=�3=��Y<���c��G��V�*��ea�`��m���u ��b��\Kž�B�� b���΢�?��;ea��C*�2�kX��(��� �y<�[<=���=�@�=�|�=D��=���=�[�=L��=���=�A�=��=@1�= ��=�^�=�˹=8��=�s�=v1�=�߶=^4�=)��=�Z�=Lv�=��=��=�   �   >)�=Zr�=�|�=���=@t�=��=N�=38%=��	<�=���f��&[ �68��^q�R��2ꬾ7b����̾�HѾ;ǅ�����%K����p�x87���~ᕽ�t��T/<F/=HQ�=��=���=��=V/�=�P�=�4�=6�=�,�=RS�=��=
��=s��=��=T��=p��=3�=v/�=L��=p��=8��=�G�=���=F��=�   �   ؎�=���=��=���=޶=�@�=^�-=���;T�������(!���l�����Siʾ-��b4����W	$��D'��$���4��z�9�ɾ(���X�j��������vc�X�$<j\:=@��=�.�=V�=�y�=*D�=Z:�=��=� �=���=(p�=��=�<�=&g�=��=f��=ny�=E�=�ž=�Z�=�+�=d2�=HG�=�1�=�   �   �"�=��=�/�=���=�_�=8��=��1=�<~J��	��*��ng��]���]ƾ���	����!!��=$��!����a�	������ž����r�e��}�����Vt���=<�k>=n=P��=|��=@��=l��=|��=���=�7�=�7�=L�=���=���=0<�=���=�$�=���=Y
�=P��='�=K��=�o�=4L�=2��=�   �   ���=��=�L�=���=Pɸ=�V�=�?=�[<���%��t��W���������b�������1`�aq�Zz��������ᾰ���D2���BV�Ǣ�ɳ����ּ�H�< AJ=��=��=���=|�=n��=��=�^�=�n�=�=>��=lR�=F�=���=1
�=�8�=�L�=(1�=|�=�m�=\�=��=bO�=f`�=�   �   ~�=4c�=0�=�7�=�Ǻ=a2�=T�S=仫<(l���������,�>�z@��zI��� ̾2�y����
�5��z�
�r������̾է��YW���c>����8���l������<��\=z$�=��=���=N �=l��=vI�=<`�=���=�[�=��=�'�=�=�s=H�c=L�\=��_=�pl=2׀=�֎=��=�=8-�=3�=�   �   a��=���=���=�e�=ڼ=�v�=��m=l�<�덻�vA�`�Ƚ`[��_�G�������;k����L��H��}:�üξ&!���ۑ�?�`����ϋȽ<,?��sY��4=��t=�q�=�U�=�f�=�!�=t
�=���=���=�^�=���=4�}=�gQ=*=��
=8��<���<`��<��=��=��C=�ln=B��=���=/9�=�   �   �ů=�H�=�)�=P��=�m�=9U�=ڡ�=&�*=��8<d�ּ`���k��t�3��am�Қ���y���4��=�˾7�о��̾�;���ʬ�����p�@�5�ؘ��F��D;ټ@?<<��-=Xˇ=u9�= �=�H�=I:�=�&�=Fs�=z��=�a�=�R=�S=t��<��#<  �5@K׻x����� `�P�;�1�<�,=�B=��|=r=�=�   �   �9�=☫='ӻ=��=
��=��=F��=��Z=��<P|����*��������}6�#�e�mȇ�Co���A��6���壾V����V��pi�n�9���������1��o����<��Z=�ӕ=���=���=��=s;�= ��=U��=�w=��0=�-�<@z�; zY����¾.��Q�2Z_���V�&A8�`���#��@��:|#�<� =pwh=�   �   ��b=,��=
��=�3�=J�=���=iģ=��=�B5=�y�<P�T��E�b	���� �LU'���I�*e���v�C�}��Bx�f�g��,M� 4+�|���]��:hR�H�}�p,�<n0=Ę�=Kg�=h^�=访=n��=�$�=֥�=T�n=��=���<�5 �����qg�����u��5�׽��m�ڽ�ƽ������w�^
��ND�@�M<T�=�   �   nD=d�m=���=��=j��=��=�5�=S:�=\2u=�A =��g<�1j�ȁ8��Ĝ���ڽ5	�����0-���2�<�.��}!�4��h��?��P�H�g�� 6<bI= �m=Τ�=ȴ�=���=x�=5�=�8�=2.u=4< =��g<Uj�t�8��ʜ��ڽ5	����5-��2���.��!���I�E��V�H�dw��@�5<�   �   �!�<�0=t��=�f�=(^�=��=(��=&�=���=@�n=.�=��<X ����feg����~n��k�׽3�཮�ڽ�xƽ7�����w���� +D��N<"=��b=���=��=X4�=T�=^��=jã=��=H>5=�m�<�T���E�:��� �EY'�\�I��e���v�I�}��Gx��g��0M��7+����.c��qR���}��   �   ������<ځZ=�ҕ=5��=ח�=N�=�<�=���=p��=�w=.�0=�=�<�Ī;�OY�x��F�.�֝Q�M_���V��48���������:�2�<T� =||h=�;�=F��=Ի=���=���=~��=4��=h�Z=���<P�����*�����1��p�6�T�e��ʇ��q�� D���8��裾ɠ���X��]i���9����-����1��   �   �Eټ@0<<&�-=�ʇ=9�=�=I�=$;�=(�=u�=���=nd�=h�R=h[=�ȸ<8�#< `<7��ֻ���P�������N�;�B�<4=,B=�|=�?�='ǯ=�I�=^*�=���=�m�=�T�= �=��*=H�8<��ּd���p����3�hem�霒�/|��u7���̾؝о�̾8>���̬����
p���5�6����I���   �   �0?� �Y��2=�t=xq�=�U�=�f�=H"�=p�=��=p��=a�=��=�}=fnQ=h*=x�
=�
�<�<���<d�= �=@�C=hrn=Ľ�=��=�:�=���=p��=6��=f�=�ټ=Rv�=��m=H�<����|A��Ƚ�]�ʥ_�����!��ݾ;Wm�K�FO�����<�Ǿξ�"��~ݑ���`����َȽ�   �   ����Ä����<��\=0$�=��=,��=� �=$��=nJ�=�a�=8��=�]�=�=m*�=��=��s=D�c=\�\=��_=Tvl=�ـ=;َ=��=���=�.�=T4�=�~�=�c�=t0�=�7�=�Ǻ=�1�=��S=���<�s��������0�>��A���J��W"̾
�u����
�;��w�
�_����쾔�̾���\X��Be>�9���   �   ���X�ּTF�<P@J=��=��=��=X|�=��=���=�_�=�o�=L�=���=T�=�G�=z��=*�=�:�=�N�=3�=�}�=No�=��=��=hP�=0a�=t��=:�=$M�=���=ɸ=\V�=t?=��[<$���&��Bu���W�r���/���dᾡ��V���`�r�{�1��X���ᾍ����2��DV�����   �   ���u���=<`k>=^=N��=���=f��=���=���=���=n8�=N8�=�=r��=���="=�=~��=�%�=z��=F�=+��=�'�=���=p�=�L�=���=
#�= �=�/�=ؓ�=r_�=�=�1=0�<FL��
������ng�/^��g^ƾ� ��	�"���!�:>$�J!�F����	�W��Y�žֱ���e�~��   �   ����c���$<�\:=R��=�.�=Z�=�y�=,D�=\:�=�=� �=���=0p�=��=�<�=-g�=�=l��=ry�=E�=�ž=�Z�=�+�=h2�=HG�=�1�=Ў�=���=��=t��=�ݶ=v@�=�-=���;���J����(!���l����riʾJ��n4�Ķ�]	$��D'��$� ��4��z�!�ɾ���0�j�h���   �   �����r�(�=<�l>=�=���=���=���=���=���=���=n8�=F8�=��=l��=���==�=r��=�%�=l��=8�="��=�'�=���=p�=�L�=���=#�=�=�/�=��=�_�=h��=h 2=h�<�I�Z	������mg�X]��f]ƾ���t�	�n���!�~=$��!�����	�:��e�ž�����e�}��   �   .�����ּ�L�<�BJ=��=���=|��=�|�=��=���=�_�=�o�=F�=���=�S�=�G�=h��=�=�:�=�N�=�2�=�}�==o�=��=��=dP�=:a�=���=d�=pM�=V��=�ɸ=;W�=�?=��[<����#��;s���W�ۍ��F����a�d������_��p��y����%���᾽���x1���AV�����   �   ����������<��\=R%�=X�=���=!�=T��=�J�=�a�=<��=�]�=��=W*�=��=`�s=��c=�\=��_=vl=�ـ=َ=��=���=�.�=W4�=�=d�=�0�=b8�=�Ⱥ=3�=�S=<��<pf��ň��M����>��?��MH��H̾�	쾚����
�D����
����P�쾡�̾����FV���a>�����   �   ('?��4Y�8=��t=�r�=|V�=�g�=�"�=��=,��={��=a�=	��=�}= nQ=*=�
=�	�<<�<ط�<��=��=��C="rn=���=��=�:�=���=���=���=�f�=�ڼ=�w�=ڹm=�<�΍�0rA�_�ȽvY���_�������ʺ;�h侩�J����[8�̺ξc��yڑ���`������Ƚ�   �   80ټ�P<<�-=�̇=�:�=�=�I�=�;�=D(�=u�=���=gd�=6�R=&[=�Ǹ<��#<  57��ֻ ������`��pJ�;�A�<�3=�B=��|=�?�=Dǯ=�I�=�*�=Z��=�n�=WV�=#��=T�*=�9<�{ּ�\��Mg��֩3��^m������w���2����˾Ęо �̾�9���Ȭ�� ��|�o���5�p����B���   �   pB����<�Z=2Օ=���=��= �=�<�=���=���=w=�0= =�<���;PQY����в.�|�Q��M_���V��58����\�� ��:�1�<� =f|h=�;�=���=�Ի=D��='��=< �=���=�Z=���<�P���{*�+���n���z6�h�e�RƇ��l��?���3��㣾����T���i�%�9� ��+�����1��   �   �7�<�!0=���=�h�=�_�=6��=���=�&�=駗=t�n=8�=ē�<x ����eg����n����׽����ڽyƽ����Z�w�� �8-D��N<� =�b=��=���=5�=|�=¶=�ţ=:�=G5=܄�<ЕT�|�E�2���� ��Q'���I��e�>�v��|}�>x���g��(M�\0+�V��{X���_R��}��   �   �N=H�m=���=7��=핻=��=�6�=�:�=�2u=�A =нg<�2j�"�8��Ĝ�6�ڽ`	�����0-�Ŕ2�~�.��}!�s�����?����H�h��� 6<^I=X�m=4��=p��=���=�=a7�=�;�=x6u=�F =��g<�j�(x8�𾜽_�ڽ� 	����V,-�I�2��.��y!�������P9����H��V���6<�   �   ��b=���=���=�5�=��=���=�ģ=��=C5=,z�<��T�>�E��	��ǣ �tU'�#�I�be��v���}��Bx���g��,M�C4+����*^���hR���}�L,�<�0=��=�g�=\_�=V��=v��=�'�=���=�n=�=P��<p�������Yg�R���g��)�׽χ�g�ڽ�qƽ���w����`D�h1N<=�   �   �=�=��=�ջ=ʤ�=8��=���=���=H�Z=���<0|��*�����<���}6�P�e��ȇ�ao���A��36���壾~����V���i���9���������1��q����<
�Z=>ԕ=X��=���=� �=�=�=W��=z��=#w=P�0=L�<��;�(Y���򼪦.���Q��@_�̍V� )8���`���@��:�A�<�� =��h=�   �   �ȯ=7K�=�+�=���=�n�=�U�=F��=��*=��8<t�ּ`���k����3��am�蚒��y��5��^�˾_�о��̾�;���ʬ����p�|�5�4���_F���;ټh?<<�-=�ˇ= :�=�=J�=P<�=q)�=�v�=֭�=�f�=h�R=pb=hظ<(�#< P�7P�ֻ�q��L���(�p��;�R�<;=ZB=D�|=�A�=�   �   ��=���=B��=�f�=�ڼ=rw�=L�m=4�<pꍻ�vA�y�Ƚv[�	�_�X�����ʼ;k����L��n��:��ξI!��ܑ�v�`�����Ƚ~,?��sY�D5=(�t=Tr�=^V�=�g�=>#�=��=h��=��=c�=x��=��}=�tQ=B!*=��
=��<��<��<��=�=��C=xn=.��=��=�<�=�   �   ��=�d�=F1�=�8�=�Ⱥ=�2�=ЗS=l��<�k���������>�>��@���I��� ̾G쾅����
�D����
������<�̾򧨾pW���c>����Y���p������<h�\=�$�=2�=���=x!�=���=tK�=�b�=���=a_�=�=�,�=/�=��s=Мc=�\=|�_=�{l=f܀=�ێ=��=���=F0�=�5�=�   �   ,��=��=�M�=r��=�ɸ=
W�=(?=��[<p��%��t��W�����"����b�������:`�lq�ez������Ϗ�ƍ��W2��CV�ޢ�峟���ּI�<dAJ=,�=|��=���=�|�=n��=T��=l`�=�p�=p�=���=�U�=xI�=:��=��=n<�=�P�=�4�=��=�p�=&�=	�=jQ�=b�=�   �   j#�=R�=0�=&��=�_�=X��=" 2=��<rJ��	��0��ng��]���]ƾ ﾼ�	����'!��=$��!����h�	������ž������e��}�����dt���=<�k>=�=���=���=���=��="��=T��=�8�=�8�=��=.��=`��=�=�=_��=�&�=\��=#�= ��=�(�=���=�p�=6M�= �=�   �   ,��=���=�/�=!��=�=zK=�]^<v����½�+/�"4���ۻ��������f�6���P���d�$�q��}v��r��e���P���6��6��n��0_��y��m+�!?������4�<�jY=��=�b�=���=�l�=�	�=(��=FD�=á�=ً�=j\�=�X�=���=6�=$�=8�=�"�=
n�=NO�=ø�=�c�=���=��=�   �   ���=�[�=(�=�[�=.ƛ=H�N=x�v<�n�bW��J�*�:0������4������{3���L��`���m��Cr���m��a��L��\3�\k�C���������!'���x�缐�<�\=`��=��=@��=�G�=���=(��=�4�=f��=�{�=-`�=���=z0�="0�=�+�=�[�=l��=܈�=�2�={��=�2�=���=��=�   �   H_�=���=~^�=���=:֝=Y=8��<�ϼ�)��hy���t�C������pa�z�)�^1B�~^U�/�a���e���a��U�'bB���)�J�k@�ͫ�-rr�h��n ��܏�� ��<(�e=:�=��=� �=���=��=��=|��=�2�=��=�2�=��=�Ky=.�h=��a=��d=|�q=Q��=���=�ȡ=�}�=n)�=v�=�   �   �l�=���=>��=^��=ٲ�=li=���<�u��)��d���Y�l0���ξ�W�4���Z1��*C���N�=�R���N���C�t�1�m#�c���ξ�ښ��<X��	�������M���<`$t=Lq�=	��=�R�=���=:��=���=��=��=���=~=^=B7=f	=@?=hO�<���<>�=b�+=��O=��y=��=#�=v�=�   �   S��=	��=�<�=c?�=8��=V�|=~�=�3��h�I�ݽb�6���p��E��И����N�+��H6��9���6�|,���9A�&�⾒*���H����6�� ܽ\�D� Ո�\W=�̂=ʐ�=��= H�=�g�=��=�I�=�&�=�\]=�!=�:�<��R<��8;`�y��Ի�ȣ��:�c<Dɰ<�=��K=��=B'�=�   �   
��=�@�='�=���=��=��=�6=|U<��q/��&��(�W�OI��B&�������W��~���������>�?n���徐ֽ�������Y������p�㼈�a<X�:=��=�ީ=�i�=|s�=��=P�=�xz=<5=� �<0��;�=S���0��T��Kb��Y�|�:����XE�� ��:��<t�"=��i=�   �   �KZ==Q�=���=���=�Φ=W�=��^=@��<`z��ZH�Y�ͽ�z#���e��:�����%TԾ��R��u ��-��-��c`־�̸�rd����i��&��)ҽ�M�0Pѻ@3�<��`=��=|��=gl�=���=@T�=H�h=��=0hl<�S.��~�*�{�o���Ͻ��k�𽞐�dս�h��5K��,�)� :~��!<=�   �   P =0�Y=�f�=���=��=B��=��=j54=��<L����z�����w&�2�^��u���â����¾JZǾ��þ�·�����X|zc�z+�RI�8p��������s<��0=.x�=\��=\o�=<q�=�i�=\�d=�_=�Q<�r���<^��u��������Tz1�A�tG�żB�|�4�^���� �B񾽞�r�P�Լ���;�   �    ��;�Y=�h=�˒=�Q�=Tߢ=�}�=F�n=��=�<�ǼV��%w׽LO��~C��j��f��~o��V2���P��
��N�n�e�H�ӌ��c὘鉽0����;x^=@�h=�̒=�Q�=�ޢ=�|�=��n=$�=��<D�Ǽ]%��~~׽�S���C�nj��i���r���5��T������n�6�H�����j�*�*��   �   Գ��@�s<N�0=1w�= ��=�o�=3r�=uk�=,�d=Df=�s<�]��0^�Cn��dw����u1��A���F�\�B�^�4����d� �꾽��r���Լ�Λ;8=n�Y=Gh�=���=��=���=o�=614=�Ӆ<h���n�z�1���{&��^�Vx���Ƣ�|��v�¾�]Ǿ=�þCƷ����� �
c�=+�aO��t���   �   X�M�Pzѻ,�<��`=v�=���=%m�=Z��=IV�=Ĺh=�=��l<).�<r�Ĳ{�g��T�Ͻ|�N�𽫇��vս�`��3D����)��~���!<�=�PZ=S�=���=��=�Φ=��=��^=t��<�����H���ͽB~#���e�B=������uWԾ����U���v �|1�����c־�ϸ��f��t�i�3�&��.ҽ�   �   d�����㼠�a<:�:=�=�ީ=Vj�=�t�=���=��=�~z=n
5=�<pF�;@S����N0�2T�j=b��{Y��x:�:���.����:H�<V�"=,�i=��=*B�=�=Y��=��= �=�6=XjU<d�弪3�������W�yK���(����㾒�� ��Z��n��v �?@��o�o���ؽ�������Y�8���   �   �ܽ��D� d��dU=Ẑ=���=~��=�H�=$i�=o�=L�=c)�=Vc]=��!=�L�<�R<`�9;`Dy��bԻ�p����:`�<�ڰ<̛=<�K=p��=n)�=�=,��=�=�=�?�=�=ľ|=�}= ���>�I��ݽ��6�F���r�����3��g����+�sJ6���9�)�6��},�Q��zB�G��R,��;J����6��   �   B�f�����M���<�#t=:q�=O��= S�=Ƞ�=��=U��=�=d!�=z�=D^=4I7==8G=�_�<���<̺=x�+= P=��y=T�="�=�=	n�=���=���=p��=���=�i=���<x�u�P,����W�Y��1��Dξ�X�a��\1�B,C���N���R���N���C���1�u$�D��ξ�ۚ�H>X��   �   D�����,��� ��<��e=�9�=C��=0�=J��=���=4��=���=84�=��=�4�=k�=�Py=\�h=8�a=��d=h�q=���=���=�ʡ=x�=�*�=��=
`�=���=�^�=���=�՝=�Y=l��<Hϼ�+���z�f�t�W�����6b�Z�)�U2B��_U�:�a���e���a��U��bB���)��J�jA��ͫ�Usr��   �   "'���������<�\=b��=��=p��=�G�=<��=���=^5�=7��=�|�=8a�=��=�1�=j1�=-�=8]�=���=���=�3�=b��=I3�=Z��=���=���=\�=@�=�[�=�ś=��N=��v<Rp��X���*��0��v������p��_|3���L���`���m�Dr�3�m�[a�o�L�]3��k����n���Z����   �   �l+��>��������<DkY=4��=�b�=���=�l�=�	�=6��=JD�=ʡ�=��=w\�=�X�=��=<�=$�=8�=�"�=n�=LO�=Ƹ�=�c�=���=��= ��=���=�/�=��=��=*K=\^<��)�½,/�F4��ܻ�і�����|�6���P���d�,�q��}v��r��e���P�q�6��6��n��_���x���   �   !'���H����<�\=�=��=���= H�=J��=���=f5�=4��=y|�=2a�=��=�1�=^1�=-�=,]�=���=���=�3�=^��=D3�=X��=���=���=0\�=p�=�[�=^ƛ=��N=��v<�m��V����*��/�������񾹹��{3���L���`���m�Cr�.�m�ca���L�P\3��j���𾆣�������   �   B������������<��e=�:�=���=��=���=؝�=@��=���=54�=��=�4�=Y�=�Py=2�h=�a=��d=:�q=���=���=�ʡ=h�=�*�=��=$`�=���=_�="��=�֝=4Y=(��<�ϼ�(���x���t���������`���)��0B��]U�B�a���e���a�(�U�IaB�4�)�aI�A?�,̫��pr��   �   v�A�����M����<�&t=Ar�=���=�S�=��=���=l��=�=_!�=l�=�C^=I7=�=�F=_�<���<��=2�+=�P=L�y=E�=�=�=,n�=���=)��=4��=���=Di= ��<h�u��'����b�Y�P/��ξW�3���Y1��)C�@�N��R�5�N�L�C�C�1�Y"�t�� ξDٚ��:X��   �   ,�۽��D� ��Z=(΂=���=P��=tI�=|i�=��=L�=d)�=Dc]=��!=,L�<�R< �9;�Jy�0fԻ�t����:��<ڰ<~�=�K=a��=t)�=��=��=$>�=~@�=N��=��|=\�=������I��{ݽE�6�@�Tn��2�ᾚ��}����+�*G6�m�9��6�|z,�x���?���⾼(��]G��m�6��   �    ����b<��:=" �=:�=@k�=(u�=��=��=�~z=j
5=��<�D�;�S�`��0��T��=b�L|Y�vy:�����/��@ԯ:��<*�"=>�i=I��=�B�=��=W��=�=0�=�6=�U<���+�����"�W�mG���#��F��k�����ƚ��������<��l���3Խ�������Y�Z���   �   (�M�0ѻ�<�<|�`=��=��=n�=�=�V�="�h=<�=p�l<�).��r�&�{�Wg����Ͻg|罣����FwսGa���D����)��~�x�!<�=QZ=`S�=\��=��= Ц=��=,�^=<��<@L���
H���ͽ�w#���e�c8��T���QԾ��뾘N��Ks �J*��Ї�J]־ʸ�b����i��&��$ҽ�   �   @�����s<~�0=#z�=��=q�=s�=l�=ƍd=�f=�s<�]��L0^�ln���w����Hu1��A�%�F���B���4������ �b꾽�r�\�Լ�͛;^=�Y=�h�=���=���=���=��=�94=`�<����x�z����t&�ʂ^��r�����������¾�VǾf�þĿ�������댾�uc���*�-C�Lk���   �   ��;,d=��h=�Β=�S�=��=�~�=T�n=.�=��<�Ǽl��Ow׽iO��~C��j��f���o��v2��Q��-����n���H���4d��鉽��p��;�^=H�h=�͒=NS�=��=��=��n= =��<��Ǽ���mp׽KK��yC��j��c��~l��H/���M��*
����n���H�����\��㉽ ��   �   �=��Y=jj�=f��=Զ�=s��=��=B64=���<������z�����w&�R�^��u���â�7���¾lZǾ�þ÷�����|�zc��+��I�hp��������s<��0=�x�=���=5q�=�s�=wm�=�d=xl=��<4J��H$^�Kg��Yo��\��4p1��A���F�-�B�i�4���G� ��⾽x�r��}Լ��;�   �   tVZ=YU�=���=���=;Ц=Y�=��^=���<�w��LH�g�ͽ�z#���e��:�����ATԾ+��=R��(u ��-��Y��`־�̸��d��Əi�A�&�;*ҽD�M��Nѻx4�<�`=��=��=�n�=&��=rX�=.�h=��=��l<P.��f�^�{��_��7�Ͻ�s罞��꽲nսRY��Y=���)�@�}���!<�=�   �   |��=$D�=��=Է�=�=��=�6=x~U<d��n/��/��:�W�^I��T&�������h������������>�Vn�ܟ徶ֽ�Χ���Y����P��X�a<^�:=r�=�=�k�=v�=���=��=0�z=85=,"�< ��;(�R����R�/���S��/b�nY��k:��������:�'�<X�"=��i=�   �   ۟�=ï�=�>�=�@�=<��=��|=H�=�$��8�I�%ݽo�6���p��V��ۘ����_�+��H6�"�9���6�|,����NA�K�⾲*���H����6�� ܽZ�D� ��� X=u͂=Б�=���=+J�=�j�=2�=:N�=,�=�i]=J�!=d]�< �R<`<:;`�x��Ի0�� 3:�<�<b�=¯K=2��=�+�=�   �   xo�=���=���=t��=���=hi=���<��u��)��f��%�Y�v0���ξ�W�=���Z1��*C���N�P�R���N���C���1�#�t���ξ�ښ��<X�
�������M�8��<X%t=
r�=��=T�=ܡ�=���=���=�=�#�=,�=J^=�O7=D=�N=�n�<���<"�=R�+=<	P=�y=��=&�=��=�   �   �`�=P��=x_�=E��=�֝=�Y=��<Hϼ�)��ly���t�J������va���)�h1B��^U�<�a���e���a�$�U�6bB��)�J��@�0ͫ�Crr�v��p ������̬�<��e=v:�=���=��=��=���=F��=��=�5�=� �=�6�=��=�Uy=<�h=(�a=��d=&�q=ښ�=Ī�=�̡=��=,�=��=�   �   Z��=�\�=��=\�=hƛ=��N=P�v<rn�_W��L�*�<0������9�� ���{3���L��`��m��Cr���m��a��L��\3�bk�N�� ��� ����!'���\����<N�\=���=��=���=6H�=���=<��= 6�=���=X}�=/b�=.��=�2�=�2�=B.�=i^�=Ц�=��=�4�=G��=4�=��=,��=�   �   X	�=���=�]�=�j�=��r=g�<t���k쭽T+��u��qʾ�
�\2���[�����B���u��6"��c!��(��>w��ђ��\���[���1�K	�.Ⱦj��j{&�������i�<��=Ju�=NR�=L��=�F�=H�=�i�=��=��=Fz�=X��=�Ä=�oy=T�r=��u=��=}�=`�=.��=�e�=��=���=�   �   ��=p"�=���==,�=�t=X!�<�b��j���ɟ&�|[��$Lƾ�r��/���W�*�~�e���ɝ�9Y���O���c���ԝ��a��\~�:W��V.����6ľ�*��T@"��D���k��lA�<��=��=���=>0�=�a�=n#�=���=�.�=���=z:�=pg�=�Aq=�`=��X=(&\=0�i=�
�= ��=�`�=�=H?�=���=�   �   � �=[��=�P�=�<�=ȉz=��<��c��������|�-F��:n���%�s[L��q��+��?���<����pS���&���H��_�q��,L��%�%��󮸾�,y����*T����*�H�=@��=V�=��=�=T��=Q��=}�=���=ME�=�0l=,
F=�^'=��=�c
=�=�$=:{:=<%^=�x�=���=�b�=л�=�   �   ,޲=�=�C�=��=�/�=vD=�͟���r� [���`����P����:�Q']���{�iΉ��|��6/��У������7|���]�A�:�y���������S^���|�g�����=�8�=�Q�=x޽=���=���=r&�=^g�=��q=�9=��=č�<0�"<@(e; mi: \;PW�;���<Ll�<��'=��_=d��=H�=�   �   Е=�=��=��=�>�=&9*=@��;�M+��3׽�=��ȏ���Ⱦޟ���#�"C�ԟ^��Pt��!������X���u���_���C���$����ɾ2���� <��;Խ��#���<�3=�e�=_��=�i�=ݔ�=>��=nB�=��G=���<�qG< �Ļ�5��B;�DX3�JA��8�d��<�Ӽȍ(��2�;L5�<L5=D"w=�   �   (�^=�I�=4J�=��=�g�=��E=��<�ƴ�Q�!���j�uF���jܾ�D
��i%���=�	�P�C�\��Ea��`]��Q�z�>���&��W�z޾�p���]k��T��Y���孼���<��L=[��=� �=��=P'�=h�n=$=���<P�Ի��4�g�����Ž��ܽR�|�t,˽�q��p�{���XQ?�(�V<P�=�   �   (O�<�Q=�N�=LՏ=���=>t`=F�= �ƺ>C@�p(ֽv2�d~���㯾c
߾cf������*�Cr5��A9��6�D,��"�
�����9��R��@5�'hٽvhC� gҺ��=z�d=���=#�=��= �^=��=`�<�$���]��´��������LA3��<C��]I��E���6�4������g����s�8JռG�;�   �   `�;���<\R=�ˁ=iN�=�aw=tM6=�ʗ<L䑼�0��RW��EF?�>����⪾5/о'����W������>����Y��KӾ�򭾜I���C�����j^��Tq��pl�<�G5=ƾx=w#�=�ӄ=��Z=z�	=�y�;t��Ƌ�5��/e!�έN�b<w��΋��i��\k��*o��a���jn|��T���'��|�&v���-��   �   p���В�;�W="�_=�ރ=
y�=�c=��=�Z<4$߼2���o����"9���u�^N��a���ƻǾSyվ%�ھ�־{�ɾ�u��p��
|�5?����X��q�����;\=b�_="߃=vx�=�c=��=><�7߼���������'9���u��Q��>����Ǿ�}վ��ھD�־��ɾ�y��Ts���|��?�<�)	���   �   "c���~��`c�<HE5=�x=�#�=�Ԅ=��Z=��	=���;X��������`!��N��5w�'ˋ�f���g��vk��޶���g|�`�T�є'�mt�o��~#� ;���<�	R=�́=yN�=�_w=J6=���<���:6��a^���J?����H檾3оs��*�Ŭ����HA�(��]���NӾ����,L���C������   �   mٽpoC���Һ��=Hd=б�=�=���=(�^=�=x<l��~]�����0���@��v;3��6C�NWI�pE�3�6���I��]_��V�s�44ռ���;<\�<��Q=qP�=�Տ=k��=Zr`=��=��Ǻ�K@�".ֽ�y2�ˀ���毾�߾mh����H�*��t5�>D9�16��,��$��������;��BT���5��   �   W��\����<8�L=]��=��=*!�=j)�=0�n=�$=���<p�Ի�����g����nŽ��ܽ����߽W#˽\i��l�{����%?���V<h�=v�^=�K�=VK�=��=Sg�=t�E=��<�Ҵ�������sj��H���mܾxF
��k%�و=�t�P���\�RHa�_c]�2�Q���>�՞&�*Y�޾�r��ak��   �   $#<��>Խ��#�8�<��3=�e�=���=�j�=|��=��=XE�=�G=�<КG<@gĻ���F-��I3�B;A���8�����qӼ�_(�Ѓ�;XF�<P5=�'w=ҕ=f��=� �=��=|>�=7*=��;8S+��7׽�=��ʏ��ȾB����#�C��^��Rt�#��A���Z���u���_���C�l�$���ɾ�����   �   �U^���ʑg� ���=�8�=R�=4߽=��=���=�(�=j�=�q=9=z�=`��<H�"<@�e; l: ;���;,ӆ<�|�<��'=�_=���=S�=�߲=�=bD�=��=b/�=�B=�矻��r��\���`�����R���}�:��(]�e�{�Wω��}��*0���������h9|�\�]�s�:�t����5����   �   .y�V��?U����*���=0��=��= �=��=b��=���=�~�=���=�G�=6l=&F=Le'=j�=~j
=̢=+=*�:=�*^=�z�=���=�d�=$��=�!�=��=$Q�=�<�=��z=x�<�c�쪕���ָ|�[G���o���%��\L�F�q�},�����K=�����T��F'��I��X�q�_-L�M%�&�������   �   +���@"�8E���l�� A�<��=��=���=�0�=:b�="$�=���=�/�=2��=�;�=�h�=$Eq=�`=,�X=|)\=R�i=V�=J��=�a�=��=@�=D��=`�=�"�= ��=&,�=t�t=@�<f��������&�\���Lƾ�r�/���W�ט~�te��0ʝ��Y���O���c��՝�b��z\~�c:W�W.� ���6ľ�   �   F��4{&����$����j�<)��=iu�=dR�=Z��=�F�="H�=�i�=��= ��=Pz�=`��=�Ä=py=`�r=�u=��=
}�=]�=0��=�e�=��=���=L	�=���=m]�=�j�=��r=(f�<�����쭽�+��u��Bqʾ�
�\2��[�ƈ��O���u��>"��e!��(��8w��ђ��\��[�s�1�4	��-Ⱦ�   �   J*���?"��C���h���C�<���=6 �=���=�0�=Lb�=4$�=���=�/�=/��=�;�=�h�=Eq=�`=�X=^)\=8�i=J�=C��=�a�=��=@�=N��=y�=�"�=@��=�,�=��t=t"�<la��ﴧ�v�&�@[���KƾIr�D/���W���~��d���ɝ��X��>O��Pc��nԝ�ua��g[~�t9W�NV.����6ľ�   �   O+y�N��XR���*�f�=��=,�=� �=�=���=đ�=�~�=���=�G�=�5l=F=&e'=D�=Rj
=��=�*=�:=|*^=�z�=���=�d�=6��="�=F��=�Q�=�=�=�z=��<��c�ϧ�����޵|�aE��,m��c�%��ZL�$�q�O+������;��m���R��&���G��I�q��+L��%��#��㭸��   �   �Q^�K����g�@]�� = :�=�R�=�߽=t��=ˊ�=�(�=j�=�q=�9=L�=���<p�"<`�e; l:`�;P��;�҆<�|�<��'=��_=�=h�=�߲=t�=E�=��=�0�=�F= ���.�r��Y��`�熧��N����:��%]��{��͉��{��O.��ꢑ���26|�|�]���:�b����澡����   �   �<�78Խ�#���<h�3=�g�==�k�=疭=���=rE�=�G=�<��G<@iĻD���-�J3��;A���8����hrӼa(�P��;�E�<>5=�'w=Nҕ=Ћ�=�!�=��=5@�=&<*=���;�H+��0׽�=�qǏ�غȾ���k�#�wC���^��Nt�� ������W��pu���_�
�C�o�$����ɾ�����   �   R�}U��X٭���<|�L=(��=��=�!�=�)�=��n=�$=���< �Ի����g�%���Ž�ܽ��*�߽�#˽�i��ڢ{� �x&?�x�V<��=�^=L�=L�=3�=6i�=�E=(�<໴��윽���sj�_D��Chܾ C
��g%���=�ʎP���\�aCa��^]��}Q�\�>��&��U��޾�n��bZk��   �   �bٽ@`C�@�Ѻ��=��d=���=I�=~��=�^=��= <d���]�����Z���^���;3��6C�xWI��E�`�6���q���_����s��4ռ���;�\�<��Q=<Q�=:׏=Z��=x`=�=�?ƺ�;@�e#ֽ�r2�F|���௾0߾�d������*��o5�6?9�@6���+�� ���<��S6���O���5��   �   :Y��Ha���x�<�L5=>�x=�%�=�Մ=,�Z=|�	=���;��������)`!��N��5w�<ˋ�3f���g���k������5h|���T� �'��t��o���#��;��<^R=�́=VP�=�ew=R6=L֗<TՑ��+���P��4B?������ߪ��+о!�����"���<���vU��mGӾ�ﭾ�F����C��z���   �   �]�� �;b=L�_=\�=�z�=6�c=��=p]<�#߼(���{����"9�αu�nN��x���߻ǾpyվE�ھ�־��ɾv��'p��[
|�c?����~���p�����;^]=��_=���={�=��c= �=�v<�߼X������9�2�u�'K������ѷǾ&uվ�ھ��־x�ɾ+r���l��q|�w?����4����   �   ��;$��<fR=�΁=�P�=�dw=PO6=�̗<(㑼�0��SW��NF?�J���㪾I/о?����i������>����Y��>KӾ�򭾹I��-�C�Ӂ��n^���p��tn�<�I5=��x=�%�=�ք=��Z=�	=p��;��缠������W[!�d�N��/w��ǋ��b���c���g��n����a|���T��'�6l��h�����   �   �j�<��Q=�R�=؏=z��=�v`=�=��ƺ�B@�a(ֽv2�l~���㯾u
߾nf������*�Vr5��A9��6�\,��"� �����;9��9R��_5�>hٽ8hC��LҺ�=�d=���=�=��=��^=�=�3<����8�\��������"���53��0C�SQI��E���6�������>W����s�|ռ֗;�   �   ��^=N�=rM�=��=3i�=��E="�<tŴ�'����j�}F���jܾ�D
��i%���=��P�X�\��Ea�a]��Q���>��&��W��޾�p��
^k��T�sY��\䭼��<��L=���=A�=#�=�+�= �n=�%$=(��<�-Ի��Z�g�����
Ž��ܽ$潗�߽l˽a����{�����>� W<��=�   �   �ԕ=l��=~"�=T�=@�=�:*= ��;M+��3׽=��ȏ�ǼȾ����#�.C��^��Pt�"��&���Y���u���_���C��$����ɾG���!<��;Խ>�#��<��3=<g�=8��=rl�=S��=Ĵ�=)H�=��G=� �<��G<�Ļ�����;3��,A�n�8� ��`XӼ�1(� ��;�W�<�"5=�-w=�   �   ��=��=�E�=,�=�0�=�E=�ȟ���r�[���`����P����:�\']���{�qΉ��|��@/��ݣ������7|�
�]�V�:����������T^���6�g����=�9�=S�=V�=x �=J��=�*�=�l�=�q=9=l�=��<��"<�of;��n: �;@��;P�<t��<<�'=Z�_=���=��=�   �   *#�=
��=R�=�=�=��z=
�<0�c�𨕽����|�2F��@n���%�y[L��q��+��E���<����yS���&���H��p�q��,L��%�%������,y����T���*���=���=6�=� �=��=���=��=k��=���=�I�=8;l=�F=nk'=��=q
=@�=L1=�:=�/^=@}�=���=\f�=���=�   �    �=B#�=���=�,�=��t="�<Pb��Z���ş&�|[��(Lƾ�r��/���W�.�~�e���ɝ�<Y���O���c���ԝ��a��\~�:W��V.����6ľ�*��V@"��D��xk��B�<L��=( �=��=1�=�b�=�$�=���=�0�=L��==�=Pj�= Hq=`=X�X=�,\=^�i=��=���=�b�=��=�@�=��=�   �   ���=���=˱=��=Fy$=��<�����W�Z���cȾ&���?�Kzt�n��9���_�Ŀ�ֿ`�῅�忁��s�ֿ��Ŀ�V��{����Js�O<>�]O��ž��~��o��`r� ��:h3=�f�=�~�=$��=���=���=֞�=V�=$�=i�=�a=NDD=H�0=)=�-=&�<=�zV=��w=\�=�p�=k.�=
��=�   �   �=m��=��=(<�=r.'=@0��2]y� @��L~��BľH��T<�s*p�ې������|���ӿJ(޿E ⿀4޿�ӿ����儫�1��� o���:�t�
�J���7>y�&���Rh�`� ;
~5=��=죶=OX�=�$�=���=���=�2�=`̊=k=h�D=��%=��=\=P�="�=��9=�]=�u�=���=���=2+�=�   �   iD�=zf�=fV�=�(�=��.=��K;nPZ�F`�8m��H��~ ���1�k�c��+���J�� q��Sɿ��ӿ_W׿q�ӿ�/ɿZ����K����� c��0����~&���h� U��,K�p��;`<=\��= �=&B�=ć�=�)�=D�==ҍP=Z=���<lv�<�:<�&<8�(<�|<\��<�=|�@=� u=�1�=ns�=�   �   ��=0 �=nm�=ࢉ=H�8=h!<R3*���彠AR�W������!�P��%�w��+ǩ�<���%ÿ��ƿ\ÿv����%���T��`h�!�O�ۉ!�}��;��"7O�:�߽���WQ<��D=�Ï=6�=��=U��=.�=ڂc=�� =�W�<���;h=#����`7���%�J> ��Nȼ��Y����:4��<f�=&�Q=��=�   �   8hm=ͯ�=|s�=䲄=��C=`~�<t�ۼ��G0�� ���{ϾG��� 7��~a���Q����������<���S��V���Ւ��=����Xb���7�%���RϾ�p����.��貽��ɼ8��<��M=<G�=Ԩ�=f��=�H}=�4==���< �k;@Ӥ�>�0� ǂ�M����ẽ�ýJ载3Y��������C��mͼ�6���$�<6m+=�   �   ��=�ES=hy=r�x=�(L=���<�+��Z���
�N�f�G諾hj�
����?�gc�6t��؍��ҕ�����o-���w��58���d��A�`�����𧬾�Mg�x�	�c����{�<D�<�_T=�8�= f�=1a=�%=PLy<@�S���5��ǝ���޽4��F�#��W3�?9��"5��e'��R���齻]���iL�D����L-<�   �   �-�; ��<4B=$=_=��O=�;=���;r��Ľ2�/�s��rս��0��L`�g�:�8sU���j��Yx��T}��y�Gl�5+W�l<�\�������U����1�'tƽ������;�==\�U=xgg=��L=2�	=�<��ż�ր���ؽ��@�F���n�1J��Ǒ������Ւ�aH��Yt�,�L��� ��H�)I������   �   �5��]�;P��<��;=�WL=TE,=��< �:�F�n����YF�����}���	�� ��T�(��:��uE���I�J3F�Fr;�MV*��k�9���þ6<��skJ�s����0v�&K��w�<�-=T
P=�4B=�P=p��;k�� ������>:��w���������r�ɾ& ؾ9BݾN9پLC̾)���`3����~��@�JO�}���   �   
���MԼP�+<h�=��@=�;B=�=�G<<z���ΐ�4D��J�Ȉ��&���)�ھ���K������L�۝�v�u� ���޾�j���􎾝�O����t���=Լ ,<@�=X�@=b:B=J�= �G<����Ր�^H��J���������ھ7���������O����.�� �D�޾kn��������O�f 	��   �   �����9v�@=K��p�<ʐ-=8P=�7B=*V=��;TU伙��ӳ��
9:�*�w����8�����ɾ0�׾0=ݾ`4پ�>̾㗷��/��=�~���@�K�����+��;T��<�;=XL=\C,=�ز<;�v�n�����]F�����0���u�󾭄�+�(� :��xE�7�I�s6F�Eu;�	Y*� n�>=��z�þ�>���oJ��   �   P�1��xƽ�����;:<=ĺU=�ig=ֽL=��	=` <0�żπ�}�ؽ8��F�h�n�TF��Ñ������ђ��D��\ t���L�B� ��?�B���z��o�;���<�!B=�>_=N�O=�9=�f�;��d�Ľ�/�����ؽ��4���b��:�3vU���j�]x��W}��y�al�.W��n<���������������   �   �Pg���	�a���x���@�<�_T=�9�=�g�=\6a=�,=`ry<P�S��5�:�����޽���:�#�tQ3��89��5��_'�-M���DU���[L�xn���p-<R�=>JS=8y=~�x=(L=P��<��+��^��|
��f��꫾�m����?��ic��u���ٍ��ԕ�T���/��zy���9��}�d��A� ���������   �   `r����.�4벽��ɼ얦<��M=�G�=��=c��=�N}=�;==P
�<�Fl;����&�0�����=���xغ�ߎý�޽�8P��5����C��Sͼ�۳��6�<,t+=`mm=���=�t�=-��=��C=�x�<��ۼs�RJ0����O~Ͼȝ�z7��a�Y��������)	��l>��U���������Y����Zb���7�i���TϾ�   �   �<���8O�`�߽����QQ<B�D=ď=�=���=X��=�0�=��c=�� =lj�< �;�#�h���������0 �5ȼX�Y�@ݙ:�Ґ<<�=��Q=E��=�
�=s�=n�=�=(�8=h� <�7*�����CR�䡥���h�!��P��'����Mȩ�S=��7'ÿ��ƿ�]ÿ�����&��hU���i�k�O��!����   �   C'���h��U��.K���;,<=���=��=C�=��=j+�=:F�=�Ă=�P=a=��<І�<p�:<XI<x�(<`�|<|��<��=��@=�%u=�3�=u�=�E�=Kg�=�V�=�(�=��.=�qK;�SZ��a��m��I��F���1���c��,��nK���q��3ɿ|�ӿBX׿L�ӿ�0ɿ���*L��y��� c���0����   �   �����>y�h��6Sh�`� ;~5=��=C��=�X�=�%�=v��=���=4�=�͊=xk="�D=�%=��=X`=~�=�=H�9=\�]=7w�=Ȑ�=� �=�+�=��=���=/��=<�=�-'=@[��V_y��@��M~�XCľ����<�"+p�@�����������ӿ�(޿� ��4޿ӿ���1���U1��L!o��:���
��   �   �žx�~��o�@`r�@˅:�3=�f�=�~�=<��=���=���=䞻=f�=$�=i�=�a=dDD=Z�0=$)=�-=�<=�zV=��w=Y�=~p�=_.�=���=���=p��=�ʱ=߅�=�x$=`�<�Z��X�����cȾG��)�?�rzt����K���m�Ŀ�ֿg�῅��}��j�ֿ��Ŀ�V��k���uJs�0<>�@O��   �   ����5=y�i��tPh��!;X5=`�=���=�X�=�%�=���=���=4�=�͊=xk=*�D=��%=��=D`=b�=��=8�9=T�]=6w�=͐�=� �=,�=��=��=t��=�<�=/'= ��^\y��?�]L~�KBľ��<�*p�����L���%����ӿ�'޿���4޿EӿK��������0��F o�5�:��
��   �   e%��b�h��S�H)K�  �;�<=p��=�=oC�=H��=�+�=QF�=�Ă=��P=a=���<���<��:<�H<��(<��|<0��<��=n�@=�%u=�3�=&u�=�E�=�g�=WW�=d)�=>�.=��K;NZ�x_�m��G�����0�1���c�e+��J��mp���ɿơӿ�V׿��ӿ/ɿ�����J��O���b�,�0�@���   �   -:���4O��߽4���eQ<��D=:ŏ=��= ��=���=�0�=��c=�� =pj�<�;8#���������&1 ��5ȼP�Y�@י:xҐ<,�=��Q=^��=�=��=�n�=&��=��8=�!<�/*�6���?R�'������!�� P�+$����)Ʃ�;���$ÿU�ƿT[ÿU���s$���S���f���O���!�����   �   Ho���.��䲽��ɼ��<��M=,I�=���=괒=O}=0<==�
�<�Gl;���D�0�����X����غ��ý߽�dP��`���N�C�TTͼ@߳��6�<bt+=�mm=��=iu�=���=ڹC=셓<�ۼ�붽�E0�Y����yϾ���6��|a������K��F���;��BR��������������Vb�C�7�����PϾ�   �   5Jg�̳	�i����c�DN�<|dT=D;�=�h�=�7a=�-=�sy<��S��5�C�����޽���O�#��Q3��89��5��_'�IM�M��rU���[L��n���q-<�=`KS=*!y=��x=�,L=���<x�+�9W��]
��f� 櫾�g�L����?��dc��r���֍�cѕ�����+��wv���6����d�sA����������   �   ��1��nƽ̊����;"C=l�U=�lg=̿L=��	=�<��żπ�~�ؽD��F�~�n�`F��Ñ������ђ��D��� t��L�d� �#@�B���z��s�;���<�#B=�A_=$�O=�@=��;
���Ľ�/�B���ҽ�g-��(^��:�npU���j��Vx�XQ}�my�3�k�X(W��i<� �N������������   �   ����`&v�K�p��<��-=�P=�:B=�W= '�;@T�{��ͳ��9:�4�w����G�����ɾE�׾H=ݾz4پ�>̾�����/��h�~���@�K�����+�Н�;���<<=�\L=\J,=<�<��:���n�����TF�뎏���������(�:��rE�ٞI�10F�No;��S*�i��4����þ\9���fJ��   �   ,��� *Լ�+,<��=��@=@B=��=��G<tx���ΐ�(D��J�Έ��0���7�ھ*���W�����M������� ���޾�j���􎾼�O����\��<Լ�,<��=��@=�@B=��=�G<,h���Ȑ�]@��J�����u�����ھ:��������J�
������ �m�޾�f��]�t�O�����   �   � �pے;8��<�<=�]L=I,=8�<��:���n����YF�����������(��^�(��:��uE��I�^3F�[r;�`V*��k�:9��,�þL<���kJ�o���:0v�� K�L|�<��-=P=�<B=�\=0_�;l@����V����3:�ԍw�\������#�ɾ_�׾E8ݾ�/پ :̾�����+����~�F�@��F�����   �   �;���< (B=D_=x�O=*?=���;X���Ľ&�/�t��wս��0��S`�q�:�DsU���j��Yx��T}��y�`l�M+W�.l<�o�-������d���"�1��sƽ������;�@=8�U=�ng=��L=��	=�#<��żȀ�Šؽ�ԜF���n��B����������͒��@��]�s���L�ߑ ��6彚:���b��   �   �=�PS=z$y=,�x=�,L=د�<��+�UZ���
�H�f�K諾pj���ɽ?�!gc�<t��؍��ҕ�����|-��x��B8�� �d��A�s��	������Mg�n�	�����u�TI�<�cT=�;�=2j�=*<a=@4=(�y<�|S��r5�����/�޽B��c�#�MK3�^29�s5��Y'��G�C�齸L��ML�pV����-<�   �   �sm="��=�v�='��=��C=\��<�ۼ��G0�� ���{ϾK��� 7��~a�$��Y����������<���S��c���咗�J����Xb��7�6��SϾ�p����.�C貽��ɼ��<��M=xI�=���=���=,T}=C==��<@�l;ԟ����0�����x���CϺ�{�ý�ս�PG�������C��9ͼ@w��,I�<�{+=�   �   $�=^�=�o�=���=��8=!<�2*�w�彔AR�X�����!�!�P��%�{��2ǩ�'<��&ÿ��ƿ�\ÿ�����%���T��vh�3�O��!����;��"7O�
�߽���\Q<��D=Vŏ=��=?��=t��=^3�=�c=�� =||�< g�;��"��u������
��# ��ȼXtY� 3�:��<N�=N�Q=�=�   �   .G�=�h�=�W�=�)�=�.=��K;�OZ�4`�3m��H��� ���1�p�c��+���J��%q��Yɿ��ӿhW׿{�ӿ�/ɿe����K�����* c��0�����&���h�U�L,K�0��;�<=p��=��=0D�=x��=-�=PH�=:ǂ=��P=�g=���<���<X ;<k<� )<��|<���<��=��@=+u= 6�=�v�=�   �   v�=p��=���=�<�=(/'= #���\y�@��L~��BľJ��V<�u*p�ܐ���������ӿO(޿K ⿇4޿�ӿ����鄫�1��� o���:�y�
�N���:>y� ��fRh�`� ;�~5=L�=���=XY�=<&�=D��=���=N5�=Kϊ=�
k=��D=̖%=��=fd=��=��=��9=��]=�x�=��=��=�,�=�   �   *-�=��=��=�^=H{�<r��Q��P8]��˵�~�ɭ>�V�|�H���#l��9o�i���j
�(l�����m��
�������\����ힿn{���<��y��ײ��X���ڽ0x��4״<b�k=)�=��=�l�=(=�=LQ�=��=��r=�C=�=|��<h��<S�<���<�]�<V�=�j7=�Ke=`�=�w�=���=�   �   �@�=��=���=TV^=�H�<���\�ܽ��W� ����v�v(;�V[x�k���:����ݿa���,��������p�����yqݿ%����P����v�n�9����/���	S�h@Խ�XＤ	�<�j=l��=\ �=���=�{�=��=�*�=Z�V=(�#=���<�ѡ<��a<8�:<��Q<���<�{�<�!=V�H=8 |=�~�=�ç=�   �   �@�=���=,��=��[=��<�d߼Sɽ��H��⦾�����0��bk�O!����|'ӿ^��8h�:9�ƞ
�HN�L��_��,ӿ�������Dj�r�/�Z��v���$�D�2y��0+ļ��<��g=��=2��=��=s�=x�}=�B=��=��< �;��\����i������ �0� ��X�Q<���<f_2=�[n=�=�   �   ���=���=���=4V=��<|ڙ����1�������G� �2W�����Hb����¿�Aۿ����P�����������5�e�ۿr�¿a��������V�(F ��������-��i�� ͂�$��<�Ga=^ߌ="�=O��=@,]=̎=\t�<@q����˼��1���n�$g���4����޳x�x�?��o�ء
�@�O<��=T�M=�   �   �(=�[=Էi=&rJ=�'�<��
�W��<+���Iž���H7=��q�����A����ÿ�@տ�࿞�� �2�տ�qĿ�����C���vr�j=����tľJ�}�@$�<����ͻ !�<��T=�5u=2�h=�+7=8A�< �D:T� �h��\��@+体/�V�Tf�����1
�oi콚����}����0׀����<�   �    �C<$=��6=�Y6=8��<��;�]4����B�N��ᢾ������v�M�.�|�픿����Y7���7¿#�ſ��¿�	������_啿��~�YO�� ��w�v&��RN����Z/�`�;�=$y?=F�A=�=��<�T��E��L�����`	-���Q��o��v��%��ro���0s�N�V���2��	�v��|�Z��㏼�   �   ��ͼP�;���<m=�:=0Q<�7��L㞽����~�/���^��(��P�(ev�q#��Fy��2���6������W��L7���x��
R���)�֗��ٽ�ƀ��>���P��(�� �_<>�	=�'=�C�<��(<����p`~�kj��x)��c��T��৾EK��(�ɾرξ��ʾ ����ت�2���8�j�� 0�`RｙS���   �   ����\�ͼ ��;��<�. =��<@�n� �9�ֽa:�J!���AǾ�$���#�LsC���_���u�������v���tbw���a�H�E�d�%��	<ʾ�[���}=�k�ٽ��=� ׂ���<�=�$�<�<��I������ƫA�E����߭�MFԾڱ���	�]	�"_�V���b
�-��Q.ؾ�ͱ�=(��6H����   �   )a���u��TW��8�N<$��<`�<��^<X6��x"x������G�����¾ü������\*�6(<�һG��L���H��=��U,�  ������ž�ɓ���L�Z���p��HJ��xO<���<d\�<@�^<�E���-x�|���ڽG�����#¾�������`*��+<���G��L�3�H�g�=�'Y,��"�������ž"͓���L��   �   ��=��ڽ&�=� ���<��<��=0,�<�/<pߴ�C��yy����A����nۭ�IAԾ9����	�,��[�+���_
��'��t)ؾ�ɱ��$����G����g{���ͼ���;@�<�. =��< Jo�Ɨ9�zֽ�e:�E$���EǾF'�q�#��vC�.�_���u�������u���>fw�+�a�`�E�&�M��?ʾu^���   �   ւ��%�mT��D��X�_<��	=�*=dN�<H�(<4����Q~��`�s)��c�vP��|ۧ�KF���ɾ��ξg�ʾ}��tԪ�8���f�j��0�aI｣L���ͼ J�;���<o=�:=0Q<�C��螽u�m �62���`�](��
P��hv�R%��G{��H��	9�������X��9��7�x�ZR���)����Vܽ��   �   }(���TN����r_/��;�=8{?=j�A=6�=
�<x�S��E�OC��7��-���Q�Zo��r��� ��fk���(s�F�V���2���	����0�Z��͏�0�C<�)=��6=�Z6=X��< �;�c4����N��㢾ڤ������M� �|������P9���9¿0�ſ��¿���m����敿>�~��O��� �~z��   �   �vľ��}��%�Z����ͻ� �<�T=�8u=�h=�27=TS�<�[G:p�j�h�\S��� ��)�L�6`����,
��^�E��\u}�"t���� ɭ<�(=8�[=B�i=�rJ=d%�<@�Z���-�Z���ž5��49=�m�q�e���{C��L�ÿwBտ���}������տsĿC���)E���xr��k=�O���   �   �������{�-��k���Ђ�`��<�Ha=p��=��=ė�=�2]=��=,��<`����˼��1�|�n��^��j,�������x���?�XU켸s
�%P<��=��M=ڄ�=z��=P��=\V=��<����Ɓ���
1�!���Ձ㾗� ��W�����nc����¿Cۿ}��UR��2������7￮�ۿ��¿Z���箈���V�*G ��   �   Y��%����D�Rz��x-ļX�<r�g=��=\��=N�=��=Ē}="
B=�=�<��;�������4T��pr����0� ���Q<d��<�e2=�`n=�ď=fB�=�¡=���=��[=�<�i߼iɽA�H��㦾������0�0dk�"����s(ӿl���h��9�Z�
��N�΅�F���ӿc�������cEj��/��   �   M��.0��.
S��@Խ�Y＜	�<��j=׼�=� �=V��=�|�=T��=�,�=�V=Z�#=��<�ۡ<p�a<0�:<��Q<���<���<�%=��H=4|=��=�ħ=fA�=@�=⾙=V^=�F�<v����ܽ~�W����� w�);�\x����7;��o�ݿ����z���V��(���������qݿs����P����v���9��   �   �y��ײ�;X���ڽ�v��ش<Ăk=P�=��=�l�=@=�=\Q�=��=��r=(�C==���<���<$S�<���<`]�<D�=�j7=�Ke=S�=�w�=���=-�=��=��=��^=,z�<&��ϱ㽦8]�&̵����>���|�_���;l��Po�{���p
�,l�����m��
�������G����ힿD{���<��   �   ���B/���S�?Խ�T���<��j=.��=2!�=y��=�|�=]��=�,�=�V=d�#=(��<�ۡ<8�a<�:<H�Q<h��<p��<�%=��H=<|=��=�ħ=�A�=x�=<��="W^=,J�<����ܽ"�W�����Tv�.(;��Zx�-��i:����ݿ������r������&�������pݿ����DP����v�ފ9��   �   ���d����~D��v��`$ļX$�<v�g=5�=���=��=��=��}=@
B=�= �<��; �����dT���r���0� ����Q<P��<�e2=�`n=ŏ=�B�=�¡=M��=��[=x"�<`߼�
ɽ��H�%⦾�����0�bk�� ��񴿳&ӿy��g��8�:�
��M�Ƅ�c��Gӿ��c���YCj���/��   �   *��h����-��f���Â����<^Ka=X�=r�=��=$3]=<�=���< ����˼��1���n��^��},�������x�ܧ?��U�t
� %P<��=֏M=,��=��=C��=LV=��<hә��|��1�����N~�@� ��W�ӿ��Oa��r�¿Q@ۿ���HO��������64��ۿ:�¿N���*���%�V��D ��   �   �rľ�}��!�� ����ͻ�*�<j�T=;u=r�h=j37=@T�<�jG:(�h�h�`S��� ��)�Y�E`����,
�_�^���u}�,t� ���ɭ<�(=��[=z�i=BvJ=0�<8�
�*T��B)�J��hžl���5=��q�Խ���@���ÿ�>տ��Τ�Q��z�տ�oĿj����B���tr�@h=�����   �   #$���NN����.S/�0%�;f =�~?=��A=��=��<��S�rE�@C��6��-���Q�go��r��!��qk���(s�\�V���2���	���� �Z� ͏�H�C<>+=^�6=�^6=��<�1;W4�P��8�N�tߢ�ٞ�
��<�M���|��딿񯨿5���5¿&�ſ��¿��ꬩ��㕿��~��O� � ��t��   �   q~�����dK��,�����_<l�	=D.=S�<��(<�~��Q~��`�s)�	�c�wP���ۧ�TF����ɾ��ξv�ʾ'}���Ԫ�F�����j��0�gIｅL����ͼ U�;���<�r=h@=�.Q<�)���ޞ����d�~�/,���\��(�(P��av��!��\w��/���4������U��z5����x��R�H�)�ߕ�vֽ��   �   [y=���ٽ��=� ����̲<��=\3�<�8<�ܴ��B��Ly���A����oۭ�NAԾC����	�3��[�6���_
��'���)ؾ�ɱ��$����G����${����ͼp��;�!�<f4 =D��<`�n�څ9���ս]:����5>Ǿ�"���#�>pC�#�_���u��	�����|���^w�(�a��E���%����P8ʾ�X���   �   �Q��}j��P7��P%O<���<,j�<��^<T2��^!x�;���z�G�����¾ʼ������\*�>(<�ݻG��L���H���=�V,�. ������žʓ���L��Y��!p��`F���O<4��<8l�<��^< %��2x������G�𔐾�¾�������Y*��$<�:�G��K��H�v�=��R,�=������ž�Ɠ���L��   �   bt��$�ͼ���;�(�<h5 =��<��n�J�9��ֽ�`:�E!���AǾ�$���#�RsC���_���u����
�������bw�§a�Y�E�s�%�(�<ʾ�[���}=��ٽ6�=�@���8Ȳ<�=9�<�O<`˴�|<���p����A�F|��T׭�~<ԾѦ���	���X����\
��!���$ؾyű�D!���G�R���   �   <�ͼ@��;��<�u=�@=�&Q<�2���➽�����~�/���^��(��P�/ev�w#��Ly��:���6������W��W7���x��
R�Ľ)����ٽ�Ȁ�����O�����8�_<�	=\0= \�<�)<j��TC~��W�tm)�R�c��L��ק�tA��ӡɾU�ξ@�ʾ*x���Ϫ�,���p�j�0��?�E���   �   �C<�1=r�6=�`6=��<�;�[4�;��$�N��ᢾ������{�M�4�|�픿����`7���7¿/�ſ°¿
������l啿��~�jO�� ��w�~&��RN����Y/���;�=(�?=(�A=Z�=�<��S�Z�D�{:�������,���Q��wo��n�����bg��<!s�1�V�b�2�G�	�U����Z�@����   �   �(=x�[=|�i=�wJ=\/�<(�
�`V��+���Gž���M7=��q�
����A����ÿ�@տ�࿪��+ �A�տ�qĿ����D���vr�j=����tľE�}�$������ͻ�(�<�T=�=u=��h=�97=�d�<�J:��߼��h�,J��L�4$�d�.Z����X&
�`T������d}�f��"��ܭ<�   �   ���=ԣ�=Y �=,V=8��<י��~���1�������H� �5W�����Kb����¿�Aۿ���P�����������5�s�ۿ~�¿l��� �����V�0F ���������-�}i���ɂ�h��<�Ka=&�=��=X��=.9]=�=t��<���ԙ˼"�1�Ȝn�uV���#��^��x�Ԙ?��:켠D
�8MP<�=r�M=�   �   ED�=ġ=��=B�[="�<�b߼ɽ��H��⦾
�����0��bk�Q!����'ӿc��<h�@9�̞
�NN�R��j��5ӿð������Dj�x�/�c��w����D��x��$)ļ8"�<X�g=��=���=��=��=ؗ}=BB=F�=�$�<� ;��(|��?��h]��0�0��, �hR<|��<"l2=>fn=2Ǐ=�   �   aB�=�=���=�W^=XJ�<B��:�ܽv�W�����v�w(;�X[x�m���:����ݿc���.����
����r�� ���qݿ+����P����v�r�9����/���	S�I@Խ�W�8�<b�j=R��=�!�=��=�}�=���=.�=��V=T�#=��<h�<`�a<��:<�R<h��<���<4*=��H=l|=y��=Ƨ=�   �   �:�=��=G��=�= E��A��`'�c�����/���r�^r���ȿ+��l��g��-���6��W:���6��-��:���B�%�ƿ�^��n�p��-�n��ₓ���"���� P���D)=⁉=��=<[�=���=�P�=��l=�5=0��<d��<X6<��%; �8�P�:��;T�<���<�.)=�`=�x�=�}�=�   �   08�=LO�=��=�+=`R����T�"��͒�����:,�4�n�%���d�Ŀ�<� 
�����#*��3�T7�X�3��$*�r����	��z��ÿ����e�l��*��x]��b��ua�� �й�q(=��=�B�=�w�=`Ř=0��=�<P=t�=� �<�Z<��`�� D��&�L��Pz�;$,�<�(=��C=>0{=��=�   �   ��=\Ƌ=�%t=�q= �ƹt�u�:��oP���ܾ	�"���a�͔�1������^+���!�j�*�R�-���*���!��@��s��z�م�������`�0W!��پ�=����"�i� �;ba%=�}=�=�z�=�ly=�&@=@��<4<���ü0P���:�6YH���>�4L���ؼ�g,�>�;���<��2=m=�   �   �H=fe=��W=��=�l;�>K�x���+u�Κƾ���i@N�b������п�o���x��T��v�����������n2п�竿���wM����'�ľdr��� �A�@��;x<=��a=jBp=��T=�=pR�<@������k��F��h�ǽ�߽����Y�̽͡qީ�2�z��l�н3��0Y<�(=�   �   ��<��=4�,=a= ��;zx�7Tؽ�P��n��A� ��25�Sq����M^��.fؿ�����V���f����7�����EEٿ9�������@q��5��� ������9N�rԽ���x> <=(�6=^\'=�;�<��D;��ۼ��y�mPƽ��`J'��	A���Q��MX���S�y	D��\+����+Fн	��� ����~a��   �   h�E���_<`��<�{�<(�6<����$�����&�$���n-׾�����L�8����t���ɺ���ҿ����
�I�������Կ�����j���j����M�'P�}׾�����&�{b��Ӷ��P<�F�<���<<�<�
�D2����t�	�~�=�:�p�����U���C���'E���7��,���4yv�"�C�~��(_����C��   �   �i��s�����;�ƕ<@�N<��4���`�8���0[�&��@����:'��W�P��~������R��.�ʿ#�οog˿�b��h���̜��8����X�V�(� ����:��XI\�m����_��(� .b<Ą�<�"<�s��Y���ӽ �'���l�Mv���ý��qݾ����П�$��^A��������J�����_s�I�-��ݽ�   �   ���|zi�h䎼�`�;h�;< ~Ź P���������|���%|��DR�v)���Q�|�x�=������:գ�u	���a�����ǎ�S{��ET�F~+����ӿ��*��� ��@���� � (@�� H<0��;(�{�Ƅ]��޽^c6�|P��6,��I"�Qj
����U�0�ҿ;���?���<�@%2���!�����F�Y�<���p�;��   �   �7��EԽ�.D�8�6����;P��;P�&�^9=���ν03�����&���YS��V7��C>�B�Y�ͻo��}���J�~�stq�;\���@��!��0�� ľ���*7��?Խ�&D��n6����;��;�'��B=���ν53�8���d����X��}:�lG>�M�Y�%�o���}������~��xq�'\�t�@��!�G3��ľ����   �   2-��\� �E���� � �A� &H<��;��{��x]���޽�]6��L���'����2g
�����0��;���?�̃<��!2�"�!��~��A�﷾܆��E�;����oi��֎��{�;H�;< �ƹ]��V������C�������T�y)�_�Q�y�x�r��� ���ף�����c��R���Ɏ��V{�IT���+�B��׿��   �   J=���L\�/�����_�P�(��/b<���<��"<�s�B�Y���ӽB�'�>�l��q������Blݾ}������ڭ�$>�������E������Xs���-�Z�ݽ��i�Pb�� �;�˕<(�N<0�4���`���5[�)��8���='��W�#��%���4��:U����ʿ��ο�i˿e��?j���Μ�3:����X���(�}����   �   �׾n⌾
&�Se��hض���P<LK�<t��<��<p�	���1�����	���=�N�p�v��Q���>��͵��@��3��΢��}qv���C���hV���C��bE���_<���<p~�<��6<���󊤽��&�P���s0׾���3�L�»���v���˺�=�ҿ��t�΁��.����8Կh���Xl��)l����M��Q��   �   Ƌ �[����;N��tԽT���< <�=־6= b'=(L�< wE;�ۼ|�y�NFƽ ��C'�eA�g�Q�FX�$}S�mD�~V+�&��?<н�~��l��� �^��'�<��=&�,=�a=���;�|��Wؽl"P��p���� ��45��q�q����_��hؿ+��������g����8������Fٿ��������Bq��5��   �   ���t�ľ#r��� �4A� ��;�== �a=�Fp=��T=�=Pf�<�1仈��F�j��=����ǽ��߽��nO���̽lթ�qz��^� �3�hVY<�/=��H=�ie=��W=��=��l;�BK���l.u���ƾ��BN�c�����пCq���n��X��|�����d��W��3п�諿���
yM��   �   �W!��پ>������i���;b%=��}=x�=�|�=�qy=.-@=���<H%4<P���¼�C���:�LH���>��?���ؼ(?,����;���<��2=�m=�=zǋ=�&t=zq= �ǹ� v����iQ��<ܾ��"��a��͔����Ὺ�
,�z�!�,�*��-���*�2�!�xA�t�S{ῄ�����ʇ`��   �   T�*�Z羬]������a�� �й^r(=�=�C�=�x�=�Ƙ=Ĩ�=\@P=��=�*�<�p<�B�����C��v&�������;�5�<-= �C=3{=�=�8�=�O�=��=�+=`#R� ��0�"�7Β�l�龇;,��n������Ŀ�=�!
�V��T$*�P�3��7���3�%*����8�	�F{�^�ÿ3�����l��   �   ��-�.�뾱�����"�]���=��E)=��=�=Y[�=���=Q�=�l=5=���<���<�6<@�%; �8�P�:P�;,�<���<�.)=�`=xx�=�}�=�:�=��="��=��=@J������'����ծ�/���r�{r���ȿ,+��l��g��-���6��W:���6��-��:����B�	�ƿ�^��>�p��   �   ��*�2��\�����)`�� �Ϲ�s(=��=�C�=�x�=�Ƙ=Ҩ�=p@P=��=+�<�p<�B�0����C��v&� �����;�5�<-=*�C=&3{=,�=(9�=
P�=N�=�,= R����	�"�^͒�5�龲:,�ۄn�鸜��Ŀ�<�x 
�����#*���3��7��3�V$*�����	�Vz쿓�ÿ������l��   �   JV!���پ�<������i�@�;�d%=V�}=��=�|�=�qy=r-@=���<�%4<����¼�C���:�LH���>��?��ؼP?,����;���<��2= m=��=�ǋ=v(t=�s= �Ź��u�V���O���ܾh�"���a�w̔����+�ῒ~��*��!���*���-�D�*���!�D@�s��y� ������΅`��   �   ���g�ľ�r��� �rA�p��;�@=T�a=�Gp=h�T= =�f�<p0�l��<�j�=����ǽ��߽��uO��̽rթ�"qz��^���3�PWY<T0=^�H=ke=�W=<�=��l;�:K����)u�p�ƾ���#?N�Ca�����gпCn�<�����`��z��������p��1п�櫿+��EvM��   �   B� ������6N��mԽ��pU <� =d�6=�c'=�M�< �E;d�ۼN�y�;Fƽ��C'�jA�l�Q�FX�-}S�uD��V+�,��I<н�~�������^��)�<��=��,=�e=P��;�r��Pؽ$P�;m��� �\15�R
q�Ȼ���\��|dؿ.�����8��he����6�����yCٿ����F��W>q�25��   �   z׾}ތ��&��]��Ķ���P<(T�<�<�<8�	�B�1�����	���=�M�p�w��Q���>��ҵ��$@��3��Ң���qv���C���QV����C��^E���_<8��<p��<0�6<������:�&�B����*׾���r�L�ٸ��s��Ⱥ���ҿQ�忊��|��I��b���Կ�����h��Qi��D�M�:N��   �   �7��E\����D�_�Ȏ(��Kb<���<��"<(ys�@�Y�R�ӽ.�'�1�l��q������Dlݾ�������ݭ�(>�������E������Xs���-�*�ݽ��i��^����;�ԕ<P�N<@�4�
�`�� ���,[�{#������A8'��W����"|�����pP����ʿ��ο�d˿W`���e���ʜ��6����X��(�#����   �   �'��Ϸ �p:��� � �7��@H<0%�;��{�Rw]�9�޽�]6��L���'����2g
������0��;���?�Ӄ<��!2�)�!��~��A�﷾ކ��5�;����dni��ю�@��;8�;< ����>��k����������x��P�es)���Q���x�!���Z���ң���_�����XŎ�O{�RBT�d{+����п��   �   *�6�8Խ(D��I6��9�;0�;��&��6=���ν�/3����� ���WS��W7��C>�F�Y�ѻo�	�}�Ə��U�~�~tq�F\��@��!��0�� ľ
���7�?Խj$D�p_6�@)�;`�;�&��.=���ν|+3���4���iN��]4�U@>�a�Y���o���}�~�����~�$pq�;\�^�@��!�4.���þ���   �   Y�潒bi�����;H�;< �¹DI������x��l���|��CR�v)���Q�~�x�?������?գ�y	���a��	���ǎ�S{��ET�O~+����ӿ��*���� ��?��X� � �:�BH<p@�;��{��l]��z޽�X6��I��}#����6d
�!���0���;���?��<��2���!��{�N<龢귾B�����;��   �    xi��K��O�;Dە<0�N<H�4�Ĺ`�k���0[�&��=����:'��W�R��~������R��4�ʿ*�οxg˿�b��h���̜��8���X�a�(�����:��1I\�����N�_��(��Ib<T��<x�"<XVs�ƠY���ӽ��'�N�l��m�������fݾn���]������:����R���@��r���Qs�և-��ݽ�   �   �3E��	`<��< ��<Ȥ6<���������&����j-׾�����L�:����t���ɺ��ҿ����
�S��Ŧ����%Կ�����j���j����M�/P�}׾����k&�ja���˶�`�P<,W�<<�<�'�<��	���1�尽R�	�"�=���p�%��XL���9������;��7.��]����iv���C�L��M���C��   �   T:�<h�=f�,=pg= ��;�u�hSؽZP��n��@� ��25�Vq����P^��3fؿ�����Z���f����7�����QEٿD�������@q�5��� �����x9N�PqԽ���O <�!=J�6=�h'=�\�<�"F;8�ۼwy�z<ƽs�f='�j�@�
�Q��>X��uS�P�C��O+�B��2н)v�� l���	\��   �   T�H=Doe=��W=@�=��l;=K�2���+u�ƚƾ���j@N�b������п�o�
��z��Z��~�����������x2п�竿&���wM����$�ľFr�M� �"A���;&A=.�a=|Kp=��T=H=ly�<��㻼��f�j��4��һǽt�߽���E��̽@̩��`z�~P�0^3�HY<B8=�   �   ��=bɋ=4*t=�t= �Ź2�u���bP���ܾ	�"���a�͔�2�����`+�©!�n�*�X�-��*���!��@��s��z����������`�4W!��پ~=������i���;`d%=p�}=�=�~�=�vy=L3@=���<XH4< J��¼�7�Ƙ:��>H���>�v3���ؼH,�@��;X��<r�2=:%m=�   �   *:�=�P�=��=x-=@R����B�"��͒�����:,�5�n�&���d�Ŀ�<� 
�����#*��3�Z7�\�3��$*�x���	��z��ÿ����i�l��*��u]��O��0a�� 8й^s(=��=BD�=vy�=�ǘ=6��=�CP=�=�4�<p�<��������C��]&��샻�ҿ; @�<�1=��C=^6{={�=�   �   ��=�ˋ=rZ=�ɻ<���'�ֽ*^�������X����P
��&�Z�N�)��+A���T�4&b�L�f�%b���T��@��)����'���Ͽ�S���:V�2J�<����YZ�M�нLмp��< �`=].�=��=R&�=,�o=
%6=��<�\< Ϲ k;����x��� ���=R��~�`8<PO�<h�,=��f=q�=�   �   �=1Q�=)T=P�<�ؼ�нq�X��	������%T�/����ѽ�w3�����'���=���P�L�]�eb�>�]���P���=���&�|x��񶼿���KnR�����θ�7hU�r+˽H�Ƽ��<p�Z=nʉ=輎=�w�=T\T=6�=��<�c ;��O��ʼ|��P��8����ּ`�p� ��8���<�
=t�J=Hu|=�   �   r�d=�k=��A=�c�<�j��
���",J�����V�	�z�H���Et����ῒ	� ����3��rE��\Q�\�U��Q� �E���3�N�������[����I��bG��z�C����'G��㺽�8��h��<8�H=�r=�l=��C=�W=�=<�&�0� ���N�蚆�c��������ڜ��"����X�����mU���<t3�<�(:=�   �   ��=1=�0!=���<p2��29�� �3�B᝾1d����6�}�|��ƥ�e�Ͽ����� %�d�4��
?���B��M?�~�4��f%�hV�����"�Ͽ�q����{�56�����肜�
11��5���҆�@}�<|(=D9=�*=|��< �b��E�b�{��߹���ｪC�rI�� �)u��v�`���%���f"���T��oػX�<�   �   �N�;��<���<� �< �W��Q���[������ؾ�A ���^�S��_����߿�T����JT �Z7)��t,��)�B� �d������^�v��y����^����/�׾�Ά�����L��H?�4O�<��<�J�<@��;������a���ý�f�\8�y]^��|��w��B.��89��x���*b�9n<����D̽Ƌq������   �   8R��ʻX�#<x�!<�+�րM���𽪞]����s��}=�H>{����	���\�����Xd
�X��*��V9����p���⿝¿@ٟ��)|��=�F���
��$ ]��>ｮI� l��3:<��B<�ks��}��F��X� ��	<�&(z��v��<�����̾k�ھ��߾�۾3\ξ�0��-;������]A�Z��65���   �   �����91��0W����0/�D2�⬲�6�*�dW��C|ؾ����IN�����ǳ���^��w�Կ����k������!��s.�25ֿ�ӽ����j�����O�	��ߙپg+��}����0Cл AG:x�7��p&��s����<�_�A����ľQ��
�
���#�&#'�u($������>���'Ⱦ�s���*e��8��   �   ����}��N�.�8%���pI��`�q�}9���T�+E�� ���""��Q�����-���G諿;㻿#9ƿ��ɿz�ƿ3���>E�����,ׁ�S���#���ߦ��'V�����R�s�܉������k�.a'�s�����"q�Z?����QF�e�+��]E���Y�y�f��~k���g��[�9NG�[�-��V��a�\��lv��   �   ^�p����+m��~���`��v[�.��
&���"�rm���������d�t�D���i��Q���C��x������t'���0���~��~Tl��'G��p �9���
���p�Ҭ�ph��f���`��[�����+���&�Y
m��Ǩ��g�7�D�F�i�4T��`F��'���ʶ��*��n3��%����Xl�e+G��s ���������   �   {⦾�+V����\�s�������k��W'�`�����fq�;����C���+��YE�@�Y�Ŭf��yk�~g�~[�'JG���-��S��\�X��6v����lw��`�.�`����P���q��?��Y!T��H������%"�qQ����������꫿滿
<ƿ�ʿY�ƿ�����G�����ف�G S���#����   �   ��پ>��i+�$������>л�:H:�l7�e&�uk��z��1�_��<��O�ľ1ﾤ�
�Q��1�#�1'��$$�M��F�I���"Ⱦ�o��$e��3����\/1��W�����46�7�����*��Y���ؾ���LN�ҩ��ﵠ�a��+�Կ����n������$��D1��7ֿֽ�������l�O� ���   �   �������"]�B���I��l��>:<�C<@�r�q�F>���� �<��z��q��⺶�с̾O�ھ��߾�۾uVξ�+���6�����DWA�!��7-��xF��Iʻ0�#<0�!<h1���M�`��<�]�i��C���=�IA{����1��_�q����e
��������:�4�s��H�⿊¿�ڟ�d,|��=��   �   7��"�׾?І�7���N���?��R�<<�<\X�<�!�;�}��d�a�p�ý�`�T	8��U^���|�ns���)���4�� ���"b�Xg<�8���:̽|q�li��Е�;���<���<D"�<��W�qT��^�Ҝ��+�ؾHC ���^��������߿V�����U ��8)�v,���)��� ��������`࿁w�������^��   �   P6��������V21�/7�� Ԇ���<(=�H9=�1=���<�7b��7�v�{��չ�����=�@C��� ��n��p���������)���F��ػ��<�=$1=�2!=(��<�6���;���3��❾]f��S�6�j�|��ǥ���ϿS����>%���4� ?���B�O?�� 5��g%�@W�����L�Ͽ�r��R�{��   �   �bG�B{������(G��亽�9����<:�H=:�r=��l=t�C=H_=0(=<��%�� ���N������򚽵����Ҝ�z��RyX�����DU���<|A�<@.:=l�d=:k=,�A=pc�<�n���¿��-J�؜��-�	���H����+u����6
������3��sE��]Q�d�U���Q���E���3���j��]�����?J���   �   �nR�م�ϸ�|hU��+˽0�Ƽ��<��Z=Eˉ=��=gy�=`T=��=t*�<�� ; �O��ʼ����������ּ�p� �8���<B�
=��J=�w|=��=�Q�=p)T=O�<�ؼl�нv�X��
��{��D&T�����Wҽ�4�J��'�r�=�n�P���]��eb���]�.�P� �=��&��x�f�5���*����   �   �9V�J�����zYZ���н�м���<��`=�.�=<��=w&�=\�o=>%6=<��<��\< 	Ϲxj;��򘼰x��| ���=R� ���8< O�<D�,=f=P�=��=�ˋ=Z=�Ȼ<0�ἱ�ֽ�^�����B��BX���q
��=&� Z�^�)��+A���T�<&b�L�f�%b���T���@� �)�n���￲Ͽ�6����   �   �mR�'��θ�*gU��)˽��Ƽ��<��Z=�ˉ=G��=�y�=2`T=��=�*�<�� ;�O��ʼ����������ּЊp� �8ȳ�<Z�
=��J=x|=*��=	R�=j*T=4R�<�
ؼ��н�X��	�����F%T������ѽ�3���L'���=�p�P�ȿ]�~db���]�6�P�*�=�.�&�"x�u�p�������   �   
aG��y����:&G�<ẽ�0�����<
�H=b�r=B�l=�C=�_=)=< �%�̲ ���N������򚽴����Ҝ�y��JyX����DU�(�<�A�<�.:=&�d=bk=�A=@i�<�e��x���+J�욯�Ο	���H��
���s��)��	����(�3��qE��[Q�Z�U��Q�4�E��3����T���ῂ���I���   �   �6�h���_����.1��2���ǆ����<��(=�J9=�2=���<@1b�x7�L�{��չ���ｼ=�=C��� ��n��p������������F��ػ��<�=�1=T5!=D��<*���6��|�3�����b����6���|��ť�5�Ͽ3���2�%�<�4��	?�V�B�|L?�L�4��e%�xU�����źϿ�p���{��   �   /����׾,͆����H��`?�d\�<L�<\�<�*�;�|�� �a�L�ý�`�L	8��U^���|�ns���)���4�����"b�Wg<�2���:̽�{q�8h��О�;X �<���<�+�<�mW��N���Y�������ؾ+@ ���^�$�������߿�S�����R ��5)�s,���)��� �*�����]�tt��#����^��   �   ���&��V]�9��vI��L�XS:< !C<�r��o��=���� ��<��z��q��ߺ��ρ̾O�ھ��߾�۾xVξ�+���6�����:WA����,��@E� :ʻ��#<(�!<��RyM���k�]������m=��;{���"��vZ�<����b
��������7�b��m����⿎¿{ן��&|���=��   �   S�پt쎾,c+��w������ϻ��I:�_7�c&��j��N���_��<��H�ľ*ﾢ�
�Q��1�#�2'��$$�P��H�L���"Ⱦ�o���#e�u3�����t-1�`
W����@��*�ۧ����*�U��yؾ���GN�N���ȱ��\\���Կ����h���������+鿇2ֿPѽ��򡿜���ĪO�����   �   0ܦ��"V�,����xs�xv�������k��T'�w ��K��@q��:��w��C���+��YE�?�Y�Ƭf��yk�
~g��[�+JG���-��S��\�X��v�����v��F�.�`�H���8��B�q��2��"T� B����_ "���P�����𘗿�嫿�໿I6ƿ��ɿ��ƿm����B��a��� Ձ��S��#�l��   �   �p�J���a��rz�h�_�pZ[�����$��)"�>m�쉯�����d�r�D���i��Q���C��z������v'���0���~���Tl��'G��p �>������p�r��g����8�_�0U[�������v���l�M������a���D���i�O��KA��֡��b����$��V.��m|��/Pl�$G�hm �$������   �   Ɔ��o���.� �~�`���<��r�q�V8��HT�E�����""��Q�����-���I諿<㻿%9ƿ��ɿ~�ƿ8���DE�����1ׁ�S���#���zߦ��'V�q���h�s�P}��`��(�k��L'�/������q��6��b���?��+�~UE�؊Y� �f�uk�Vyg��	[��EG���-��P�-W羷S��jv��   �   i����!1���V���� ��-�F�����*�GW��7|ؾ����IN�����ǳ���^��y�Կ����k������!��y.�85ֿ�ӽ�
���o�����O���ۙپ��f+�6|�����л <J:@F7��X&�xc��D����_�{8��A�ľD�L�
����V}#�@'�� $������"��Ⱦ.k���e��-��   �   �8�p�ɻX�#<�!<���|M����Q�]����p��=�I>{����	���\�����Zd
�Z��.��Z9����p���⿦¿Eٟ��)|��=�G���
���]�t=ｔ{I��Q�8Z:<�3C<�;r�Nd��5���� ���;�z�Vm������|̾G�ھ��߾�۾�Pξ0&���1��S��fPA����T$���   �   ��;�< ��<�/�<0pW�]P��h[�������ؾ�A ���^�U��`����߿�T����LT �`7)��t,��)�H� �h�����_�v�������^����)�׾�Ά�0��mK��h	?�^�<��<�g�<`p�;�d����a���ý�Z��8��M^��|��n��%%��D0��i���b�B`<����0̽,kq�0N���   �   ޖ=�1=N8!=���<H+��8��І3�.᝾)d����6���|��ƥ�g�Ͽ����� %�f�4��
?���B��M?���4��f%�lV�����*�Ͽ�q����{�86�����؂���01��4���ˆ�至<��(=�N9=�8=ع�<��a��)��{�;̹�	���7�=�p{ ��h��j������������n8���׻$,�<�   �   ��d=� k=�A=�j�<Pf��R����+J�����U�	�{�H���Et����῔	�"����3��rE��\Q�`�U��Q�$�E���3�T�������^����I��#bG��z�9����'G�㺽D4��T��<6�H=�r=&�l=D�C=~f=K=<`�%�� ���N�F���뚽엢�0˜���~kX� ��U���<Q�<�4:=�   �   O��=�R�=�+T=�S�<t
ؼԜн[�X��	������%T�/����ѽ�x3�����'���=���P�L�]�eb�@�]���P���=���&�~x��󶼿���NnR�����θ�"hU�'+˽0�Ƽ�<��Z=̉=(��=�z�=lcT=��=D4�<�!;�{O��qʼ΅�X��r��t�ּ pp� 8�8H��<��
=��J={|=�   �   z��=�r=�-=` <UL���{���y�S1��~��k���Ὺr� *��H��^f����0��J4�����%���f��H�W)������߿SX��X%}���/�������P ��G�D<.G0=�v=��=��q=|B=Z�=�i< =G�����]��F��:
+�<F!�����b��`9����M<��<<n<=�Km=�   �   :q=ؐf=H�&=�B�;~�F�a�
�삆�����-�~Uz��z���WݿN"
�\'���D�
�a�:�z����.�������z�j�a��xD�F�&��	��3ܿV����x�m�,����9�����2�A�J<��)=��i=�Hu=(�Y=N?#=���<�V;l1�� ����<�F�`�^�m��c�*aA��������*�:��<*-=��T=�   �   �9=.�@=�=�@�;r�6�,� ���{���Ծ�/$��0m��졿C�ҿ�s�z���{:��U���k�f�{�%�����{�X2l�~6U�Zc:��p��ѿQ2����k�:6#��Ӿ��y�z���`�1�p��;@�=��D=�y>=v�=���<�
���%��tV_��㛽S��g�սj_޽Jw׽�������&h�Ҁ���@�u<��	=�   �    ��<��<���<��;����� �a�:���T0���X�4�������.����*��JB�nV�0�c�6�h���c��V�@�B�D,+�"�v�i��w!���W�݌���`����H�����;���<�T=�b�< �;�̽��9b�_&��Z���ӟ�T5��E��J��F���6����� �k弽m���м`v;�   �   P� �;p�T< �N:����P����@�����6�1u>�lc���>��!�׿2A�N����+�`o<���G��K�h�G�.=��,���О��Pؿ\��hY���:>�Z��������?�[���J� ��:�g<8W<�/��h,��㨽����E6���g��ى��x��e�>#������ݱ���z���3k�4	:�F������6��   �   ��t��ͼ`�ֻ�Hڻ2輽���*��C����پ�� �l�_�����"��J�t?����!�П*�:�-�r
+�XP"�|�����5�亿�.���N`�-!�(�پ0��*������`g�P��������-��V�j�P׽�(���l�EO��e����.ݾ�_��"a�3\�������Y߾H�������6q�$,��ݽ�   �   ����2����|ϗ��Gּ��n��>�g�W�����+�c7�|�s�c�������ۿ����*�^e���N��.���k���Dݿ�E��ᦛ�& u���7�.������LXX�n��.�m��Ѽ�
� ��ꅽ���O
@�����7*�����jt��u%���6��BB�~_F�2�B��8���&������0����[��.�C��   �   DJ�`j��jȈ��������[3�ې��B��>ヾ��Ⱦ�&��@���v��-��������ȿ�8ۿ翷k�ٽ�K[ܿFDʿ����l��uy�=[B��@�Xʾۄ�X� ����2�3�?߼�:��������j�F�M��xоX���+�[%L�v�i�df��`ꇿã��bO����nek�� N���,�|�
���Ҿq;���   �   �/��N�=��޽n�n��V	�bR��k�(۽�U;�D����Ծ
���<���h�+͉�����aw��N��܄�������b��ʝ�I��s1k�w>���A?׾�,���=�4
޽��n�FU	�BU�r�k�s.۽�Z;�������Ծ����<���h��ω�v���Tz��a�����������e���̝�����5k��z>�N�xC׾�   �   �[ʾj݄�t� �������3��;߼5�W���q���F�h
��mо5��8+�!L���i��c���燿����L��~���`k��N�4�,���
�F�Ҿ�7��J�c���È�2��l���_3�R�������僾��Ⱦr)�c�@���v�40��Y�����ȿ�;ۿn�o�)��o^ܿ(Gʿ?��o��3y�B^B��B��   �   ���E����[X�T�򽆳m�ЬѼ<돼�� �Z䅽a��@���%������p��q%���6�K>B��ZF���B��8���&�J����R����W��L�C�}z��-����Dɗ��Iּ��n��C�p�W�����-�$7���s�~���&����ۿ������$g�L�������n���Gݿ�G��̨��E#u�6�7��   �   �!���پ�1��(�������g�0����Ǫ�D����j�7F׽�(�҄l��J��ۉ���(ݾY���]��X�&��Y����S߾��������q��+�̬ݽ(�t��	ͼ0cֻ�9ڻX5輐������E����پ�� �/�_�P��� $�����@��	�ڞ!���*��-�D+�R"����\���7��庿30���P`��   �   �<>�}�������?�4�����@�:�g<0v<��/�Z,�*ڨ�����>6�eyg��ԉ��s��*����ŕ��𬜾nv���+k�a:��~����6�6���O��J�;��T<��N:���S��6�@����98�-w>��d��5@���׿XB����4�+�q<���G���K�:�G��=���,���ҟ�tRؿm]��xZ���   �   X�W�ȍ��񾾈`�0����@��;P��<Z=|r�<`q�;0����)b����
������z5��
E���J��F�.�6�h��� ��ۼ�Tm�`�м@;h˲<|��<���<��;���h�M�a������1�J�X�O���n����0��(�*�ZLB�V��c���h�:�c�j�V���B�L-+��"���j��Q"���   �   ��k��6#��Ӿ��y�z�����1���;��=*�D=>=(�=�҉<෿����JH_�ܛ����w�ս_V޽in׽P���L���l�g��t� ��(v<��	=��9=�@==�>�;��6�D� ���{�
�Ծ�0$�?2m���L�ҿXt�<��r|:��U�<�k�ĳ{�ձ���{�z3l�p7U�d:�������ѿ�2���   �   1�x���,��:������A��L<�)=��i=,Ku=��Y=�C#=��< W;�#��n~�v�<���`���m�fc�2YA����Ј�� ��:X"�<�0=p�T="<q=
�f=��&=P>�;�F��
�������ᾣ�-�JVz�{��kXݿ�"
��'�2�D���a���z�u��/��	��P�z��a�yD���&�F�	�4ܿ����   �   %}�r�/�k�侭�� ��G�xF<�G0=�v=:��=�q=�B=��=�i<@9G�X����\��*��2
+�@F!����,c���:�� �M<���<�m<=VKm=T��=��r=�-=� <�UL���J{��z澃1�B�~��k���῾r� *�&�H��^f����5��J4��������f��H��V)������߿1X���   �   �x�֖,���V9�����f�A��S<6�)=l�i=�Ku=��Y=�C#=8�<@W;�#��^~�b�<���`���m�hc�.YA�����������:�"�< 1=��T=�<q=ƒf=ʋ&=L�;h�F��
����������-�'Uz�Wz��{Wݿ"
�'�H�D���a���z����\.��P���z�Φa�4xD�ډ&���	�)3ܿ�~���   �   f�k�F5#��Ӿ��y�������1����;��=v�D=�>=��=\Ӊ<ൿ����*H_��ۛ����p�սYV޽an׽H���A���T�g��t�x��@v<d�	=t�9=f�@=(=�Y�;r�6�F� ���{�͕Ծ/$�0m�졿��ҿ>s�����z:��U���k��{�x���b�{�1l�p5U�xb:�R~����ѿ�1���   �   g�W�����t�_�˓����ҿ;0��<�[=�t�<w�;@���L)b�}�����w��p5�~
E���J��F�*�6�`��� ��ۼ�m���м�;�Ͳ< ��<���<��;����� �a�����b/�F�X�W�������x-�6���*��IB��V���c�z�h���c�^�V��B�++�"!���Sh��h ���   �   9>����~�����?�Ȃ�������:��g<�~<��/�HY,��٨�����>6�Wyg��ԉ��s��&��������jv���+k�X:��~����~�6���O��[�;h�T< P:v��XM��@�@�����5��s>�Zb��?=��r�׿.@���6�+��m<��G�0�K���G�|=���,��������Nؿ�Z��)X���   �   !��پ�-���������U�0n���������T�j��E׽`(���l�wJ��щ���(ݾY���]��X�$��T����S߾��������q��+�m�ݽЇt�ͼPEֻ`
ڻ�"�y���p��A���پ�� �
�_����. ���&>�|�p�!� �*�\�-��+��N"�������a3�⺿-���K`��   �   �������SX����Z�m�H�Ѽ8ߏ�Բ �8ㅽ����@���%������p��q%���6�I>B��ZF���B��8���&�I����L����W�� �C��y���+����`����6ּP�n��8򽇹W���*��7�Z�s�u���d���t�ۿ�������c���������sh��BݿCC��̤���u��7��   �   /Tʾ؄�� �t��� y3��)߼V/�����a��W�F�S
��`о/��2+�!L���i��c���燿����L��|���`k��N�3�,���
�?�Ҿ�7���J�b���������0R3����z������\�Ⱦ�$��@�
�v��+�������ȿ�5ۿ��Xh뿂��XܿIAʿ����vj��p�x��WB��=��   �   [)��Ǔ=�J޽�n�RJ	�BJ�ʚk�u&۽�U;�&����Ծ���<���h�)͉�����`w��M��܄�������b��ʝ�J��u1k�w>���9?׾�,����=��޽|�n�0M	��H�ޔk�� ۽=Q;������ԾI����<���h��ʉ����~t��C����m����_��Cǝ�����-k�gs>����:׾�   �   �J��Y��ͼ�����D�⼺T3��������ヾ��Ⱦ�&��@���v��-��������ȿ�8ۿ翷k�ڽ�M[ܿHDʿ����l��yy�@[B��@�Xʾ�ڄ��� �٠��(}3�`)߼�*����'���F�����о=���+��L���i�@a���䇿H����I������[k�MN�o�,�^�
�0�Ҿ�3���   �   {p��d%����������5ּ��n��<��W�����+�a7�z�s�b�������ۿ����(�^e���N��0���k���Dݿ�E��㦛�, u���7�+�������WX����Z�m��Ѽُ��� �_݅�-����?��> �����im��m%�i�6��9B�UVF�.�B�>�7���&�������-񽾰S����C��   �   &yt�p�̼Pֻ��ٻX#�b���u
�\C����پ�� �n�_�����"��J�t?����!�ҟ*�<�-�t
+�\P"�~�����5�亿�.���N`�.!��پ�/��x��Q����X�p_���~������j��<׽k(�7}l��E��w���y"ݾsR��Z� U��������RM߾K�M����q���+���ݽ�   �   @�O�Й�;��T<��P: ��7O�� �@�����6�0u>�mc���>��#�׿2A�L����+�bo<�G��K�l�G�4=�"�,���Ԟ��Pؿ\��lY���:>�V��s���j�?����������:��g<x�<�c/��K,�Ѩ�/���76�qqg�yЉ��n���禾����������q��l#k�F�9��x�6�����6��   �   tݲ<@��<4��<0#�;z��|佨�a�&���Q0���X�7�������.����*��JB�pV�4�c�8�h���c��V�D�B�H,+�"�|�i��{!���W�ی��𾾴 `�i��R���ӿ;���<�`=���<�Á;\����b�&�����N���5�cE�j�J�a�E�H�6��I� �Ҽ���l�Īм@�;�   �   ��9=�@=d=�`�;ܑ6��� ���{���Ծ�/$��0m��졿E�ҿ�s�z���{:��U���k�j�{�'�����{�Z2l��6U�^c:��t��ѿS2����k�:6#��Ӿq�y�������1����;�=J�D=>�>=��=�<0h��$����:_�Kԛ�h�����սYM޽{e׽����T����g�jh��a��/v<"�	=�   �   8?q=��f=�&= R�;:�F�4�
�߂������-�~Uz��z���WݿN"
�^'���D�
�a�<�z����.�������z�l�a��xD�H�&��	��3ܿW����x�m�,����9�������A��Q<��)=��i=�Mu=��Y=lG#=l�<�hW;��� w���<�V�`�&�m��c��PA����z�� ��:�,�<V5=*�T=�   �   ��d=��R=:�= ���l@��j�,��Ӡ�̡���I��Y����ÿt%���H�0�@���e�$���3�����������?������Z��^oe��C@�,������¿/����I�x
�#����+��捽�r�� �=Z�Q=B�d=ޏM=�L=�4�< ��:H\��.1�P�C�^-g���s�"�h��F�ҩ��ԗ� ��9а�<��=��L=�   �   ��P=�E=T��<���������(��~�����EF�Q֍�j<��������hs=�dwa����^�����������[��옂�a���<�@������m���;���mE����ۜ�F)(�	��������j�<V~D=	Q=P�2=D��<�%<�)3�h���rM��Ƅ��4���0�����oA��zJQ�F��(�B��8<|2�<��1=�   �   b�=��=p7�<`Qѻ���E���哾51���;����󼶿S����V�3�X�T�֏u�����ܒ�hf�����M(��j�u���T��^3�Ш�*G쿊'�����8�:��U��e��P[�����0�һ���<��=��=�< &o;����:9F������6ʽ�����)p	��t�x���̽�D��$�K��Է��;8;�¾<�   �   ��'<���<��<��
��dj��A��!���޾�*�+)v�uڧ�&/ڿ�A�V�$��B��_^���v�}у�n��j����Iw���^�TRB���$�f1���ٿr�����u��[*� �ݾ;҄����F�i�� 
� ـ<�%�<��1<�.�f�&�f2�����(�t>=�gX�>j�gWp�*�j���Y�S�>�l�-��=���&,��n>��   �    }�� �:�S�0O�d�q�e�&���<~�(�X��Ӕ��H¿"󿜯�n�+�NC��>W���d���i�jDe���W���C��D,�~�Cg�k¿�֔���X�/d�����[e��'򽬳N�XCQ���i:�آ���ۼ��|�!�ڽcg"���Z�4׈�����1��6���хƾ9r¾��ῢ�W1���O]�#�$��޽�����   �   ���*��髼Dʬ��	9��5ȽhV=�����A���7��M~�h��C�ѿ�b�����,'�7�"�A��E��(B�2�7���'�(���h��gҿ�z��!�~�z48������̠�D=��IȽ��8��@��L覼��%�Nᠽ�;�'�J�Pދ��R����۾&K��������.��1��^��} ���ݾ++�������M�2h	��   �   v�����|M�����.�m���H��S�Qʾ-����P��U��Hݮ�R�ӿv�����JD�>� ��#��� ���^H�r���cտ����>�Q���ϸʾ���f��6����C.��2
�t�I��Բ�#����e��!���TپM
	��$�QB=���P�0U]�c�a�C�]�N�Q��i>���%�^C
���۾򤾱�h��   �   �o���������Y�~�5�Jg�U�߽��@�Pǚ�	`�26$�z�[��-��	���kȿ�Z�S���\�0y��]�����^��j�ɿ@��5��.]�&%�6��c���v�A��������4���W��౽T�0$m��c�����;L��C���h�鳄�������윿�G��1:���x���Bj��,E���� �&���   �   m���r�a�B�	�hǠ���P�V�O�]|��:��d�_�Cd��E%����&�.W�dc��t%��;��
���I+̿�ϿО̿�[¿����-���U���X�d5(���������a�0�	�Ġ�f�P���O�����҉���_�h��p*��?�&�.2W��e��9(��J��R����.̿��Ͽ5�̿(_¿���J0��X����X�y8(��
���   �   �������A�
��F���4��~W��ڱ����m�__����H�ՙC��h�9���7�����霿�D��Z7��[v���=j��(E�=�������9�o���������Y�,�5��k�L�߽ �@�hʚ�bd�9$�*�[��/������nȿ:^�����>�{�p_�,������H�ɿ���K��s1]��(%��   �   ����ʾc���������B.��-
���I��Ͳ������e�^��Oپ�	��$��==�&�P�"P]�F�a�>�]���Q�)e>���%�@
�8~۾���h���������wM�(�|�.�7���!�)X��ʾ�����P��W���߮��ӿ-y��j��:F�L� �$�#��� ����J�i����տB���L�����Q��   �   w68�]����Π���=�LȽ��8� :���٦�8�%�/٠�v6��J��ً�@M��G�۾$D��������$��-�[�Jz ���ݾ &��Q���S�M�c	�����*�ޫ� Ƭ��9��8ȽZY=����pD��k�7��P~�T����ѿne��f���-'�"7�V�A�0�E��*B�.�7���'����Zk��w�ҿv|����~��   �   ��X�we�����^e��)�|�N�h:Q� 1k:����$�ۼH�|���ڽ�`"��Z��҈�����S,��S����ƾ`l¾~��Ӻ���,���G]���$��޽㈁��f伐��� �:`�S��O�Wg�Q�e�c�����]�X�cՔ��J¿K�����+��OC�AW��d���i��Fe���W���C�hF,��	�i�l¿�ה��   �   3�u��\*���ݾӄ����0�i��
����<�1�<X�1<�.���&�D)�������^7=�b_X�*�i�4Op�$�j��Y�^�>�D�����x���,�@C>�0�'<乧<H�<�
�|gj�SC�"#���޾v�*�+v��ۧ��0ڿ�B�|�$�&B��a^���v��҃����u����Kw�Z�^��SB���$�*2���ٿe����   �   C����:��V���e���[�������һ���<��=j�=�'�< �o;�����+F����*.ʽ]����k	��o��򽃫̽=��yK�Ⱦ����8;$о<X�=�=h:�<�Sѻ��~���擾�2���;�҇��ྲྀ�x�����:�3�v�T�6�u�h���ݒ�Cg������)����u���T�<_3�X���G�-(���   �   �;���mE���2ۜ�j)(�����`����m�<��D=�Q=�2=���<�&%<3�ē�vjM�&��/���+�������<��VBQ�����B�M<�:�<,�1=�P=E=0��<`��������(����q�AFF��֍��<������h���s=�xa�岂�{^��G����( ���[��8����a��<�~�U����m���   �   ���|I�O
��"��0�+�Q捽 m����=̶Q=��d=.�M=�L=h5�< ��:�[���0�*�C�B-g���s� �h�$�F� ��`՗� ��9T��<V�=:�L=h�d=��R=��=�����@��,�Ԡ������I��Y��ۀÿ�%���H�J�@���e�0���<�����������:���螕��Z��Doe��C@������d�¿�   �   Q;���lE�?��Rڜ�@((���������Hp�<B�D=fQ=\�2=��<0'%<�3����^jM���/���+�������<��FBQ���� �B��M<;�<|�1=��P=�E=���< ���>��x�(��~����QEF�!֍�&<���������s=��va�1����]��^�����@��+[������ta�H�<���R���m���   �   ��&�:�\T��d���Y������һ0��<b�=`�=()�<`�o; ���N+F����.ʽO����k	��o���u�̽=���xK�d�����8;@Ѿ<@�=z�=?�<�6ѻ3��F��7哾=0��;�;�����M���|�쿄����3�f�T���u��
��ܒ��e��?���'���u���T��]3�"��F쿥&���   �   �u�ZZ*��ݾ�Є����H�i��
���<�5�<��1<إ.��&�)�������O7=�W_X��i�&Op��j��Y�R�>�8�����P����,�H@>�((<콧<P�<��
��_j�B@�� ��t޾��*��'v��٧��-ڿ�@�Z�$�|B�B^^���v�sЃ�W��Y����Gw�"�^��PB���$�~0�K�ٿA����   �   ��X��b������Xe��"��N�`"Q� %l:����4�ۼ\�|�N�ڽ�`"��Z��҈�탡�L,��L����ƾZl¾y��ͺ���,���G]���$���޽z����c伀�����:P�S�FO�`�Ďe�E����|�X�X��Ҕ�CG¿A	�r���+�`LC��<W���d�H�i�"Be���W���C�tC,�8�'e�Fi¿+Ք��   �   '28����4ʠ��{=�6DȽΔ8�-���Ѧ���%�cؠ�76���J��ً�3M��=�۾D�������� ��-�[�Fz ���ݾ�%��F���/�M��b	�J���d*��ի�����9��0Ƚ_S=�����>���7�9K~����1�ѿ0`��P��X*'�7���A���E�r&B�&�7��'����(f��}ҿ�x���~��   �   {�Z�ʾ������6󠽦8.�'
���I�D̲����K�e�L��Oپ�	���$��==�!�P�P]�A�a�9�]���Q�&e>���%�	@
�.~۾���h�P��@���fsM���2�.�J����OO�Pʾ����P�T��$ۮ���ӿs����hB�:� ���#��� ����F�M����տ̴���슿0�Q��   �   ˦� �����A���ཿ��:�4��xW��ر�3�dm�F_�����H�ϙC�ݙh�7���4�����霿�D��X7��Xv���=j��(E�9��������o�������n�Y�`�5��\��߽Ɲ@�lĚ�\辐3$��[��+��� ���hȿ�W�������Fw��[������e�ɿ����	��f*]� #%��   �   �����a�ƫ	�-���F�P�h�O��y��^����_�"d��2%����&�.W�bc��r%��8�����G+̿�ϿϞ̿�[¿����-���U���X�c5(�
��ػ��,�a�X�	�X�����P���O�Av��P���_��`��{ ����&�@*W�a���"��D��ӊ���'̿��Ͽc�̿�X¿����*��SS���X�2(�� ���   �   o�o�o��������Y�|�5��_���߽D�@�ǚ��_�-6$�v�[��-�����kȿ�Z�P���Z�.y��]�����]��i�ɿA��6��.]�&%� ��5���ĵA��������4��sW��ӱ�*��m�@[�����bE�ЕC�8�h�����_����뙿�朿�A��q4���s��9j�W$E���������   �   ��癵��iM������.�+���H�S�.ʾ&����P��U��Hݮ�Q�ӿv�����JD�>� ��#��� ���`H�s���cտ!����?�Q�����ʾ<��n������9.��#
���I��Ų�ƻ���e�����Iپ�	�%�$�y9=�b�P�K]�$�a�+�]���Q��`>���%��<
�lx۾餾�{h��   �   �����)�tǫ�D����9�3Ƚ�U=������@���7��M~�j��B�ѿ�b�����,'�7�"�A��E��(B�2�7���'�(���h��hҿ�z��&�~�y48�x����̠��~=�\GȽ��8�)�� Ʀ���%��Р� 1�2�J��Ջ�H��7�۾H=����������)�3W��v �X�ݾ� ��Ѐ���M�M]	��   �   K� [�� �:H�S�O�.b��e� ���6~�'�X��Ӕ��H¿$󿜯�l�+�NC��>W���d���i�lDe���W���C��D,���Gg�k¿�֔���X�)d�����s[e��%򽔭N��Q� +m:PF��,�ۼ0�|�Y�ڽxZ"�q�Z�$Έ��~���&��x����yƾxf¾�������;(���?]�&�$��޽6����   �   $(<<ʧ<�<0�
�n`j�$A��!���޾�*�,)v�wڧ�)/ڿ�A�V�$��B��_^���v�}у�n��k����Iw���^�VRB���$�h1���ٿv���Ũu��[*��ݾ҄�S����i�P
��<�?�<h�1<@{.�<�&�l ��E�齪�f0=��WX� �i��Fp��j�\�Y�6�>�������*���,��>��   �   ��=x�=�C�<�.ѻq������哾*1���;��������T����V�3�X�T�؏u�����ܒ�hf�����N(��n�u���T��^3�Ҩ�-G쿍'�����8�:��U��e���Z�D����һ���<j�=0�=�6�<�Mp;����JF�x���%ʽ�����f	��j�z�򽕢̽5��kK�<��� f9;4�<�   �   t�P=�E=��<����(����(��~�����EF�S֍�k<��������js=�dwa����^�����	������[��혂�a���<�B������m���;���mE�����ڜ�)(�\��������p�<��D=�Q=j3= ��<�;%< �2����DbM�����N+��'��7���e8���9Q�P��H�B�xd<�D�<6�1=�   �   ��L=�9=P��<����N���DD�m䲾���]��N��,lԿ$t	��n,�"�S���~�����1���)F��/����E��ͬ��Xޔ��;~�^/S�.�+��	�D�ӿ����\���E���E�.���������<��3=�fH=b�/=��<�z6<(�����Ξ@��gz�����X;��X���z{��RA���0W���;<�t�<jg3=�   �   ��7=��*=p�<%���Ω�	$@��H���D�Y�S�����пB2��{)�<�O��gy���������0��〴�L6���������*y�SO�j)�X��usп�Q��8�X��1�u����@�� ��$9����<��%=�f3=�d=H��< �#9���_5�Z ��pܢ�MV�� ��훷� Q���}��<6���� A�9���<��=�   �   ���<��<`�<P����	�� M4�0㤾Y2�N|M�b���ұƿ�� �	!���D�ȶj��|��@&�����z��������>��ш���j�p_D��� ��w �dƿh����NM��/����5�`���ߑ�,��<�U�<x�<��p<M���	�F��M���q�����2�����j�M�t�､_��uр���	�0ڻ�{y<�   �   �D�:� H< ��;X�������V"��┾@Y���_;�Kn��ñ����� ���3��U���u�z@��	�������4���r���Mv��XU���3���쿋���e^��	Z;����/���'#������C��P��;�J<<��M:`��b�_��T��H	��2���V�St�vl��輆�������t��W���2�Z�	�H���`������   �   �q"��À�(�`2��KB��@��� ����վ�h$�nm��=��9Dӿ������;���V��m�Ƈ}�������}��5n��)W��'<����7�-nӿ�T��ŏm�O�$�P-־�]��be�ׄ� Ǽ�W�\���v�"��x�����j:��Aw�Ji����kNɾ( ׾��۾"I׾��ɾĴ�R���x�%};�ּ��%���   �   �MĽ$c^����P8��~n�>�뽌mV�~в�f�
�}�I��ꊿ����#�v�	��!�֣6�h�H���T�r?Y� #U��+I�87�:�!��%
�'��)P���&���J���
�8A��Q7W�>��P�p�F�������]��Výh�"jf�eޜ���ȾL�����_-�2�%�nn)�f1&�ߑ�{|�������ɾ�ĝ���g�����   �   ��-��P׽�+��.�=�Qc�����E�*�R����߾��$�O�d����tx������������%��>/�d�2���/�Jl&��s����c�_������^ne�V%���ྣ���ک+�o���x�d��Q>�WՁ��9ֽ��,�V����!��D�J��05���O���d�jLr�lw�S�r��]e���P���5�i��P��-���s���   �   U��ܗ-���ս�ֈ���j�SJ�����EZ�B���t| �x�4��p�����a���"ڿg4���9��q������Ș�����ۿc%��E����q�DI5��� ��Z�� @[�P��	���*k�}����Խ��,�P���HE¾�6��C-���V��~�o��u�)ާ������[���������,�W�#.�����Qþ�   �   �ʿ�]�}�0m�J������^ǃ���\���r|��ܾ�����7�S�k�۾��]_��������ҿ�޿���a޿H:ӿϠ������c���l�`�8�N���ƿ�*�}��i��������Ƀ����;���x|�&ι��4�7���k�w���Yb��8���9�ҿ޿��oe޿�=ӿ���c��f��1�l���8����   �   �� ��]���C[�<R�t���(k��y����Խ�,�͔���@¾�3�@-�%�V�ѽ~����X��ڧ���������X��⎑������W�p.�����Mþ�Q��t�-��ս?Ԉ�,�j��L�����^JZ������~ ���4��p�����d���%ڿ8���;�t���������y���ۿ(��������q�L5��   �   �%���ྮ���@�+������d�LL>�DЁ��1ֽL�,��������	���F��,5���O���d��Fr��w��r��Xe��P���5����J�8)���o��ӏ-��I׽6'��r�=�Rc�����I�*����}�߾A�$���d�����z�����ԓ������%�@A/���2� �/�bn&��u�V�Df翮��ׂ��Pqe��   �   J�G�
�CC���9W���콺�p����F��J�]�Nýv��nbf��ٜ�üȾ���0��@)���%�j)�-&�Ѝ��x������ɾ鿝���g�"���EĽFX^�0��6���n���뽼pV�Ӳ�?�
��I�]슿�����%���	�N!��6���H�|�T�BY��%U�.I��97�ޑ!�"'
�c���Q��l(���   �   ��m���$�//־�^���f��ׄ�L�ƼA� q��H�"��o��� ��c:�(9w�Nd��v��SHɾ��־x�۾�B׾��ɾ����y����x�Wv;�r������e"�l�����`0���C����s��.�վ�j$�vpm�B?��"Fӿ��`��P�;�ڤV�T�m�r�}����N�}��7n��+W�2)<�J���8��oӿV���   �   ,_��([;������0���(#�����@����;pd<<��O:���p�_��J��d	��2�@�V���s�h��w���7�����t���W��2���	��>���x`�T����P�:H<��;���p��mX"�P䔾e[��a;�So������
��!��3��!U���u��A��H��Π���5���s���Ov��YU���3���n�쿒����   �   쎒��OM�0�f���5�����ݑ�h��<`^�<|�<`�p<@��p�	��>����������J-�9��\e�H�)z�bW��cʀ���	�0�ٻ�y<<��<���<|�<���F��rN4�K䤾.3�{}M�*���Ҳƿ_� ��	!� �D��j�R}��*'������u���v���g?������.�j�:`D��� �x ��dƿ�   �   �Q����X�2�Mu����@�� ��t7����<B�%=�i3=�h=X��< �)9D���V5������ע�!Q���y��֖��WL���y��t6���� �9tʫ<�=$�7=:�*=q�<|&���ϩ��$@��I��SE��Y�̛��+�п�2�6|)�صO�`hy������c1��k����6��,������y�~SO��)�����sп�   �   ����;\������IE��������$��<4�3=gH=��/=���<�{6<���(��@��gz�����Q;��a����{�SA�x��0X��;<t�<g3=r�L=�9=,��<(����N��2ED��䲾��]�O��VlԿ:t	�o,�>�S�ơ~����<���/F��/����E��ì��Jޔ��;~�B/S��+��	��ӿ�   �   !Q����X�\1�Yt��o�@����H3��H�<�%=,j3=�h=Ȝ�< �)9���V5�����uע�Q���y��̖��OL���y��b6�d�� �9�ʫ<H�=��7=�*=�s�<L"��OΩ��#@��H���D��Y����G�п2�v{)�ڴO�gy�;���)��[0��^����5��;��K���jy��RO��)�����rп�   �   �����MM��.����N5�����Ց�|Ņ<�a�<|�<�p<����	��>�����֏����A-�0��Qe��G�z�OW��Hʀ���	��ٻ��y<8��<���<L�<8���2��L4�t⤾�1��{M�ݾ��"�ƿL� �f!�.�D���j��{��k%��������������=�����֧j�t^D�&� �w �#cƿ�   �   b]���X;��|��;.��B%#������5����;@m<< /P:�����_�{J��K	��2�.�V���s�
h��o���0�����t�~�W���2���	�>��`x`�Ĩ��@{�:�H<0��;8z��0��U"��ᔾ�W��e^;��m�������� ���3��U���u�b?�����B���C3��yq���Kv��VU���3�����A����   �   i�m���$��*־�[���b��҄�P�Ƽ�0��k����"�qo���� �nc:�9w�Bd��l��JHɾ��־r�۾�B׾��ɾ����q����x�:v;�H��6��d"�l��� ���#���>����r�����վfg$�!lm�p<���Bӿ������;���V���m�(�}�[����}�23n��'W��%<�����6�KlӿJS���   �   SJ���
�~>��V3W��콸�p����Γ���]�@Mý0��@bf��ٜ���Ⱦx��*��:)���%�j)�-&�ˍ��x������ɾۿ��p�g�����DĽ�U^�ƽ�/��un�)��JjV�:β�Д
�R�I�H銿��� ��	��!��6�&�H�r�T��<Y�� U�v)I��57�v�!�L$
����N��[%���   �   �%�΍�瑏�ͥ+�������d�4E>�΁�l0ֽ�,�_����������F��,5���O���d��Fr��w��r��Xe��P���5����J�()���o��n�-��H׽ %��l�=��Fc������*������߾��$�Z�d����&v�����~����v�%��</��2�r�/�$j&��q� ��`�����~��ke��   �   "� �W���:[�"L�V��Jk�-v��~�Խh�,�����l@¾�3�@-��V�˽~����U��ڧ���������X��ߎ�������W�k.����oMþ�Q��ڒ-��ս�Ј���j��D�����WAZ�!���Nz ���4�j�p�?��7_��lڿ�0���7��o�r����Ж�[����ڿ�"��ٶ�� �q�F5��   �   p¿���}�e�>���
�������o��:r|��ܾ�����7�M�k�ؾ��[_��������ҿ�޿���a޿E:ӿ͠������c��
�l�]�8�G���ƿ���}��h������������u�� ��	m|�پ�@
�B�7�,�k�a����\������4�ҿ#޿*�^޿�6ӿ~�������`����l�8�x���   �   ,N���-���ս\͈���j�&F����� EZ����f| �r�4��p����a���"ڿe4���9��q������Ș�����ۿb%��E����q�AI5�z� �aZ��>?[��N����k��s��}Խ�,�r���<¾�0�w<-�̼V�Ƹ~����Fힿ�ק��������fU������|��@�W��.�����Hþ�   �   ��-��@׽���8�=�NFc����2�*�����߾��$�L�d����tx������������%��>/�b�2���/�Jl&��s����c�`������^ne�N%�k��Y���Ш+�
���ܼd��A>��Ɂ�l)ֽ��,�ԧ��'����KC�\(5��O���d��Ar�Xw�l�r�jSe�	}P�D�5��aD�&$�� l���   �   <Ľ8I^���|+��un���뽼lV�Eв�Y�
�z�I��ꊿ����"#�v�	��!�ԣ6�h�H���T�r?Y�#U��+I�87�8�!��%
�)��+P�� '���J���
�A���6W������p�x�������]�HEý��� [f��Ԝ� �Ⱦ��u��,%���%��e)��(&�����t����
�ɾ�����g�����   �   �V"�؛��h�����?��<��� ����վ�h$�nm��=��:Dӿ������;���V�޲m�Ƈ}�������}��5n��)W��'<����7�/nӿ�T��Əm�J�$�+-־s]��_d��ӄ�p�ƼH�\���u"�?g���� ��\:��0w�q_�����MBɾf�־��۾^<׾��ɾ帴�p����x�o;����P���   �   ���:�9H<��;,w�����V"��┾+Y���_;�Ln��ı����� ���3��U���u�y@���������4���r���Mv��XU���3�� �쿏���f^��Z;����/���&#�G����5����;��<<�BR:�궼�_�!A���	�52���V���s��c������Α��L�t�ƘW��2���	��4��Xh`������   �   ,��<L��<���<���x���L4�㤾S2�M|M�b���Աƿ�� �	!���D�ʶj��|��@&�����z��������>��҈���j�r_D��� ��w �dƿi����NM��/�����5�����֑�lȅ<h�<�%�<��p<���v�	��7��yw���������'�����_��B��p��N����"�	�`gٻp�y<�   �   ��7=X�*=�v�<� ��;Ω��#@��H���D�Y�S�����пB2��{)�>�O��gy���������0��䀴�N6�����£��*y� SO�j)�Z��usп�Q��9�X��1�u��T�@� ���4���<d�%=fl3=&l=|��< ^/9���O5�]����Ң�L���t������\G���t���5���� *�9 ի<J�=�   �   �q==b�(=<��< 8���k��/�R��޽��-���h������޿��.5�|~_��4��yݞ�+��dU�������V���
���Ӟ�r$��h[_��5���A�޿4���h�ƨ�����.U�_RŽ� ɼ�<�h=Z�4=�Q=D��< �;�����5�0�a� �������򧽹0���ލ��z_�� �X�t��;P��<�#=�   �   �\'=X=��<p���ü�EkN����+D�Kld��F����ڿ ��V2�v<[�_]���Q��5�����#����������M���R���"[�h�1�����ڿmg��Y�d�;��-����P�Y����ʼ���<$�=��=Ts�<�o< -ӻ���2�V�r!��A����ʽҽc�ʽ�N�������S���꼠T���e�<$?=�   �   lY�<��<8aK<(A��M���TB��;��V���UX����!Nп����)�5O�N�x��M���p���������j����~���W��"�x��1O��)�����dпA��f�X��O�iF���?D�F�� aϼ(�'<��<,�<��<Hd���*��)���Ͻ���A2���%���*��%����*u��~ν({���p&���M��z&<�   �   �=�����;�X�:t�ϼ����9F/��������5sE��I��ר���|���p�^O=��Pa�����1��eߜ��������&J������sa��e=����͛��3ο�Dw��:�E�7��z���H1�����߼ A���Ĭ;�» @��D���[Խ�����@�Z�f�w����a������\��C���)�f�S@��Q�޺ҽ*h��Lw��   �   �E@�V���w�����m��5��𷉾���|-�s�y�^`��>�ݿ��
���'�4�E�Fc��5|����6Չ�DΆ��s|�:Qc��F���'���
��ݿ����|<z�c�-��v�喊��N��ڗ��\�d2���U����D�r/��(���I�����ԣ�Ӵ����վ �@���5�վH����ϣ�E����KI�����T���   �   �#ؽt�~��I �@� �Kڇ�D� ���e�u������,�T����h��Cd�����X)��x@�H�S�d
a��e��.a�� T�ʻ@��)����=��TN���M���U�b�������Vg�V������%�$�$�1-��\�ٽ\�*���w�~�����վ ;��C�(%��H/�s�2�/U/� 2%�A]�LR��վB�����w��z*��   �   ��:��
�+��B�\�H���Խ
d8����}X���-��q��ٞ�ȿ�P���P�.��s8�f�;�ґ8��.����4��,l��\ȿ����wq�t<.���4��{9���ֽ�΃�j�_��[�����N;����e¾�����- �Tw?�@[�!q�#�C��� ;�$Lq�Ru[���?�N] �� ��=¾����   �   �4��7�:��W�&:��'���"ͯ�2b��8j�����>�	�}�����ÿ忞@�t���|��#�����^n��p��-ĿNX���A~��?��d��=��Bk�:�+鰽k̆�%�N����:�%
��Q�ξ�6��27��b�:�������"���`��7���Wt���E���ט��g��T�b�Vy7��l�1Ͼ�   �   �j˾�w��(?+��ս����X����Խ�*��)��h�ʾ?�tB��x�Ga��'���ʿ 1ݿ��'�?'��fݿ*�ʿ�j��E����!y��^B�Aa�g˾2u���;+���Խ�~��~Z��L�Խ#�*��,���˾. �8B���x�d��&*����ʿ�4ݿ���*�+鿗jݿ��ʿ�m��ڡ��3&y�JbB��c��   �   �f��@��@k�{��갽nˆ�{�����꽾�:�y��Y�ξb3��.7�C�b�]7������C��!]��ː���p���B���Ԙ�Ke����b��u7��i���ξ�1����:�R�P7�� ����ϯ�e�.=j�q���%�4�>�0�}������ÿ�忄B�����~�,&�����4p�'t忟0Ŀ�Z��XE~��?��   �   �>.���76���9���ֽ�΃��_��V��x��d
;��	��+¾@����) ��r?��:[��q�S�`���x5��Fq�cp[�G�?��Y ��
 ��8¾���:��콟&��h�\����B�Խ2g8�����H\�u�-�?q�ܞ��ȿ�ZR�&����.�`v8���;�>�8�L�.������o�@_ȿ����zq��   �   U����ܹ��jYg���僊�F�%�"�$��&��-zٽ$�*���w�r���w�վ�7��?��%� D/���2��P/��-%�]Y��N�&�վp����w��t*�_ؽ�~�.C ��� �[ۇ�� ��e�������ЬT�F������f�r��|Z)��z@���S�&a���e��1a�4#T��@�ږ)�J�����9P��AO���   �   �>z���-��x����P�Hۗ�Z��&���B��8�D�8&��.����I������ϣ�򮿾g�վL��v��q���վ�����ʣ�򑄾�DI� ��L��,9@�`E����w�����xn������������~-���y��a��<�ݿ��
�Z�'��E��c��8|�x����։��φ�<v|�`Sc��F�,�'���
���ݿ����   �   x��h�E��7��{���I1�O��ȉ߼ 5��P��;���8&�������PԽz��V�@�J�f����@]��g���SX��򒂾G�f�L@��K��ҽP`�� _� ������;���:L�ϼ.����G/�!�������tE��J��6���p~���q��P=�`Ra����I2���������3��UK�����Dua��f=�x��1���FϿ��   �   �A��-�X�P�G��(@D�����^ϼ(<��<��<��<��c��*�"��#�Ͻ����,���%�څ*�u�%�5��Np��uν�s���d&�H�M�@�&<Dd�<��<�gK<�A�������B��<��5���VX�a��+Oп����)�"6O���x��N���q���������i�������X��N�x��2O�<)�:��[eп�   �   �g����d����.����P�J����ʼ躃<��=��=�{�<�3o<��һ����V����𵽞�ʽ�ҽ�ʽ�I������S�ģ� &���n�<�B=
_'=�=��<䦶�#ļ�3lN�E���D�md�VG��A�ڿd���2�=[��]��7R�����y������f��5��N���R�� #[���1�R��6�ڿ�   �   �3����h���������U��QŽ ɼD�<i=ʳ4=�Q=���<��;X����5���a�쓎�������0���ލ��z_��h�t�P�;���<@#=q==��(=��<�9��l����R��޽�
.�ݕh����޿��8.5��~_��4���ݞ�7��kU�������V���
���Ӟ�a$��J[_��5����޿�   �   �f����d�>��-��`�P������ʼ���<^�=��=p|�<�4o<��һ4��j�V����	𵽑�ʽ�ҽ�ʽ�I�� ��x�S�����$��o�<C=�_'=�=x�<����t¼��jN�B���C� ld��F��W�ڿ̯�2�
<[�]��SQ��� ��d������Q��2��*M��=R���![���1����K�ڿ�   �   Q@��,�X��N�"E���=D�\��xVϼ�(<��<��<��<�c���*��!���Ͻ����,���%�Ѕ*�k�%�)��Dp��uν�s��Rd&��~M���&<\f�<<��<�qK<�9��t���7B�
;������TX���hMп���T)�,4O� �x�4M���o���������`����}���V����x��0O��)����cп�   �   5v����E��5�:y��hF1����D~߼ b�� �;���8$������~PԽ^��>�@�6�f����7]��`���MX��풂�8�f�
L@��K�аҽ`��d]�p쎻��;�'�:��ϼ����xD/�|�����rE��H��Ƨ��U{���o�0N=�Oa������/��ޜ�P�������H�������qa�^d=�������̿��   �   :z���-��s������K��՗�4S����$=����D��%�������I�z����ϣ�箿�]�վC��m��h���վ����ʣ�瑄��DI�����K���7@�@����w� |��2i����p������u{-�l�y�_����ݿ��
�x�'�z�E� c�X3|������Ӊ��̆�q|��Nc��F�L�'�h�
��ݿ+����   �   5U�i��ش���Rg�"�~��ܡ%�j�$�R%��Cyٽ��*�y�w�]���e�վ�7��?��%��C/���2��P/��-%�WY��N��վ`���ޠw��t*��ؽ@�~��> ��� ��Շ��� �]�e��������T�������a�p���V)��v@���S��a�D�e�&,a�6T���@�<�)�H�����2L��L���   �   �9.����41��={9���ֽ�ȃ���_�UT�����	;��	��¾,����) ��r?��:[��q�L�]���r5��Fq�]p[�@�?��Y ��
 ��8¾�����:�3�R$���\���Z�Խm`8�����U�|�-��q��מ��ȿ!
��N����.��q8���;�^�8���.����f��i�7Zȿx��9tq��   �   Cb�:���	k��Gⰽ�ņ�򺚽g~��:�E��9�ξX3��.7�<�b�Y7������A��]��Ɛ���p���B���Ԙ�Ie����b��u7��i�~�ξ`1����:��O��3����Aǯ��^��3j�����n��>�7�}�����ÿ���>�r���z��!������xl��m��*Ŀ�U��`=~�P?��   �   �b˾�q���6+�%�Խ�w���S��n�Խ�*��)��@�ʾ3�nB��x�Ea��'���ʿ1ݿ��'�;'��fݿ(�ʿ�j��C����!y��^B�8a��f˾�t���:+���Խ�y���R��ĄԽ��*��&��S�ʾ���B���x��^��$��ıʿ~-ݿ��"#�\#�>cݿ��ʿ�g������<y�[B�H^��   �   �-����:�CI�#0��x����ȯ��`��7j��������>��}�����ÿ応@�t���|��#�����^n��p��-ĿMX���A~��?��d��=��|k����䰽�ņ�8����x꽄�:������ξZ0��*7���b��4���������Y��Z����m���?���ј��b���b��q7��f���ξ�   �   ��:����
����\�� ��x�Խ�b8�����TX���-��q��ٞ�ȿ�P���N�.��s8�b�;�Б8��.����4��-l��\ȿ����wq�n<.����3��k~9��ֽGɃ���_��O����콑;����/
¾ ����% �bn?�6[�Dq���z����/�HAq�Lk[���?��U �L ��3¾����   �   Kؽj�~��6 �� ��Շ�ִ ���e�;������(�T����g��Ed�����X)��x@�H�S�b
a��e��.a�� T�̻@��)����=��UN���M���U�V��~����Ug���;����%��$�����pٽ�*���w�������վ4��;��%�~?/�C�2�&L/�j)%�[U�HK���վR�����w�pn*��   �   �)@��,���w�w���i��$���������|-�s�y�``��?�ݿ��
���'�4�E�Fc��5|����6Չ�DΆ��s|�:Qc��F���'���
��ݿđ��}<z�^�-�zv㾙����M�aח�XR�����,��(�D���b��s�I�,����ʣ�*����վ��㾣�辵�㾀�վ�����ţ�h���#=I����<B���   �   𞎻0;�;@��:�ϼ<���xE/�v������2sE��I��ڨ���|���p�^O=��Pa�����1��dߜ��������%J������sa��e=����Л��5ο�Fw��8�E�7��z�� H1�\��,~߼ ���0:�; j��h��ˁ���FԽt��P�@�X�f������X�������S������$�f��D@��E�~�ҽ�W��XC��   �   �r�<@��<�|K<�7�������B��;��O���UX����"Nп����)�5O�N�x��M���p���������i����~���W��"�x��1O��)�����dпA��f�X��O�IF��?D����|Wϼ�(<�!�<�)�<p�<H�c�z�*����s�Ͻ���'�A�%��*�ĵ%����Dk��lν�k��^W&�8TM��&<�   �   �b'==��<젶�^¼�kN�v��)D�Jld��F����ڿ ��X2�v<[�`]���Q��5�����#����������M���R���"[�j�1�����ڿmg��Y�d�ʾ��-��P�P������ʼd��<��=��=<��<Go< �һ`��d�V�
��
뵽L�ʽ6ҽ��ʽvD��9����S����P򨻌y�<.G=�   �   \�7=\-#=�ߙ<�ļ�ŽJyV�~���Z&�5Uk��즿���Λ��C7��\b��$���M���׵�KH������K��b��_`���@����b���7�����Ῥ��� pl�W0�B�¾�>Z�;�̽�Z��y|<P�=Pb+=��=ʯ<� ";Ĥ��
�!��@m�IZ���3��g���W�������Nh����؈��U�; ��<r�=�   �   ��!=t==�
�<D\Ƽ����� R��̼��6��$g�g���MݿJ:�\4��^��B��ᵝ�����������������Pȱ��ĝ�[��"L^��a4���3�ݿ?���57h�B:����`�U��$ɽ�3���]<X7=g=4��<�F<p�R��d�b�9L��+��ѽC�׽u1н�~��@٘��\� =���"Ỡ�o<��<�   �   �<$��<��0<Lͼ
���l�E�*ر�����Z�A�����ҿ�X�X+���Q��L|� ����
���u��-̶�3t����e����j|�*R��F+�z��y!ӿ�b��g�[�l��ʣ��CI��g��"�g�;�.�<��<@u�;��R7�ޙ���ֽ�����*�)��5.��8)��+�ec���ӽ($��v�.��j��B<�   �   @�ǻ���; �Ը�}߼G���2�����.���G�H��������S���G��?�dyd�̏������_��y6���Y���y�����8�d���?��m�!���G¿Zf����H�j[�t�����5��������@*<� 41;g��L�w`����۽c�fLE�8�k�	.��&�8��뷎�;ń���j���C��]���׽섽�3���   �   ��H���ü������\��E��������/���|�pn���<࿦6�>�)���H��_f����̈����bÈ�����Hf���H��)�JJ��z����ޠ}��w0�$>�,Y���p�[p��P���/���IּʭQ����"���N�v��N���@þ�UپΔ羘k쾉\�Q�ؾ�¾>��������L����tP���   �   �ݽ�����(��V)�������� j�����/��
|W��gq��~`�hx���+�>#C���V��>d��h��+d���V�fC�T�+��n�i�E����#��a�W�L������$l� ��5���~1�D0�5����ὂx/��V}��ݪ��dپ�`����֑'��1�[@5�F�1�EX'��L�B�ҝؾ���o�{�c�-��   �   Dd>������ f��솽�ڽ�2<�-5����V0��Pt���ʿ1���*���!���0���:�\Y>�n�:�X�0���!�2�Q����ʿk����t�N�0�����曾��=�VuݽO���P\k�뭚��O����?�KB�ž*���"��_B��n^��zt�6D�����b2��X9t�`^�� B�\"�����ľ$G���   �   ��R�>�)<��f��s	��!l����,�n��׺�X1
��~A�R���F��&|ƿ�������RW�����G�p��>�����$Oƿ�*��J����A��K
�$��{o����?ٶ��l��	���ڑ�H?�g����_Ҿ���:��f�-$���Ě��W��g����ĵ��k1��
�������Ģe�_�9�A���Ѿ�   �   -eξtÉ� �.��ڽꚽ!嚽��ڽ+�.�ɉ��zξ�e���D�O|�A�������vdͿ�࿒�����{����߿a,Ϳ�_���S���|���D��J�2aξ������.�P�ڽ 隽�暽��ڽA�.�#̉�
ξxh���D��S|����Ě���gͿ��}�����Y��i�߿�/Ϳ�b��FV��|�j�D�@M��   �   (N
�6'��"o�����ڶ��k��X������B?��ܑ��ZҾ����:��e�i!�������T�������������3.�����H1�e���9��=�G�Ѿ�{����>�Y6�d��@	���n�������n�0ۺ��3
� �A�l����H��'ƿ!��������Y�����I�z��������QƿQ-��6����A��   �   ��0�H���蛾l�=��wݽ����Vk������G����?�:덾��ž��ȸ"�T[B��i^�ut�TA��4����/���3t�e^�c�A�TX"�͵���ľ]C���^>����9��"f�톽K�ڽ�5<��7�����X0�8Tt��󠿋�ʿA4���,���!�>�0�2�:��[>���:���0���!���=���ʿf���;�t��   �   ��W�������N'l�@��v����1�<0�ƛ���
�9r/��N}��ت��^پ]����x�'�{�1��;5���1��S'��H����ؾ�����{���-�i�ݽb���ֻ(��T)��������j�{���!���~W������s��!c��y�p�+��%C�p�V��Ad���h�T.d�D�V��C��+�8p�wk�/���K%���   �   �}�iy0�%@�dZ���q��p������#��h6ּ�Q�?v����b�N��z���LþOپ�羹d��U���ؾ�y¾�8��;�����L�2���G��4�H��ü��������]����\�������/�i�|�p���>��7���)���H�8bf�����͈�V���Ĉ�d���Jf�H�H�|�)�bK�\|�\����   �   /g���H�9\�w�����5�+������ �;�`�1;0@��?�X��/�۽ � EE��k��)��鎾;4��O���������j���C��W���׽"䄽T����ǻ�$�; �θ�}߼�����2�v���N����G�\��������U���H���?�*{d�琄�\����`���7��[���z�����Ђd���?��n�����-H¿�   �   c��4�[����s����I��g���缀}�;�7�<0��<P��;و�rE7�>֙���ֽ������l�)��/.�.3)��&�~^�۷ӽ����.���j��`<  �<8��<��0<ͼj���ѩE�Uٱ����Z�᛿ȞҿZY�.+��Q�JN|�ዓ�����v��;Ͷ�6u�����*���,l|�R��G+����6"ӿ�   �   w����7h�u:�Q�����U��$ɽ(2�`�]<�9=\j=���<0'F<��������b�aG���%���ѽ��׽,н�y���Ԙ�؆\�(/�����0�o< ��<�!=�>=��<�]Ƽ�����!R�xͼ�o7�S%g����^Nݿ�:��4�T^�AC��e���±�%���$�������ȱ�Gŝ�_[���L^�b4�8����ݿ�   �   �����ol�(0���¾4>Z���̽�Xἐ||<��=�b+=P�=�ʯ< ";����!��@m�5Z���3��g���W��	����Nh��dو��S�;���< �=��7=�,#=�ޙ<��ļ��Ž�yV�ƙ���&�qUk��즿�����C7��\b��$��N���׵�QH������K��W��P`���@����b�n�7��������   �   ����r6h��9�J���7�U�#ɽ�-� ^<�:=�j=\��<0(F<�������b�OG���%���ѽ��׽,н�y���Ԙ���\��.��0���o<���<��!=�?=h�<XYƼ���h R�t̼��6�C$g�1��qMݿ:�4�@^��B��~���	������	��������Ǳ�_ĝ��Z��zK^�6a4������ݿ�   �   �a��*�[��������_I��d��t����;,;�<`��<���;؈�E7�֙�_�ֽ���~��a�)��/.�$3)�|&�r^�Ƿӽ���̚.�ؒj��c< "�<h��<H1<��̼+���J�E�dױ�w���Z��ߛ��ҿ8X��+��Q��K|�;��� 
���t��˶�%s��
�������i|�
R�F+�ԗ�o ӿ�   �   Ge��A�H�<Z�Ɛ���5�� ��������;���1;�9�v>��W����۽�EE���k��)��t鎾24��F���������j���C��W�p�׽�ㄽ���Ёǻ7�; lǸr߼Q���2�����S����G�u������bR���F��?��wd�ʎ�����.^��5��SX��Jx�� ���pd�Z�?��l�h����E¿�   �   ]�}�v0�j;�5W���m�zk���������0ּ�Q��u�����4�N��z���料@þOپ��羲d��U���ؾ�y¾�8��0����L���>G����H���ü,�����X�����1����從�/���|�m��;࿐5���)�ޕH��]f�4���ʈ�K��������8Ff���H���)�I��x�e����   �   ��W�J�����w l��������<1�470�:����	��q/�\N}�|ت�t^پ]����r�'�u�1��;5���1��S'��H���ڗؾ�����{�E�-���ݽ����.�(�M)�L���$���j�j�������yW���o��!^��v���+�!C�\�V� <d�,�h��(d�.�V�$C�l+�,m�uf����"���   �   ��0�����㛾��=�~nݽ���@Ok�,���F��%�?�덾ۢž����"�J[B��i^�	ut�RA��1����/���3t�`^�]�A�OX"�Ƶ���ľ>C��`^>�2������ f�=熽G�ڽ�.<��2�����S0��Mt��s�ʿ0.��()���!���0�>�:��V>���:��0�ޣ!�^�.	����ʿ9����}t��   �   cI
�T ���uo���CҶ�f������؈�3B?�yܑ��ZҾ���v:���e�f!�������T������	�������/.�����E-�e���9��=�.�Ѿ�{��	�>�(4�`�����!f��v��W�n�QԺ�/
��{A�d����C��Syƿe�(�����$U�X��^E�X��R��;��#Lƿc(��/�����A��   �   �\ξL�����.�f�ڽA⚽�����ڽ*�.��ȉ�qzξte���D�O|�=�������udͿ�࿏�����y�뿽�߿a,Ϳ�_���S���|���D��J�aξl�����.�2�ڽ䚽)ߚ���ڽ��.��ŉ�|vξ�b�j�D��J|���������aͿ+࿲����ￏ����߿�(Ϳ�\���P��|��D��G��   �   �w��Ќ>�d-�\������g�����R�n�f׺�G1
��~A�N���F��$|ƿ�������PW�����G�p��>�����#Oƿ�*��I���	�A��K
��#��Mzo�]���Զ��e������!��=?�ّ��UҾ��� :�k�e��������kQ��������������*�������뇿]�e���9��:�$�Ѿ�   �   bX>�ӱ�
��(�e��憽l�ڽt1<��4������U0��Pt�~��ʿ1���*���!���0���:�\Y>�n�:�X�0���!�2�R����ʿl����t�H�0�Ԝ�x曾ɚ=��qݽ�����Kk������>����?�S獾�ž����"��VB��d^��ot�u>��F����,��a.t�A^���A�XT"�y��f�ľ,?���   �   >zݽt��(�PI)�q���\��?j�������|W��iq��~`�hx���+�@#C���V��>d��h��+d���V�fC�T�+��n�i�G����#��_�W�@�y����#l�������� 1��00�����:�l/��F}��Ӫ��Xپ�Y����&�'��1�75�&�1��O'��D�,����ؾ���e�{���-��   �   ��H�$�ü8押B��Y��-��f������/���|�qn���<࿨6�>�)���H��_f����̈����bÈ�����Hf���H��)�LJ��z����ߠ}��w0��=��X���o��l��
�����$ ּ��Q��l��6���N�~v���ꦾq	þ�HپE���]�O�x�ؾ�s¾�3��������L�����=���   �   3ǻn�; (���n߼���"�2�����!����G�G��������S���G��?�dyd�̏������_��y6���Y���y�����:�d���?��m�#���G¿\f����H�^[�B�����5�'����� ;� "2;�p2��O���۽�>E��k�5%���䎾~/������j�����j���C��Q��׽mۄ�P����   �   �.�<p��<�1<��̼x����E�	ر������Z�A�����ҿ�X�X+���Q��L|�����
���u��-̶�3t����e����j|�,R��F+�|��|!ӿ�b��h�[�f�������I��e��|缠��;�A�<,	�<0��;pĈ��87��Ι���ֽ�!����)��).�n-)�!�hY�îӽ�����.�0hj��<�   �   ��!=B=��<�WƼ����� R��̼��6��$g�h���MݿJ:�^4��^��B��㵝�����������������Qȱ��ĝ�[��$L^��a4���3�ݿB���67h�A:����,�U�+$ɽ(/⼈^<<=Hm=D��<x:F<������b�b��B��� ��Bѽ;�׽�&нXt���Ϙ�~\������8�o<T��<�   �   �=="�(=��<p���y���O��ú�&���	e�٤���[ۿ����a2���[������ɴ���Ӽ�_]��ټ��ȯ�-��y��~a\�,
3�����wܿ_�����f�X9��h��N�S���Ž �Ѽ�L�<=:-=��=���<��t;H9��2��a�hލ�����꥽˞�_^����Z�����Yh�0��;��<�.#=�   �   Y'=�&=$[�<Hu��8帽P�J�b�����f�`��䟿��׿����Y/��W�+��8t���«�ĝ��o������0ͫ�����	>��04X���/��6�3�ؿ�Р���b�wR�������O�����xVҼX�n<d�	=��=��<�W< |������@+X�Ք�Ŵ�c�ȽCvϽL�ǽ�?���4����N���⼰5��LL�<J�=�   �   �E�<�_�<��Q<#���宽߲>��h��G��"U��ᗿ�cͿ����&�"L�$�t�$Ŏ������w�������j��t��=Ȏ��t��eL��'�vn�!Bο�����V����qɮ�#C�I\��(�ּ��<�-�<�%�<���;��v���-�����e+Ͻ������$�`a(�b#����1 ���ʽ�@���!�(�@���-<�   �   �Ot�`��;�
;�qȼ����I,���������B��N��P���:���e��:�� ^�9���]�����������������g���]���:�ʞ�����Q���ue�C��� �u��b80��6����@�����;��D��������fԽ�G�
d?��d�9L��꼊�zލ�n_��
���Qc�p =����}jν�z�L#��   �   p);�]��@l�8A�w���e����F߾�+�vv�9.����ڿ�����%��ZC���_��kx������w��6k��Tx�Z�_��C�R�%����#ۿԏ��Sw�(�+�*ιJ��$M�����������:Ƽ^�G�����M�ȠH�����zf���̽��pӾP?�/����
�ҾZ�������P����E��F
�䃭��   �   �ӽ�y�~,�@���B��&H��;{b��I�������Q�xI���Լ�����	�jq'�4*>�VQ�F�]��6b���]���P�H�=��'�������;ټ��s��DgR�V�G���ae��*��K����&�XW&�@����4ٽ�!*�:8v�F��±Ӿ��������=#�?%-�aw0���,�}�"�������_2Ҿ�ɤ�"Xs��_'��   �   Ъ7�S�罬T��sX������ѽp�5�ݒ���L�Ϸ+��4n�<����ſɒ￶��J����,�N6�>_9���5�),�ހ��w�s���ſ�윿�2n���+�G���R��Ww7��սf?��F�_������뽸�9�����0j��}�����=���X�ln�|��R��Ӿ{���m��(X�β<���������	��`����   �   M쌾�7���䷗�U�o������eg�
���B��є<�G{�il������s��'���lf����7�0��j�3����S��z��`�z��U<�u�߯��B�g�PU�����ƅ�3���P�轰R9������̾���h5�=k`�mᄿ���<N���P��T�����'ꤿy���P^���w_�n�4�c0�l�˾�   �   �\Ⱦ�u��$�(�ҽ"�������aҽ8)�R���9�Ⱦ3���@�7v��ߖ��a����ȿ�ڿ[��6꿎��OڿMȿ�°��T���]u��l?�2��XȾs����(�dҽ1�������Ifҽ2)�[Å���Ⱦ��p@��;v�B▿�d����ȿ��ڿ�^濥:�U濌Sڿ�
ȿ�Ű��W��	bu�p?��4��   �   Bw�貵�5�g��W�|���Ņ�������轞M9����#�̾����d5��f`��ބ����K��KM���P��w��礿�����[��Ps_���4�k-��˾�茾w�7�Q�����sr��M��Yjg�~�������<�c{��n������������vh����9�L��d�������U�����#�z��X<��   �   ��+�����T���y7�$ս"?���_�f��]����9�����e���v��3����=���X��fn�p|�P��<�{�h�m��#X�~�<�5�������������x�7���<P��XoX�����ѽ��5�b����P�h�+�8n�a��n�ſڕ�~��T��2�,��6��a9� �5�H+,�Ђ��y�M��i�ſ��5n��   �   iR���i����e�(,��K��:�&�tO&���+ٽ�*�<0v�A����Ӿ�������H9#�� -��r0�[�,�L�"����~���,Ҿ�Ĥ��Ps�&Z'���ӽjy�&�����C���K���~b�CL�������Q�*K���ּ���b�Bs'�b,>�� Q���]�~9b�V�]��P�X�=�r'�R��Շ�ۼ��t���   �   Uw���+���K��ZN�ᗽ���$���'Ƽ�wG�򜳽�G�n�H�����Na���ƽ�BjӾ�8�|�律��נҾ��������L����E�OA
�m{��$;��L�� l�L?��x���� ���dI߾�
+�txv��/����ڿ���%��\C��_�Dnx����_y���l���x�t�_�PC���%�&��;%ۿ+����   �   F��C�R� �p��g90�37�����@
���:�; �軤���o����\ԽdA��\?��d��G��`����ٍ��Z��ʕ����b���<����`ν��z��㼠�s���;�M
;�qȼ�����K,�0������%�B�P������<���f�@�:�x^�G�������)��S�N��Ϙ���h����]��:����5���d����   �   ����c�V�[��ʮ��#C��\����ּ(�<\6�<P2�<$�;�nv���-�����"Ͻ����^	$��[(��\#�و�,- �=}ʽ�9����!�p�@���-<LP�<�f�<��Q<�#���殽<�>�
j��"��WU��◿�dͿ�����&�0L�~�t��Ŏ������x�������k���t���Ȏ�4�t��fL��'��n��Bο�   �   �Р�J�b��R�⤹�"�O������TҼ��n<Ʊ	=*�=d��<�.W<�I�������"X�OД������Ƚ�pϽ
�ǽ�:��0����N�<��0��<U�<��=~['=�'=\�<�v��=渽9�J���r��$�`�埿��׿"��DZ/���W�����t��Kë�S������A����ͫ�]���S>���4X�B�/��6��ؿ�   �   ;���c�f�(9��h����S��Žl�Ѽ�M�<�=�-=( =T��<��t;�8���1���a�Vލ�����꥽˞�r^����Z�����Zh����;D��<r.#="==��(=��< ���y���O�ĺ�U��(
e������[ۿ����a2���[������Ӵ���Ӽ�_]��ټ��ȯ���j��^a\�
3����]wܿ�   �   Р�>�b��Q�᣹�ΖO�;���LPҼh�n<��	=Ҋ=(��<�/W<�G�������"X�;Д�쿴� �Ƚ�pϽ�ǽ�:��0����N���⼰���U�<�=\'=�(=�^�<tr���丽��J� ������`�X䟿��׿����Y/�~�W�����s��L«�B������.����̫�~����=���3X�|�/�b6���ؿ�   �   H���d�V����.Ȯ�?!C�aY����ּ �<�9�<�4�<`*�;`lv�N�-�٫��c"Ͻ��z��T	$��[(��\#�Έ�"- �'}ʽ�9��!��@�X�-<xR�<�i�< �Q<����㮽ñ>�(h�����]U�bᗿ?cͿx��P�&�LL���t�hĎ�����v�������i��s��eǎ���t��dL�$'��m�Aο�   �   g틿ξC�`� �����50��2��\�� ���0N�; ��l������P\ԽBA��\?���d��G��V����ٍ��Z��ŕ����b���<����`ν�z��	㼠�s�p�;`�
;lfȼ����$H,��������f�B�+N��@���9���d�Ƶ:�D�]�C���7�������������l����f��^�]���:����$��������   �   �Pw�Q�+���H��?J��ۗ�̷�@���"Ƽ�uG�E����G�>�H�t���?a���ƽ�5jӾ�8�s�徃��РҾ��������L����E�'A
��z��r;�<G���k� 2�s����藇��D߾t+�tv��,���ڿ���D�%�&YC���_�,ix�P���xv���i��� x��_��C�Ԩ%�����!ۿA����   �   �dR�a�o���:�d��'�&F����&��J&�d����*ٽl*��/v�A����Ӿ�������@9#�� -��r0�X�,�G�"����~���,Ҿ�Ĥ�wPs��Y'���ӽ��x�n!����@>���B���wb�PG�������Q��G���Ҽ�5��n��o'�&(>��Q���]� 4b��]��P��=��'�\����׼��q���   �   ��+�^���O��s7�:�ԽH9��p�_����ӽ�`�9�e����d��sv��(����=���X��fn�i|�P��8�{�e�m��#X�{�<�/��x�����������7�����M��hX�>v�>�ѽ��5�n���I��+��1n�J��t�ſ����Z����,��6��\9�\�5��&,��~�v�c��o�ſ�ꜿ4/n��   �   �r�.�����g�0Q���6��� ���s���L9�ɻ����̾����d5�}f`��ބ�����J��HM���P��v���椿�����[��Ms_���4�e-�ʴ˾�茾��7�.潣����都j�����ag�Ȍ����ۑ<�{�j������?�⿋���pd�̼��5���b�w��M�'P������B�z��R<��   �   JTȾ�o����(��ҽs�������s^ҽ2)����	�Ⱦ$���@��6v��ߖ��a����ȿ�ڿ[��6꿎��OڿMȿ�°��T���]u��l?�2��XȾ�r��¾(�PҽM���$����Zҽ�)�V���+�Ⱦ���<@��2v��ܖ��^��?�ȿ�ڿ?W��2꿼�NLڿ�ȿ����KR��2Yu��h?�'/��   �   1匾��7��x�𭗽�能�k��&���dg�Ǐ��/��Ĕ<�?{�el������p��&���lf����7�0��j�4����S��y��^�z��U<�u�����|�g��S����#���S������iH9�����y�̾����`5�b`�܄�����G���I��MM�����㤿����Y���n_�Ð4�7*��˾�   �   6�7�u�罳H���bX�tu�V�ѽL�5������L�·+��4n�9����ſƒ￴��J����,�P6�@_9���5�),�����w�u��	�ſ�윿�2n�}�+�"��{R��Fv7�w ս�9��ؖ_��
������9���`��Zp��u��,�=���X�Nan��|�BM����{���m��X���<�P��	������������   �   ��ӽ��x�r����c>��HE��Zzb�kI�������Q�vI���Լ�����	�hq'�6*>�VQ�H�]��6b���]���P�J�=��'�������=ټ��s��@gR�I�����e��)�KG����&�ND&�ޤ���"ٽ�*��(v�D<��ܥӾ����ת�5#�S-�Pn0���,��"��	��w���&Ҿ����|Hs��S'��   �   �;�\4����k��,�+t��������F߾�+� vv�8.����ڿ�����%��ZC���_��kx������w��7k��Vx�\�_��C�R�%����#ۿ֏��Sw�#�+��sJ��L�8ݗ���������Ƽ�iG�哳�0B�B�H�2���@\��)���dӾ2������ྃ�Ҿݭ��r��DH��J�E�=;
��q���   �   `s��;�;`�
; cȼ���"I,�����������B��N��P���:���e��:�� ^�9���^�����������������g���]���:�̞�����S���wc�C�|� �B���70�E4��`�� :��pz�;p�����T����RԽh;��U?�,�d��C��س��CՍ�`V��r�����b�q�<���iVν�rz����   �   �^�<�r�< �Q<����㮽h�>��h��@�� U��ᗿ�cͿ����&�$L�"�t�%Ŏ������w�������j��t��>Ȏ��t��eL��'�xn�#Bο�����V����Sɮ��"C��Z����ּ��<t@�<?�<e�;0Fv�X�-������Ͻ4�<���$�V(��V#�}��7( �Ztʽ�1����!�@�@�0.<�   �   ._'=+=�a�<�p��u丽�J�U�����e�`��䟿��׿����Y/��W�+��7t���«�ĝ��o������1ͫ�����	>��24X���/��6�3�ؿ�Р���b�uR�������O�?����QҼ��n<�	=�=��<pAW<�������X��˔������Ƚ�kϽ��ǽ�5��T+���N�4���ԓ�$`�<8�=�   �   l�L=�W9=���<`7d�y���R)=���i��OV�����iNοd���M'�D�L�>�u�֞��������
���Ź��ꬡ� ׏���v��M��'(��L���Ͽ�י�gRX�l%������B��b���L���*�<��$=��8=� =R�<�O<�j3������A�ttw�Rǌ����'���p�b�7�(!߼`E��XZL<���<��3=�   �   d�7=�m+=h��<�*g�6���09��u����
��wR���@�ʿ|\�D�$�d=I�Hq��������ɩ�����ȩ����8�����q��I�0L%���?̿0���eT��g��t���>��ͬ�������<�_=>h$=�B='�<`>��k¼��7�
d��t��OX���F������C0��0j{��,��[���\�:��<`�=�   �   ��<Ϋ =���<�^t�ט���-�fs��$���LG����%��H�����<�>�N\c�V���ѓ�����cq��ߑ��n���Z��~�c�~<?�J�!i��57¿�v��� I�y��4����2��Ţ�40����]<�6�<x��<@8A<��@���h��4����e��B	�*��M����������I�����t�D[ �@-���~�<�   �   �_);�X<��<��f����������9�5�������������J�2/��O��n��҄�j���R������I����+n���N��,/� ��׉翕���F^��287��V�xn��F!��d��@0��@7y;�<��ֺl�ƼX}d�g������}�/�E�R���n��4��:��Mt���l��`P�x,��^�#Զ��4T�����   �   �7���d��P���5���z�x��*�y�)oϾ���N�f����Lοw� �����
7���P���f� �u���z��Nu�$Df�VP�T�6�"���� �Lο�o����g�e� ��iѾ�}�i�,ᄽ�мh�9��i���'��z���] �jR8��|s�T���a��C�ľ3�Ѿ��վ�ѾK�þ5������o�W|4�2���ꤗ��   �   ��� S�����Tu��4d��[��O�G�������oD�An��<���k�޿\��t�^W2�ԋC�z�N���R�ғN�H�B�Z�1�����\�9�޿����g���`�D��_�g���|�R��,�l�o�t�` ��`�O�½#~�P?c��J���žs����	����`�!�t�$��{!���	���4þ5S��w_�����   �   ^N'��ν(�x�l�4��	Z��d����%�i!����پ4r �xE_�����5V�������n��|'"��*���-���*�ژ!�D��4�0��w˹�IT���!_�P� ���ھK狾�'��G���]b���=�7A��\ Խ5*��(�SᲾ�m��G�sl1��AK�'�_�&Zl��p�%�k�d�^�n5J��G0�}'��X������{��   �   �聾��'���ͽſ���^b��z���A��ָT�h������Po0���k�Hݕ�[�����տ��K��!
��d���	�4��k�"�Կ����@��Y�j�0��{���d���"U������V��f�f��a���ѽĕ)�.��@s��׊���)�qbR��xy���~a��ޣ�㫦�h���ؚ��F���x��Q���(��������   �   �㹾{�u������5��j��X����"���v�έ����s�3���f��Ǎ��㦿n輿�ο��ؿ�xܿO~ؿ�YͿ�
�����J���e�A�2��|�!๾b�u����L���*4���k������Z&���v�ڱ��N���3���f�Iʍ��榿�뼿SοS�ؿa|ܿ߁ؿ]Ϳ���������e���2���   �   ����g��@&U����*X����f�B^���ѽ��)�����n��؇��)��]R�csy� ���o^���ڣ�����C���՚��C���
x��Q��(�<�������偾D�'�S�ͽ ���R^b��|��G��)�T�Tk������]r0�ގk��ߕ�%�����տ�M��#
��f���	����	�%�Կ����"C����j��0��   �   w� ��ھK鋾z�'��I��0]b���=�I<���Խ�/*�\!�uܲ��g�AD�3h1��<K�
~_��Tl���p���k�c�^��0J��C0�$�,S�j���{�WI'�,�ν��x���4��
Z��g����%��#��M ھ�t ��H_������X�����l��P���)"�P�*�0�-���*�ޚ!��F6���࿻͹�V��f$_��   �   ~�D�qa�h ���R�6/���o��p�����`���½Xx��7c��E���	žԳ�;�	���*�!�1�$��w!�+��p	�����þ�N��op_�F���黽4�R�\����p�� d��^� �O�����r��rD��o��;�����޿̹��u�ZY2��C���N� �R�2�N�r�B�<�1�X��^�i�޿u���͓���   �   ��g�ı �\kѾE�}�8j��ᄽ��м��9��W��:�'�r��CX �zK8��ts�t����[��S�ľ��Ѿ��վhѾw�þ���딾�o��u4�����朗�>,���d��-���3��~�z�*��.�y��qϾ�����f�5��&ο�� �"��d7���P���f���u��z�Qu�^Ff� XP��6�`���� ��Mο�p���   �   _��P97�\X�ho��@!�Re��p-��@uy;@,<�pպ�Ƽ�md��z�����ʌ/���R�j�n�d0������k���l�aYP��q,�Y��ʶ��%T�d� �);`"X<��<4�Ȁ�� ��e������5�����&ñ�i���K�h/�(O�h�n��ӄ�����S�� ��R���F-n�
�N��-/�֎�(�翛����   �   zw��YI��y��5��p�2�)Ƣ�$.���^<4?�<D��<hWA<h�����a������\��=	�������������{��G�����t��O � 䥻���<� �<� =���<�_t�Mؘ�.�-�vt������MG������&��HI��`��,�>��]c����ғ�y���Sr��Ē��:��������c�F=?���j���7¿�   �   H0���eT��g��t���>��ͬ�������<�a=Dk$=�F=�0�<`���]¼��7��_��1o��BS���A�������+���a{��+��N���	�:�<��=��7=�n+=`��<�-g��6��d19�^v���
�|xR�y����ʿ�\���$��=I� q�s�������}ʩ�u��?ɩ�	������.�q�h�I�tL%���O?̿�   �   �י�0RX�A%������B�'b��XK��,�<�$=@�8=x� =�R�<(Q<pi3�����A�Ntw�<ǌ����-��&�p���7��!߼ G��HYL<��<8�3=�L=&W9=���<P:d������)=���i��OV�˨���Nοz�� N'�`�L�\�u�䞏�͓�������������߬���֏���v�λM��'(�vL�e�Ͽ�   �   �/���dT�g��s��Ϻ>��ˬ��񜼸!�<�b=�k$="G=�1�< ��(]¼n�7�{_�� o��8S��xA�������+���a{� �+�\N����:��<��=D�7=�o+=���<p%g�b5��*09�ou��f�
��wR������ʿL\��$�=I��
q���������ɩ�q��Aȩ���Ƕ���q�v�I��K%�8�r>̿�   �   3v��t�H�2x��3���2�â�&�� ^<�B�<���<�ZA<ػ����ea�����z\��=	�Ԙ���������i��-�����t��O � ᥻���<�"�<�� =p��<xPt�L՘���-��r������KG�@���!%��9G����v�>�J[c�����Г�����rp�����������D�c��;?����g��>6¿�   �   G]���67��T��l���!�	a��("����y;�5< <պؼƼ�ld�oz�������/���R�R�n�Y0������k���l�QYP��q,��X��ʶ�v%T���`�); +X<P�<�鋼�|�����	��C���5�䡂��������*J�$/�DO��}n��ф�B��aQ�����1����)n��N��+/���@��N����   �   r�g��� ��fѾZ�}�Sf��܄�Dtм�9�HR��X�'�hq��X �DK8�Xts�b����[��F�ľ�Ѿx�վaѾq�þ���딾��o��u4�l���t����*�h�d����0'����z�T��T�y�,mϾ���e�f�y���οz� ����.	7���P�\�f���u���z�Lu��Af�TP���6����g� �6Jο3n���   �   ��D�^�������R��&���o�fi�0���`���½�w��7c��E���	ž���2�	���$�!�+�$��w!�(��l	���쾾þ�N��Jp_����軽x�R�t���4c��d�c��V���O�
�����|mD��l��u���;�޿��lr�|U2���C��N��R�j�N��B�b�1���>[�ʟ޿����ɐ���   �   я �/�ھ�䋾�'�PA���Qb���=��9��$Խ/*�!�Sܲ��g�5D�*h1��<K�~_��Tl���p���k�`�^��0J��C0��#�!S�Y����{��H'���νX�x���4���Y�._����%�����پp ��B_������S��f��,�����v%"���*���-�T�*�ʖ!�d�
3�M��ɹ�AR��D_��   �   �v��la��eU����P����f��Z��eѽG�)����vn��ȇ�Խ)��]R�Zsy��m^���ڣ�����B���՚��C���
x��Q��(�5�������偾��'�F�ͽչ���Sb��t��	;��W�T� e�������l0�d�k�ە�������տ��I��
��b���	�N������ԿY����>��v�j���/��   �   �۹��u��~������-��(e��0����!�,�v�������g�3���f��Ǎ��㦿k輿�ο��ؿ�xܿP~ؿ�YͿ�
�����K��	�e�?�2��|��߹���u�Ă�W���y/��hd��ڢ��i�'�v������)�3���f�Jō��িK弿sο!�ؿuܿ�zؿ?VͿ����������e���2��y��   �   #⁾٬'� �ͽS����Qb�Jv��"?����T��g������Co0��k�Cݕ�W�����տ��K��!
��d���	�6��n�$�Կ ����@��Y�j� 0�n{���d���!U�6����R����f�?X��0ѽ�)�t
��9j�����R�)��YR�pny�;퍿n[���ף�x������Қ��@���x�:
Q�T�(�7�������   �   jC'��νf�x���4�(�Y�a����%�!����پ$r �nE_�����1V�������l��z'"��*���-���*�ܘ!�F��4�4��x˹�KT���!_�G� ���ھ 狾�'�]D��.Sb�8�=��5��`Խ**���ײ��a쾵@�d1�D8K��x_��Ol�&�p���k�H�^�,J�L?0�X �M����V�{��   �   P໽j�R�\����[����c��X�0�O��������oD�=n��9���h�޿Z��t�^W2�ԋC�|�N���R�ԓN�L�B�\�1�����\�:�޿����h���]�D��_�1�����R�9*��o��g�2�� `���½�r�w0c�]A��sž\��	�����!���$��s!�#���	���þ�I���h_�9���   �   ��p�d�@���\"��b�z�l����y��nϾ��G�f����Jοv� �����
7���P���f� �u���z��Nu�&Df� VP�X�6�$���� �Lο�o����g�_� �^iѾo�}�h��݄��rмȬ9�C��ַ'�|i���R ��D8�Vls�����:V��o�ľ��Ѿ*�վ*Ѿ��þf뮾甾��o��n4�H���ɓ���   �   @�*;�DX<��<X拼}��Ղ��
�����3�5�������������J�0/��O��n��҄�i���R������J����+n���N��,/���ډ翙���H^��187��V�In���!��b��P"����y;�J<@<Ժ��Ƽf^d�Pq�� ��4�/�S�R�P�n�,�����Bc�l�l��QP��j,�7S�0����T�hؤ��   �   `.�<ȴ =|��<XLt��՘�o�-�Ds�����LG������%��H�����:�>�N\c�U���ѓ�����cq��ߑ��n���[����c��<?�J�#i��97¿�v��� I�y��4��_�2�\Ģ�4'���^<�H�<p��<xvA<ȗ�L���Z���w��vS��8	�������`��������w��F�t�xC �����x��<�   �   :�7=�q+=���<�!g�K5��P09��u����
��wR���A�ʿ|\�D�$�b=I�Hq��������ɩ�����ȩ����9�����q��I�0L%���?̿0���eT��g��t����>��̬�,�@"�<�c=n$=NJ=�9�<���dP¼��7�?[��zj��TN��k<�������&���X{���+�t@�����:h�<��=�   �   Z^e=<�S=b&
=`0�;����t"�|q��J��|�@�+承]��Ht���6K8��[�̕}��ލ��3���ߛ�x9��z���|~�n�[��9�Fd�e�����
"����B�����͛���(�Z������\]�<NF:=0WL=R6=:�=tS�<�Һ�ќ�$ ��{?��B^�Log��Z��Q7��1� O}� �6;�R�<|`=�aN=�   �   GR=��F=�J=��;�|�����L���k���=�����{������&5�V�V��{x��׊�zٔ�{f��0ؔ����F�x���W�>�5�.��d�Z��6����?�<���C����%��7����t��<��-=�9=��=Dh�<���;��Y������K��A��O���v��O3��2Tz�~	@��R�m���:<���<��4=�   �   ��=�b=���<�ao���n�6���:��VS�r�2������{L��),�FvK��j��Q���e�������S���>��^j���K�,����s�9&��͜���4���S<��`V�� ��@g��>�<�=�X =��< ��7�z¼ *J��F����Ž�1�^���9�GX��������ǐ���8��횼 ��;��<�   �   p|J<�<���<@U����V������|��qӾA#�j�k�f���G�ѿ���t��C:���T��k�b{�@8����z��6k�F�T�z":�$��J��Nҿ����8m�6o$�D&־�ှ�
��k�X\2�h�F<Z�<��;0�`��V.�@՜�?�潐����7�B�P���`���e���_��N���4����V2޽�B��N������   �   ��ż�W>� L>;��%�f=���r�Y��췾���q�O�q⎿�캿6꿾p��y%���;�tN��Z��+_�l�Z�\�M��@;�
%��=��3�0���M����P������^^�|�HO��n� �޺ |���케U���ٽ(��KU�z܄��8��瞮��K��������k��]����߂�8�P�~��[vϽ�#m��   �   �ϗ���$��p,���C)�/3��?�3��G���g�e0�ot�Q�q�ʿ������"_!�8V0�\:�i=��9�޵/�8� �VQ�����ʿ�נ���t�>�0�ǫ񾸵��.�6���½<7��ű��S���e)�'T���(�XzF�I3�����B�Ծe���b��*��Ͷ�������&����Ҿ����܅��A�
� ��   �   ���GZ���j<������ �#������t���������H��e��u�XͿ\��� ���:��R��m�4y��W��P!̿�V��
��˾H���p3¾p�u����2����*��k	��[H��㯽�k���_�!|��=�Ҿ��;���6��3I���T���X�(fT��OH��5�
���n�5[о�H��z�[��   �   �c��U��㨽X�J���(���p�geսQ�8�o���ǟ߾B��8T����}���
¿oۿ�������s����`��p��c�ٿ6���^���҆��TS�`��� ߾4�����8�u�ֽ\u�<K.�2(Q��۬�x����e�m쨾v 龂?�lI=�k�`�p:�������B���͖���틿 �~�en_��;�v�����Y-���   �   i����V���6���F�D���E�p����z���W��h��ݰ�T!�yP����
��IH��������ĿȿMoĿn7���Y���)����~�n�N��Q �#=쾱e���V����񗽜�D���E�c����}��W�Bl��ҵ��W!�mP�B�����AK��������Ŀ_ȿ�rĿ�:��b\��^,��*�~��N�~T ��A��   �   e$߾͙����8�O�ֽ*u��I.��!Q��լ� ��l�e�:訾�<�\E=���`��7������?��
˖�:퓿닿�~��i_�>�;�F�����z)��c�R��ި�t�J�p�(��p�jս>�8�a����߾�D�y<T���������¿�ۿ$��������d��Ϣ�|�ٿ������Ԇ�XS����   �   ���76¾�u���������*�:g	��RH��ܯ��f��_��w����Ҿ���%7���6�'/I���T���X�XaT�KH�ܓ5�T���k��Uо�D��*�[�����S��.c<� ��T� ��%��,���t����ʥ���H��g�����Ϳe�ￌ�z�0��T��o��z�6Y��S�&$̿�X�����n�H��   �   -�0���񾌷��d�6���½�<7�����PF�� [)�YL��P#��sF�/�����=�Ծ�������V����ˍ�������@�Ҿ.����؅���A� � �oȗ������t(��BE)�,6���3��I���j�Og0� rt�'��ʿ����<���`!�(X0�p!:�<k=���9���/�޲ ��R�J���ʿd٠�!�t��   �   ��P�������q^�'~�.O���n���ݺ ;����켜M��bٽ�|�wCU�؄��3������'F�����}����e������>ۂ���P�z���lϽm�4�ż��=�`�>;�%�Xh=�!��.�Y��<����O��㎿S8��q�d{%�B�;�vN�2�Z��-_���Z�>�M�rB;�d%��>��5�}1���N���   �   �m�:p$��'־\‾�
��k�W2�x�F<�e�<pH�;��`�JH.�x̜����v����7���P���`���e��_���N���4�ۻ�F(޽K:�����0y�p�J<��<ԕ�<�S��Z�V���(�|��sӾ�#�:�k�������ѿ���u�:E:�4�T��k�^{�C9����z��8k���T��#:����J�*Pҿ麡��   �   G�����4�ӌ��<���V�� ��Xc�hC�<֗=^ =��< ��7Dd¼�J�2?��:�Žt(��u���4��N�����ϱ��V���8�8��ؚ�0լ;���<��=�e=t��<�fo��n�]���;���T�z�2�t���w���M㿬��),�LwK��j��R���f��{���zT��}?��zj���K�p�,�����t��&���   �   g����?�����p����%��7����0��<��-=Χ9=|�=Xq�<���;��Y�R��j�K��=��kJ��Sr���.���Kz��@�E�HU��;<���<�4=2IR=8�F=>K= �;�&��}���L���l���=������=����'5���V�P|x�؊��ٔ��f���ؔ�W����x��W���5�h�����Z���   �   �!��[�B������̛�G�(�ހ������^�<�F:=�WL=nR6=��=T�<@�Ѻlќ�����{?��B^�@og��Z��Q7��1��O}��6;@R�<0`=naN=^e=޼S=�%
=�0������t"��q��cJ����@�J承���ot�,��NK8��[��}��ލ��3���ߛ�t9��q���f~�V�[��9�0d�?��ꄼ��   �   ʱ���?�I��������%�56���
�؍�<��-=d�9=��=�q�<��;��Y���J�K�~=��ZJ��Hr���.���Kz��@��D�T�8;<(��<L�4=�IR=�F=lL=��;�<��^���K���k���=�s���;��A��D�:&5���V�{x�A׊�ٔ�f���ה������x��W���5������Z���   �   ����4�d��:;���T�!���XT�hH�<��=._ =��< �7(c¼HJ��>���ŽT(齤u���4��N����佾���>����8� ؚ�@ج;��<��=�f=���<�-o�x�n�:��;:��eR���2�L�������K�~�^(,�juK��j�UQ��)e��㘎��R��>��j���K��,�f���r�W%���   �   cm��m$�H$־����
���k�0B2���F<Xj�<�U�;��`�VG.�̜�g��R����7���P���`���e��_���N��4�ͻ�#(޽ :��~�� v���J<�<H��<0,����V� ����|�0pӾ; #��k�y����ѿ��s��B:�,�T�\�k�r{�;7����z�&5k���T�*!:���2I��Mҿ͸���   �   ��P�&��� ��^��v콴O��vn�@uݺ�$������L���ٽ�|�GCU��ׄ��3��t���F�����v����e������5ۂ���P�b���lϽ$m�0�ż@�=���>;pm%�B_=�����Y��귾j����O�JᎿ,뺿<4꿤o��x%���;�*rN���Z��)_�L�Z�h�M�?;��%�~<��1�Q.��OL���   �   ��0�f��D�����6�;�½627� ���0=���W)�PK���"�4sF��.�����%�Ծ�������P����ƍ�������:�Ҿ$����؅�q�A�� ��Ǘ�b�T�����X;)��.��F�3��E���d�c0�}lt��렿n~ʿ����H��z]!�ZT0�R:�g=��9��/�|� ��O�E���ʿ�ՠ���t��   �   ���0¾��u���>~��(�*�H`	�nNH�Tۯ�f���_��w����Ҿ���7���6�/I���T���X�SaT�KH�ٓ5�R���k��Uо�D���[�����R��_<�4���H� ����b��dt���������H�Bd��`�Ϳ}��8����P��P��k�^w��U��M�̿nT��.��ӻH��   �   e߾�����8�9�ֽ6u��?.�`Q��Ӭ�h����e�訾��<�OE=���`��7������?��˖�9퓿닿�~��i_�<�;�A��y��b)���c�zQ��ܨ�V�J���(�r�p�!_ս-�8������߾�?��5T�w}���z���¿OۿF��k�������b]�����0�ٿS���Ҏ���φ�DQS�����   �   �a��,V����&뗽��D���E�u����y�B�W�^h�����T!�kP������FH��������ĿȿNoĿo7���Y���)����~�m�N��Q �=쾐e��h�V�0��:��D�6�E�n񘽭v���W�e��2��Q!��P����u��fE��e���H�Ŀ�ȿlĿE4���V��''���~�|�N�SN �8��   �   p�b�M�ר��zJ���(���p��bսz�8�+�����߾B��8T�z��}���
¿kۿ�������s����`��q��g�ٿ9���^���҆��TS�\��� ߾ �����8��ֽ�	u��?.��Q��ά����X�e�4䨾���8�rA=�0�`�J5��}��=��Ȗ�R꓿K苿��~�De_�/�;������-%���   �   ����K���U<������� ����t���
t���������H��e��o�RͿW��� ���<��R��m�6y��W��P!̿�V����ʾH����N3¾�u�������H�*�J]	�GH�,կ��a�B�_�qs��^�Ҿ���b3�N�6��*I��T���X�w\T�nFH���5�{��Vh�pPо,@��$�[��   �   ɿ��Z��l�����v;)��0��g�3�uG��bg�e0�ot�L�k�ʿ������ _!�6V0�\:� i=���9��/�:� �XQ�����ʿ�נ���t�<�0���񾃵��n�6�`�½<47�����X2��|N)�CD����lF��*������W�Ծ�~�����������r��՗��<�Ҿ ����ԅ���A��� ��   �   ��ż�9=�@?;�d%��_=�����Y�d췾���i�O�n⎿�캿6꿼p��y%���;�
tN��Z��+_�n�Z�^�M��@;�%��=��3�0���M����P��������^�1z�<O�tn���ܺ���̞켭E��Yٽ�v�<U��ӄ��.��'����@��'��ѝ��i`�������ւ�J�P���WbϽPm��   �    �J<��<t��<� ��t�V����I�|��qӾ9#�f�k�b���E�ѿ���t��C:���T��k�`{�?8����z��6k�H�T�z":�&��J��Nҿ����:m�3o$�0&־VှB
���k��B2���F<�s�<���;hc`�&:.��Ü�_��t����7�|�P��`���e�7�_�-�N��4�����޽\1��0��HI��   �   �=�j=̵�<�o���n�Ć��:��ES�n�2��������yL� �),�DvK��j��Q���e�������S���>��^j���K�ė,����s�;&��Μ���4���8<���U�R���`V��J�<b�=�c =+�< `8�N¼�J��7��؜ŽT�-l���/�$E�����J��������t8��� �;p��<�   �   �LR=
�F=�M=@�;�"�����L���k���=�����z�����~��&5�T�V��{x��׊�yٔ�{f��0ؔ����F�x���W�@�5�.��e�Z��7����?�6���8����%�7����l��<��-=d�9=��=�y�<`��;��Y�B����K�H9���E���m��6*���Bz���?�46�;��!;<L�<�4=�   �   e�=�'v=�v4=�F><�/��U��j~�o�־��%��[o��]���{Կ�� � �V�<��ZX�"�o����G���r��dp��X�Xy=�:!�Vz���տ魤���q��'���ھ�ނ�w��f�M� �u;B�=��S=�c=PP=J$=4�<�#<@Ĳ��f��T����HB�Ҁ��wݼ�Yz� ��0p�<\q=��B=0�p=�   �   ܧt=��j=�@.=�5;<��)��_����x�Ҿc�"�')k�ƣ��vѿ��� ���9�.XT��<k���z��;��<�z�"Ok�f�T�X:�v��rJ��dҿfޡ��\m���$��,־|��Jh�D�G��as;$]=�I=�>S=b�9=N5=݋< ����p������4� R�lXZ���L���)�D�꼈M� >�;���<ʊ%=��Y=�   �   �L@=2G=.�=��.<X�fV꽘i�"0ƾ�����^�ְ��(ǿy���_��X0���H���]��l��q�"�k�^�]���H���0�$��o���t ȿ±����`������ɾ��o�8���S7�`�];@z�< E'=� =$?�<PW:<���t��~�]��ϖ�OԵ��$ɽ��νvƽՖ��
5����J�qټ`~P�p%�<8h=�   �   @��<fN	=�'�<@�<�>��Ͻ��P���>��8�K��/��fm����応�
�<3"�R8��0J�(_V�̘Z�r%V��I�
�7�Z"���
�;?�i���⌿5M�%9��ٵ�~oV�b�ڽ�����;졷<���<�X�<�Z8�|�ּdVf��L��0����/�+���9��>�Ff8�lM)�B*��-�1���hM�4۠��P�;�   �   0���@�6<�a�<@՘;���L����m2�� ���M��RY3��Nx��H��8AͿ%������#���2���<��A@���<�fN2�t#�x\������>Ϳׄ���y�bF4��T��J*��V7������� ���(<�/�;X�d���3�2��*� �00�v�]�R]���j��蒝�yԠ��ݜ����:v���5Y�Ҧ*����������   �   �5U�\6��`���*� ����X���1��8��̾A����S�'0��$��Z�ֿ���$5�6���"�L�$��!�2[���������տ�ɰ���� �S�1"�H�;��������4ἠ��Pm��ʼ�=k�|ӽ�"�T�c��ޓ�����)mҾΝ�<R��������{ ��bоC���65��(4^��Q���ǽ�   �   k����t�T�༰�g� E��V���߽@�I���������Z-�Ǎg�CQ���h����ѿ���	� �:���	��:�4\ �A�뿅�п�������f�p -������3���[K��佄N`�x{ɼh���L����₽����8��R������ۿ��g��-���7��@;�j7�)�,�.<�|k�c<�Hi������b4��   �   ��:�9*⽈u�T
��dg��f� �������:�x�'������U7�$Lk�q@�������Ͽ��ѿ��ۿc�߿�vۿ�6п�ƾ������c���i�	q6��A�m{��ax���H٣��y%�@�μ|��Xp��;��>��^��k�ƾ���)#�z�B�h^�Y t�t뀿�*��$����s��\�A���!�aC�zFľW���   �   ������/�;3̽�KX��l��dm���I[���ν��1�:-����ʾێ
�{�3�3^�)z��:`��0N������鯫�䛢�����������\��\2��	���Ⱦ������/��-̽6FX��i���r���P[���ν �1�r0���ʾ��
���3�37^��|���b��Q��p������в������
���񗂿s�\�)`2�{�	���Ⱦ�   �   �~���ex���ܣ�x|%���μ��xf�R4�m>��Z����ƾ"��U&#�W�B�gc^�dt��耿�'�������s���\�A�Y�!��@�Bľ�S����:�Q#��	u�����f��� ��������b�x��������X7��Ok��B��'����ҿ��ѿ��ۿ��߿�yۿ�9пfɾ�����e��j��s6�7D��   �   E���g6���^K�v��Q`��zɼ`���x����܂�S����8�O��0��D��v���c�Қ-�~�7��<;��e7�#�,�}8�:h��6ྵd��X����
4�O�ཾ�t���༠�g��F���V�|�߽�I�v������B]-��g�CS���j����ѿ��쿤� �����	��<��] ����п�����Ò���f��"-��   �   �#���;,����������`�� =��ʼ�/k�>ӽ�"�غc�
ړ�B�=gҾe�龁K��%��E���0�]о/����0��
-^��K���ǽ�(U� %����`�*�츾�v[��n4��:����̾9��6�S��1��&����ֿ�����6�����"��$���!��\�$��`�����տx˰�V��G�S��   �   �G4�W���+��&7��������Ń�А(<0i�;��d���3�;���� ���/���]��X���e��􍝾uϠ��؜�����q��L.Y�o�*����������	� �����6<�h�<�ۘ;������,p2����KP��-[3�)Qx�`J��
CͿI�����#���2�j�<�XC@�f�<��O2��#��]�����u@Ϳ(����y��   �   L6M�
:��ڵ��pV���ڽؠ���;��<���<|g�<��5�H�ּ�Ff��C��w������+�ϸ9��>��_8�
G)�l$��#� (���YM�|à����;���<�R	=4,�<ؽ<�@� ϽͼP����i����K��0���n���忆�
�R4"��8�2J��`V�d�Z��&V�~�I�8�7�V"���
��@�y��㌿�   �   ��`�*��`�ɾ�o�<����S7���];h~�<�H'=�� =�K�<�w:<������]�!Ȗ�9̵�wɽ/�ν�mƽ쎰��-���wJ��Zټ �O�t4�<n=�P@=�G=l�=��.<P�jX�Fi�i1ƾ�����^�����ǿ�����_��Y0���H���]��l�.q�P�k�l�]���H�<�0����Y���-!ȿR����   �   B]m��$�-־���mh�,�G� ms;`^=|I=AS=��9=b9=��< ���c�����D�4���Q�8PZ���L��)�p��(�L�`h�;���<N�%=T�Y=��t=��j=A.=�3;<�)��`����x���Ҿ�"��)k�?���ѿ���f����9��XT�>=k���z��;����z��Ok�ؗT��:�����J�Aeҿ�ޡ��   �   ŭq���'�i�ھ�ނ�.����M���u;��=�S=t�c=�P=�$=��<h�#< ²�(f�������:B�Ԁ�$xݼZz�����o�<0q=��B=��p==�=4'v=Hv4=@D><�/��U�@k~���־�%��[o�	^���{Կ"��4� �j�<��ZX�0�o����G���o��Xp�ֲX�Fy=��9!�Dz�e�տɭ���   �   ,\m��$��+־���fg�|�G�`�s;�_=HI=�AS=�9=�9=��< ���Pc������4���Q� PZ���L���)�4�꼐�L��i�;(��<|�%=��Y=6�t=~�j="B.=`:;<��)��^��T�x�u�Ҿ'�"��(k�����)ѿV�����ƨ9��WT�<k�F�z�-;����z�|Nk�ҖT��:���J�^dҿ�ݡ��   �   ��`����;ɾ
�o�Y���nN7���]; ��<$J'=� =�M�<xz:<ؤ�.����]��ǖ�̵�Xɽ�ν�mƽ׎���-���wJ�pZټ �O�45�<�n=�Q@=2G=��=p�.<^��T�ii�K/ƾ@����^�G���qǿ����~^� X0���H���]�vl��q���k�:�]���H���0�p��D���|ȿ�����   �   l3M��7��׵��lV���ڽ���`";���<���<�j�<��5�L�ּ
Ff�&C��#������+���9��>�u_8��F)�\$�z#��'��HYM�� �`��;���<�T	=$2�<��<:���νԸP����U����K�/��Xl��C��ж
�B2"�$8�L/J��]V�2�Z��#V���I�Ļ7�B"���
��=����ጿ�   �   �D4�R��C(��_7�S���8�����h�(<�;�d�@�3����_� �M�/���]��X���e��獝�iϠ��؜�����q��=.Y�Y�*�����F������|����6<�o�<��;H�༾���wk2����RK���W3��Lx��G���?Ϳ5��|��>~#�f�2��<��?@��<��L2�#�8[�m���=ͿS���Sy��   �   / �Q�;h��������D�� �� ��ʼ�-k�pӽ��"���c��ٓ�&�&gҾQ��rK����8���'�]о&����0���,^��K�t�ǽb'U�D ���x��F*�����T��W/�7��:�̾���S�S��.��A"��6�ֿ�����3����"���$�2�!��Y�@��C���G�տ�ǰ�?��b�S��   �   ����1��PWK���C`��gɼ����ؗ��ۂ�<��n�8��N����#��h���c�Ț-�v�7��<;��e7� �,�z8�7h��6ྪd��H����
4����b�t��� �g�t4���V�8�߽|�I��������NX-���g�fO��Uf��[�ѿ��x� ����@�	�R9��Z �O����п*������G�f��-��   �   �w��z[x�����ң��n%�4�μ��Hb��2��>��Z��}�ƾ��D&#�I�B�Zc^�Yt��耿�'�������s���\�A�W�!��@��Aľ�S��f�:�="�Bu�P���PU��� ����k��6�x����G���R7��Hk�I>�����
Ϳ��ѿt�ۿ+�߿�sۿ�3п�þ�����a����i��m6��?��   �   x�|�/�I&̽�9X�T���\��D[�Ưν�1�-��f�ʾȎ
�j�3��2^�"z��4`��+N��|����篫�团�����������\��\2��	���Ⱦ�����/�h,̽*AX��Y��xZ���>[���ν��1�!*��s�ʾ1�
�,�3�/^��w���]��hK����������������P���j�\�oY2�}	���Ⱦ�   �   �:���
�t������Q��� �%���L����x����x���U7�Lk�i@�������Ͽ��ѿ��ۿb�߿�vۿ�6п�ƾ������c����i�q6��A�S{���`x�h��ף�s%�H�μ���Z�2,�>�GW���ƾB���"#�R�B��^^�~t�L怿\%�������r��\��A�Ȧ!��=�2=ľ�O���   �   �����t�Й��g��2���V���߽��I�v��������Z-���g�:Q���h����ѿ��� �:���	��:�6\ �E�뿉�п�������f�n -������3��&[K����H`��iɼX���Њ���Ղ�O����8�TK��z�����%��?`���-�3�7�.8;�ra7��,��4��d��0��_��j����4��   �   ~U����@� *�@���cV��41��8����̾2����S� 0��$��S�ֿ��� 5�4���"�J�$��!�4[���������տ�ɰ�����S�."�3�;`���c�������༐�������ʼF!k���ҽ �"�z�c��Փ�봾daҾ���D��L���z����$Wо�}��Z,��u%^��E�!�ǽ�   �   �(��07<y�<�;`��r���2m2�� ��|M��FY3��Nx��H��2AͿ������#���2���<��A@���<�hN2�x#�z\������>Ϳڄ���y�aF4��T��(*���7�#�����@�����(<�;@�d���3�T
��"� ���/��]��T��Ja�����hʠ��Ӝ�6���m���&Y���*�����Q�������   �   ���<�Y	=�8�<��<�:�3Ͻ?�P����3��0�K��/��cm����忘�
�83"�L8��0J�$_V�ʘZ�r%V� �I��7�Z"���
�??�m���⌿5M� 9��ٵ�*oV�5�ڽ ��@!;���<ԣ�<�w�< [3��ּ|7f�Y:��ڍ����3�+� �9�� >��X8��@)�b��꽻���IM�,������;�   �   �V@=�G=��=�.<���U�Ui�0ƾ�����^�Ұ��#ǿt���_��X0���H���]��l��q�"�k�^�]���H���0�$��q���u ȿñ����`������ɾĨo�|����P7���];$��<�L'=� =�X�<x�:<`��:����]�����-ĵ�ɽ��ν)eƽ̆��>&��^jJ� Cټ�GO�pE�<�t=�   �   ��t=L�j=hC.=@=;<j�)�_����x���Ҿ_�"�$)k�ģ��uѿ�������9�.XT��<k���z��;��:�z�"Ok�f�T�X:�x��rJ��dҿgޡ��\m���$��,־q��h��G�@�s;�_=NI=vCS=��9===��< c��@W�������4���Q�HZ���L�P�)��꼠�L����;���<��%=��Y=�   �   �ԕ=��=�9e=�g�<0������F�򈭾�G�wG�-���k�����n�����r�3��E�<�Q���U��Q���E��&4�R���.�u��.����+��H"I�FF
�v����XO�L�˽��H��<n�4=��k=*�x=��g=�B=|=䂵<<< �
�/1��?��`�Sh���껀iY;`�<���<�:=�p=���=�   �   2X�=��=�_=���<�3��Nг�^4B�&�������yC������z��c2ݿ���@���0�*-B�X�M���Q�f�M��:B��1��U���+;޿��������rE�q��1ڭ�́J�ƽd1�h�<0=��b=��j=6�T=��)=�N�<�=Z< T{��A]�䚽�4C�����d޼������Я�;�[�<�`=�#W=���=�   �   x�n=��t=r~N=��<p�s�㧤���4������?���9�9���姿��ҿ�|��p���(�N8���B���F���B�N
8�@(��������|ӿs��������:�\���� ��B�<�έ���żp�<��!=4;F=n�?=�)=�¼<��;��b��f��G��z�&1��ks�������l�#2���Ѽ*��Xp<$8	=�G=�   �   |: =X�>=0�/=�s�<�/�����"j ��}�����K�(��Lj��b��Q¿&��D	�����(�Ja2���5��82�ο(�<|����:�S�¿暿�~k�*�o��|��'��М�����%�<
G=Θ=�<tR<������z {�Tֲ�c ��c�4���7�D$�4	 ��#ؽ
��\���Ҽ��$:��<�   �   �3<�O�<� =��<`�ϻ$d�����zv�a�ƾ�����N�V��3����ѿ����l
��{����d7!��J��#��	��u��d�ѿy3��?:���|O����R�Ⱦ�&{�[��=}� ][�H]<��<��< ��:��¼��f��@��k�
.�}WP�y?k��/|�~�����z��	h��K�Q(�kW �A����C�x�r��   �   ��߼ �:�y<�ns< �F�`�)�~�ս)bI�]W������N�/�jVj�����F���Կ�� !�L��($�`��ȼ�,Bӿ羴�!����3j��/�W���P����L���ݽ$J=���g<@X<��0	��2��8���$3��dl�����ڪ�{\����ʾ�ξb�ɾ����m���;��+�e���+�؏�﬇��   �   6i���,�@�ػ�j�; �����q�_�ゾ�ZȾB��o�@�|�v�s斿O/��?2ȿڿ�q��,�& �ZٿLǿ�U���7��h�u�P�?����H]Ⱦ&M��N������� �0��� �X�@�B� �#��ʩ�����S�A}��q޸�{ �f�� @���@��p~�|d��X ��Sݾ|ε�JM���EM�<1��   �   =���������"�p1������mT�5߽��C�	V���O޾�w���C��Oq�s��|����l���ʹ�޼��h��y���깠������o�M�B����cݾ����&�B��߽�W�����p�ǻ`�Q��D��e��w��(�b�H٠�0�վ�g��!���8�uGK� W�^�Z��yV�5MJ��s7���7����Ҿ�"��ˢ]��   �   ��Y�V�N��T��He�x�"�����ʿ��^����\�[��[�\l�W�8�rf[�z�������
���>��/o��̜x�L�Y�g7�������#����Y������`���_��"������Đ�4��.�\����Qo��8��j[��z��������k��pA���q��*�x�/�Y��7�����['���   �   [����B��	߽�W����p�ǻ�xQ�&<�5_������b�@ՠ�&�վ�d�B!���8�7CK���V���Z�7uV�IJ�(p7����V��0�Ҿ-���]� ��������!�P.�����tT��:߽��C�Y���S޾0z�G�C��Sq�Ju������no��N͹��༿8k�����I���8�����o�[�B���+ݾ�   �   4`Ⱦ5O��
��]���p� �𘿻  #���B���#�:é����l�S�,y���ٸ���-���<�]������z�a��U �mNݾ�ɵ�iI��~?M��,�Nb���"���ػ`��;������Z���@b�x傾0^Ⱦu��@�@��v�{薿�1���4ȿ� ڿ[t��/����\ٿ�Nǿ�W���9����u���?�����   �   >���\���֕L�%�ݽdM=�@�0p<�l<p�Ệ��+������3�!]l�|	���ժ�W��I�ʾ%�ξ��ɾ���������6����e���+�3�齃����߼ �:��y<xus<@G���)���սkeI��Y�������/�6Yj������H��Կ�|"�����%�ĩ���v.Dӿ��������6j���/��   �   ���1�ȾT){��\�
A}�@`[�]<T�<��< ��:v¼��f��7��be�|.�#PP�~7k�q'|�>�����z��h��K��(��Q ��7��^�C���r��23<�Z�<:� =4�< �ϻ�d�����}v���ƾ�����N�����4����ѿ����
�}�����8!��K��$�0�	�}w���ѿ�4��`;��Y~O��   �   &*��p��}��V'�DҜ�����`'�<�I="�=��<��R<�Y������z�BͲ�4��H^�n���1���� ��ؽ2�����[�P�Ҽ�$':؏�<X@ =<�>=4�/=�s�<0/������k �����侨�(�zNj�d��cR¿���(	�����(��b2��5��92���(�,}������v�¿�暿l�k��   �   ��:�b���;!���<������ż��<t�!=
>F=�@=H/=�м<�K�;p�b�x[�G�R�z��)��"l��q���V�l��2���Ѽ�ݹ��6p<�>	=�G=&o=8�t=�N=@�<�s�����0�4�����!A���9�����槿��ҿ ~����z(�* 8���B���F�޿B�8��(�F�����]}ӿ��������   �   �rE����pڭ��J�Sƽ\1�t�<"0=��b= �j=��T=b�)= W�<pQZ< �y��(]�����45���� W޼������`��;e�<�d=�&W=,��=	Y�=7�=N�_=��<\6��pѳ�I5B����� ��czC�깆�	{���2ݿ����.�0��-B���M�p�Q���M�F;B��1��U�V���;޿W�����   �   "I�"F
�<���tXO���˽���d<޲4=�k=��x=�g=F�B=�=���<X=<��
�0.1��?��,XSh�Ѕ�@hY;�<x��<��:=Ġp=v��=�ԕ=��=F9e=�f�<��{��E�F�-����G��G�G���k�����~�������3��E�B�Q���U�
�Q���E��&4�D���.�W������+���   �   �qE����|٭�ǀJ��ƽ�,���<J0=V�b=��j=��T=��)=�W�<�RZ< �y��']�(����4�ȭ���V޼���p��0��;he�<�d=�&W=S��==Y�=��=D�_= ��<�1���ϳ��3B�����s��vyC�P���Hz��2ݿ���� �f�0��,B���M�j�Q���M�^:B�&1�$U�����:޿����u����   �   �:�ˣ��j����<�Q�����ż�<��!=�?F=�@=L0=tҼ<�Q�;�b��Z��G���z��)���k��R���(�l�V2�`�Ѽ�۹��7p<?	=��G=�o=��t=r�N=Є�<Рs�N�����4�斟��>��*9�C��I姿оҿ|��܋�(��8��B���F��B�p	8�x(���g
���{ӿ����Y����   �   �*��l�P{���'��͜����,0�<�L=f�=��<�R<0U������z��̲����&^�O���1�t�� �rؽ�����[���Ҽ�E':<��<vA =��>=��/=�{�<0�.�����h ��|��d��7�(�FKj�b���O¿���t	�(����(� `2�v�5�T72���(�6{����	���¿�䚿4}k��   �   �����Ⱦ^#{��X��5}��A[�(]<���<���<�+�:�r¼*�f��6��e�@.��OP�R7k�O'|�0�����z��h�ݧK��(��Q ��7����C�h�r��73<_�<R� =�%�<�xϻ��c�����wv�o�ƾ�����N�3���1��F�ѿ���P
��z�D��6!�(I�F"��	�ws����ѿ�1���8��~zO��   �   ����ɍ��e�L�C�ݽHA=���� �<�|<��P��4*��W���z3��\l�]	���ժ��V��5�ʾ�ξ��ɾ���������6����e���+������L�߼� :X�y<�s<��F���)���ս_I�4U������S�/��Sj�r����D���Կ*	�������"����n���)�B@ӿ켴�p����0j�ž/��   �   �YȾ�J�����e���� �0U�� ����B���#�©�4��
�S� y��]ٸ�����v<�S������z�a��U �fNݾ�ɵ�]I��]?M�N,��a��� �Pfػ੘;@����缀흽�[������WȾ<��օ@�E�v��䖿-���/ȿsڿ�n�*�P��hWٿ�Iǿ�S���5����u�~�?�����   �   d���^�B�f�޽fW�P���KǻhbQ�*8��]��X����b�ՠ���վ�d�0!���8�*CK���V���Z�1uV�IJ�%p7����R��'�Ҿ��֜]���������@�!� ����dT��.߽N�C�S���K޾u��C��Kq��p�����1j���ǹ�Zۼ��e��ػ��y���♍��o��B����2ݾ�   �   �Y��� ��ج�9�8�"����� ������H�\�(��0�Gl�D�8�_f[��z�������
���>��.o��̜x�L�Y�i7�������#����Y�l�`��h���C��|"�����¹��d��o�\������㾆i��8�|b[��z�� ������N��i<���l��L�x�>�Y��7������6 ���   �   ��p��
��@�!�������riT�q3߽�C��U���O޾rw��C��Oq�s��u����l���ʹ�޼��h��x����������o�L�B����Yݾ|�����B�e߽�
W�l����Kǻ@UQ�01�&X��:��ߜb�WѠ�B�վ�a��!��8�?K�/�V�g�Z��pV��DJ�<l7���M�� �Ҿ����]��   �   Z����-ػ0Ș;� ����缈�m^��₾�ZȾ/��^�@�i�v�k斿F/��72ȿڿ{q��,�$ �!ZٿLǿ�U���7��j�u�P�?����7]ȾM���������r� �]�� �	� �B���#�g��������S�)u���Ը����
9�������)w��]�oR ��Hݾ�ĵ�HE���8M�9'��   �   d�߼�?: �y<ؔs< �F���)���ս�aI�1W������<�/�ZVj������F���Կ��!�H��($�^��ʼ�,Bӿ龴�%����3j��/�O���:�����L���ݽF=�����<Ќ<�����	#������3��Ul����Ъ��Q����ʾU�ξ�ɾ �������M2��"�e�R�+��{�����   �   H\3<�k�<T� =H)�<�{ϻ� d�.��bzv�@�ƾ�����N�N��3����ѿ����f
��{����b7!��J��#��	��u��f�ѿ|3��@:���|O����D�Ⱦ�&{��Z��:}��I[��)]<��<H�< $�:X]¼�f�.���_���-��HP��/k�|�����Czz���g���K�X	(�@L �S.��b�C� dr��   �   �G =��>=��/=D~�<�.�L����i ��}��ݫ�A�(��Lj��b��Q¿��>	�����(�Fa2���5��82�ο(�<|����<�V�¿暿 k�*�o羹|���'��Ϝ�D����/�<`N=�=�*�< �R<�-�:����z�%Ĳ����X����,���s���Pؽ������[��Ҽ �):l��<�   �   2o=��t=X�N=���<�s������4������?���9�0���姿��ҿ�|��j���(�J8���B���F���B�N
8�@(��������|ӿu��������:�Z���� ���<�&�����ż,��<��!=�AF=@=5=�޼<���;�`b�P�bG���z��"���d��2���ztl��	2�d�Ѽ ���xYp<�E	=,�G=�   �   RZ�=X	�=N�_=T��<�1���ϳ�?4B��������yC������z��a2ݿ���<���0�(-B�T�M���Q�d�M��:B��1��U���,;޿��������rE�q��-ڭ���J��ƽD/㼨�<|0=0�b=�j=��T=��)=�^�<dZ< �x��]�x����'����(I޼���� i�`�;o�<�h=d*W=���=�   �   t1�=+��=���=*8=�>�;�l[��W��׃� �Ծ'�W>\��}���p����ݿ��65���R�(��+� �(����D_�>��˱޿A��Z\���
^����Aپ=���f��5M��0@����<\M=.Ny==Ł=��u=r�W=X|0=�=(O�<� g<���;�H�;��v;��;��Y<T��<Z>=z�>=F�r=��=�-�=�   �   �ͣ=�6�=��=�?7=���;v�R�ޝ
�I󀾯�о��/XX�����q���pڿ�������2�%���(���%�|�����`��0ۿ�.���Տ��
Z����7�Ծ���L��k���7����<(�I=� r=�Vx=�f=N�C=V�=Ե�<Hk< ��; �$�P�ػ@d黠}�@�E; uU<��<t =��X=(�=Ȩ�=�   �   �X�=vڒ=���=v4=��<fh:�����`!q��Oľ�����L��ڇ������п�������m����S �z��`��	��$�)пi?��d}���jN�����Ǿ��y��	
�*�j�p�����<�?=`�[=�U=d�6=�=���<�1R;��:�X�ż�
�F"�Ҏ&�^`�Ď�X���@܂��E�<��=�(J=�n=�   �   ��]=��w=�j=~�,=0�G<��b�޽VW��&���"�7;�S$y�����7ڿ��,࿀���z�	�V����0��N�	�H�����t���;��B�y�G=<��]���<R^�Mf�Ї@� D0� P�<4Y+=T�4=�D=H��<`��; �d�x���g������䵽�|ǽ�˽�½�)���\���@@�(ļ Sչ\G�<�U&=�   �   ��<2�3=�B=��= �}<�)Ҽj��4F6��꘾�N辎�$��;\��G�������-ȿ%�� ���o����K�����c�>�ǿ(ͪ�/K����\�� %����.��v�;�S�ý���8�;4�<j�= @�< ��<�����P���}��A���i��r/�ܝ/���<���@���:�(C+�ܪ�^6� 9���'M��֘�0M<�   �   @@�x��<�	=��=<�<�xj��,��-��*�{��¾��
�]N;��p����/���:6ÿ��Կ5�߿��㿚�߿�@Կ�¿V,��7�����o��0;���6�¾�~�\��n������`<о<���<�j <�'^�r�:��?���*���1���^��?��vϜ�|㟾�ӛ�6����Y��u W��{(�)��ך��:N��   �   2w0�P��`us<h��<H�<�nz���5���ؽ�C����!d�����tE�ILs�ᑏ��̢��Ʊ��=��3a��Zﺿ">���(����!=r�ѨD��S���߾i���YD���ܽ�AB�p��hM<��<�S�;�T��tAV���ɽ�T�\��Ǝ����t�ʾ�,�,Hﾡ��l[Z߾�DȾ�C���劾N}S�T'�㶽�   �   ���8$5��9��/<<���<� �;�ż����C�h�����8~�X��|A��9e�҄��)Ɩ�0^���~��"m���ၿ��c���?��o�����-����f����x0��șʼ�.3;hLT<P��;h�i�ҕN���ν(�(�Hv�Z��D�Ҿcl������!��_+��.�h�*��� ��L�lj���Ͼw����o���!��   �   �
��m������ڞ��d4<�*<`�ڻԋ%�%����y#���z�WȰ�y��Zj�R/�[H��0\�Q�h���l�0?h��A[��G��-�N��V�������u���6h����������i4<H*<��ڻ
�%�Y��T~#���z�6̰�L��@m��
/��^H��4\���h��l�ZCh�wE[�� G�Q�-������l��J�u��   �   2�f�����4��أʼ�3;xOT<P��;P�i�h�N�a�ν$�(��Av�C��V�Ҿ�f����&�!��[+�A�.���*�� ��I��d��a�Ͼ�����o���!���R5� � =<<���<��;�ż7"����=�h�R������
���A�R=e�ᆂ�`���jȖ��`��逖�Jo���みL�c���?�&r�¥�1���   �   �k��]D�*�ܽZGB����pM<TÊ<�~�;D��l5V�Z�ɽoO�p\���b���6�ʾ�&�3Bﾔ��U�U߾�?Ⱦ
?���ኾ�vS�D"�;۶��k0��h�ȉs<��<��<��z��5���ؽĪC������g���dwE��Os�ϓ���΢��ȱ�@���c����Z@��+����J@r�u�D��U���߾�   �   ��¾C#~����<���\��H<�Ӿ<���< � <�^���:�H7���%�l�1�j�^�t;��꒾oʜ��ޟ�]ϛ������U��n�V��u(�7��ޒ���A�@�8��<�	=
�=l�<��j��/������{��¾w�
��P;��p�������Q8ÿ��Կ��߿ۣ��߿CԿ�¿.������H�o��2;�E��   �   ��龹����;���ý���P2�;T�<V�=�I�<<��<�c��D�n�}��8��2_��v)�\�/���<���@�3�:��<+�����+�0���M������r<���<�3=�!B=v�=��}<�0ҼGm���H6�t옾&Q�C�$��=\�OI��2���=/ȿ�����p���M������d���ǿ�Ϊ�ZL����\�
"%��   �   �^�^ ���S^�wh�,�@� 1�\Q�<B[+=��4=�I=���<��;��d������f�d��۵�~sǽp�˽}�½� ���T���1@���ü й�X�<�\&=��]=��w=��j=��,=X�G<V��J�޽�W�((���#��8;�+&y�����ۿ�>.�!���\�	�D�����&�	�͆���࿗��� <����y�v><��   �   7���Ǿ��y��

���j��������<8?=��[=f�U=Ϊ6=T=���<��R; �:�H�ż��
�V�!�&��T�<x꼠��������U�<��=�-J="s=dZ�=xے=��=V4=@�<&k:����#q�8Qľ؃�M�;ۇ�|����п���l 	�~n����dT ��z�ba�Z	��%��п@���}���kN��   �   ����ԾO������Qk���7�� �<��I="r=VXx=�f=6�C=қ=��<�Zk<pΚ; �$���ػp5�@�|�`�E;�U<�
�<N	 =�X=o�=Ω�=�Σ=[7�=!�=�?7=���;\�R���
���u�о��XX����Or��sqڿ����b��l���%��(��%������\a���ۿ)/��(֏�KZ��   �   ���پ���"���L�� >�d��<�M=xNy=cŁ= �u=��W=�|0==�O�<�g<0��;PJ�;��v;���;��Y<D��<N>=h�>=,�r=
��=�-�=`1�=��=���=�8=p:�;�m[�X�؃�^�ԾO��>\�~���p����ݿ���@5���V�(��+���(����:_�4����޿�@��C\���
^��   �   D��m�Ծ����t���i��x/���<�I=�"r=Yx=vf=��C=V�=��<0\k<њ;��$���ػ4�`�|�`�E;��U<�
�<p	 =�X=��=�=�Σ=�7�=��=�@7=��;r�R���
��Y�оZ��WX�\���q���pڿr�������
�ش%� �(�Z�%��^��L`���ۿc.���Տ�I
Z��   �   ���Ǿ��y��
���j��}�����<`?=@�[=� V=��6=H=T��<��R;0�:��ż�
���!�d�&�8T��w����@���4V�<̈=^.J=�s=�Z�=ܒ=ؖ�=�4=��<�e:�λ��% q�Oľc��(�L�ڇ�����п���F��8m�@�� S �dy�`�4	��#�5~п�>���|���iN��   �   �\�n���O^��b�*�@� t+�pY�<>^+=�4=�K=$��<(�;��d�v����f��򘽍۵�2sǽ,�˽D�½� ��tT���1@�$�ü �Ϲ�Y�<f]&=��]=r�w=�j=�,=��G<�����޽vW�:%���!�K6;��"y���ٿ�q+�������	�n�
��B��l�	�����%�(��9��j�y��;<��   �   ���<����;��ýL��ph�;�<��=,O�<غ�<�T��nB���}�8���^��4)�$�/���<���@��:��<+����+��/��dM�����v<P��<��3=B$B=~�=H�}<�Ҽ�f���C6��蘾VL��$��9\��F��A����+ȿO�� ����n�ԙ��J�����a῁�ǿ�˪��I����\��%��   �   h�¾�~�H������`����.<,޾<�ǹ<� <��]���:�]6��%��1��^�P;���钾Vʜ��ޟ�Nϛ������U��T�V��u(��񽏒���@������<�	=z=��<_j��(������}{�h¾�
�AL;� p�S��b���94ÿ��Կ��߿&��D�߿�>Կ��¿q*������ߦo�0.;����   �   �f���UD�d�ܽ$8B� ���;M<@Ί<���;�=���2V�I�ɽ�N��\�O�6����ʾ�&�Bﾀ��pU�U߾w?Ⱦ�>���ኾ�vS� "��ڶ�^j0�pa�ؕs< ��<T�<��y�D�5�H�ؽ8�C������`ྛ���qE�Is����wʢ�Jı�K;���^���캿�;���&����9r���D��Q���߾�   �   b�f����n*����ʼ �3;�lT<0�;�si�t�N�0�ν��(� Av���#�Ҿxf��ш��!��[+�9�.���*�� ��I��d��V�Ͼ�����o���!�����5����N<<���<�[�;L�ļ��a�g�h�����z��aA�6e�Ђ���뎿�Ö��[��X|���j���߁��c���?��l�T�쾎*���   �    ��`������n����4<�0*<ЉڻF�%�����dy#�>�z�"Ȱ�F��Aj�=/�[H��0\�D�h���l�*?h��A[��G��-�L��O�������u���hg��f�� ����4< 3*< nڻt�%�e���|u#���z��İ�ʦ龇g�	/�oWH��,\��h���l��:h�z=[�3G���-�f��w�������u��   �   B����5�(���_<<���< Q�;�ż���k���h�����~�?��fA��9e�Ȅ��!Ɩ�*^���~��!m���ၿ��c���?��o�����-��q�f�.��d/�� �ʼ��3;�kT<� �;x]i�XN���ν�(�;v�;��y�Ҿ�`�������!�7X+���.�!�*��� �KF�_��f�Ͼk����o���!��   �   �]0�=���s<���<� �< z��5��ؽu�C�ډ���cྰ��rtE�1Ls�֑���̢�~Ʊ��=��.a��Wﺿ >���(����!=r�ѨD��S���߾mi��zYD�Ǝܽ?B�����7M<|ъ<���;\/�� (V���ɽJ��	\�����������ʾJ!�4<�y��|O�aO߾;:ȾU:���݊�)pS���rҶ��   �    ��h��<(	=�= �<hj�!+�����ǀ{��¾��
�IN;��p����$���/6ÿ��Կ,�߿|�㿕�߿�@Կ�¿V,��7�����o��0;���)�¾�~���Q�������(<�߾<ι<P� <p�]��:��.��O �,�1�,z^�c7���咾�Ŝ�	ڟ��ʛ�e𐾨Q���V��o(��������3��   �   ���<&�3=�'B=(�=��}<#Ҽ�h���E6�q꘾qN�}�$��;\��G������u-ȿ�������o����K�����c�?�ǿ(ͪ�0K����\�� %����"��<�;���ýd�� Z�;`�<��=TW�<@ǃ<���7���}�U/��gT��k#�̐/���<���@�J�:�$6+���!콄&���M�(���X�<�   �   *�]=b�w=l�j=,�,=��G<�����޽W�j&���"�q7;�E$y�����-ڿ��,�v���t�	�R���.��N�	�I�����t���;��D�y�H=<��]���R^��e��@� P-��X�<l_+=��4=�O=(��<�g�;ؙd�P����f��꘽�ҵ��iǽ��˽ސ½��� L���"@��ü Mʹ�k�<�d&=�   �   �\�=Tݒ=���=�4=X�<�f:�	���+!q��Oľ����L��ڇ������п�������m����S �z��`��	��$�*пk?��e}���jN�����Ǿ��y��	
��j��������<�?=��[=\V=��6=D=̲�< <S;�|:��ż�
�^�!��v&��H�<a�u���|���f�<܏=>4J=Rx=�   �   �ϣ=V8�=��=pA7=p�;��R���
�<󀾤�о��*XX�����q���pڿ�������0�%�~�(���%�|�����`��3ۿ�.���Տ��
Z����5�Ծ���8���j�� 4���<(�I=�#r=0Zx=0 f=��C=0�=���<�lk<���; <$�p�ػ��S|��4F;��U<,�<� =��X=�=��=�   �   ┾=>�=!/�=��|=���<PҔ��(����8��c�����(�x�a�?���ݮ��̿ &翦
�����6����%"���[�Ϳ;T��_��B�b��=*��򾰔���$F�	�ҽB�@þ;\�=|@Q=�r=
y=��n=*�X=�W==Fx =z=t\�<h�<X��<W�<P�<�>=(w(=nQ= �}=��=�=���=�   �   �@�=�W�=��=��{=��<����j���V4�+��Xg�π%��]���������mɿ�m�}���(��X�������/���ɿ*e������:�^�'�FN���MA�C̽Ը� `�;:�=�qO=�#m=\�p=��b=�nI=�*=9	=@��<H��<8�{<pP\<�j<�t�<��<��=h�4=�d=�h�=��=6��=�   �   4�="�=���=�x=|q=��D�OК��T'��}����۾cw���Q�H������Oƿ�)�ؿ*������������h�ؿ�鿿�ڣ�|h���S����^߾�
���?3��P��<o��8%<8&=�uI=�]=Z�W=X4?=JP=8��<t̃<�y�;`.J��)�`�P�P\L��� �n��B <p�<2=��S=
�=�@�=�   �   �Q�=S��=*�=�Hq=f�=0T���5����\�����ƾRV���?���u�c^��Ƙ��X�ǿ��ٿ�C��0��#�5�ٿ��ǿ����9s��2&v��@��Q�٦ɾ�[���]������]��x�o<�C=��==��B=��+=\=d�<`;`�h��w򼠳/���X���o���r�~`�^9�' ���g�@�;lm�<�-=,m=�   �   �2J=��v=Lڀ=.	d=�=`�I;4�B��I��Y[��F�����Ⱥ(�[*Y�g������챿.2¿5�̿�п^̿^���)���㜿�J��-2Y��)�G����'���a�p��ttn���-��G�<$f=�4)=�=\p�<��<�DC��G�p�r��p����ѽRV��-��W�f�����������댽��.���05<��=�   �   �|�<��)= HQ=�`N=��=��=<�G��M���� 1�4i��aо1��\�8�0d�VɆ�����Q��^�� g���+����������l��(sc�fJ8��e�o�о�<��Hr4�e�Ž�� �:���<2F="#	=<.�<��n;xĳ�(TW�5���Χ��3���d=�+U�3�c��h��a�EdO�C�4��O��1ܽ叽��� x?��   �   ��.�(y�<j@=z .=��=�Ν<p`�{��M���Y_�N�����澁���C;�qw^��}��势�����*���c��<����|��]��Y:� ���m�ճ���~^�h_�Ӆ�(���xK<���<��<��< A8;8]Ӽ[����ؽ(Q��"P����J���ؿ��n���M嵾�^���[��d�����w��D���u�����B��   �   �*U�p�I���<��=>I=ܕ�<���:�l� 㸽6M$��|�B��">뾊Q�'0��{I��n]�Aj��Mn�X�i�@�\�oH��.���g��I���F:x��t �Ju����� �k:�/�<���<�H�<���;tt��������(1��0t�9	�������1ݾ�����\s�ʄ�J��Aھ�/��������i�&���ѽ�   �   ��ν�B� <���<���<���<�An<�%T��~\�x~ݽ�3�6������&ݾ����l�(���2�)6�^2���'����ɉ�"�پ+䪾�`|���+�"�ν��B�#���<���<���<�3n<�>T�.�\�E�ݽ�3�7��h����ݾ4�����(�[�2��6�da2���'����X����پ�窾�f|�$�+��   �   �x �wz����� �j:�+�<8��<N�<`��;�d��C��ݳ�1�0*t�^��v���~,ݾ������pp������<ھf+���~����i�6&���ѽpU���I�H�<ޱ=�I=x��<�&�: t�r踽Q$�T�|����bB�T�0�?I��r]��j��Qn��i���\�CrH���.�
�h��x���,?x��   �   т^�$b��օ������K<$��<���<��<�8;�JӼ
��f�ؽL��P�v���.���`��������ൾ�Y��8W��Z���b�w�ٖD���_���&�B�P�.����<�D=�".=��=0ʝ<�-`�r"��B���]_�������ĵ��F;��z^�W�}��犿�����,���e��
���[�|���]�9\:�9���p�j����   �   �>���t4��Ž����ŏ:8��<2G=�%	= 8�<`o;����fGW�C���*������|^=�$U���c�-h�w a�f]O���4��I�,(ܽݏ����@�>�ԋ�<��)=fKQ=bN=�=(�=<PR��k����#1�Tk���cо����8��d��ʆ�j���S���_��i��e-������A���n���uc�xL8��g���о�   �   �)��^
a� ���xn���-��E�<�f=�6)=��={�<�<HC��;��r�~h����ѽL�|(�vR�����b�㽐���a㌽��.�����\<`�=�8J=��v=~ۀ=�	d=6�=`�I;H�B��M��\[��H��������(�x,Y�Jh����M�3¿�̿�	п�_̿��������i䜿L��4Y�:)������   �   B�ɾ�\��_�����0b����o<D=�==l�B=R�+=�=�<`�;Мh�h`�n�/�B�X��o�~�r�|`��8�� ���g��c�;�~�<�-=�1m=�S�=���=�*�=�Hq=P�=�h���7����������ƾ~W�+�?�Ȼu�q_��������ǿ	�ٿ2E�92�C%忋�ٿ��ǿ����'t���'v�)�@��R��   �   �_߾d���@3��Q��,r���%<V&=�vI=��]=��W=�7?=�T=��<�ك<���;�I�H��P��5L��
���l��d <|��<�8=,�S=G�=�B�=��=�=��=�x=xp=�D�Қ�V'��~��D�۾Ex���Q����o���0ǿ�!�ؿ+�����+��������B�ؿ�꿿�ۣ�i���S�����   �   �N�Y��ZMA�~C̽`��@^�;b�=�rO=�$m=��p=��b=*qI=�*=f<	=���<���<(�{<@c\<�j<~�<���<��=�4=H�d=>j�=�=��=#A�=X�=��=N�{=8�<����9k���W4����,h�X�%���]�C�����nɿn����r�����\��c�����p�ɿue��٢����^�['��   �   �򾆔���$F���ҽ��@ƾ;��=�@Q=r=Ly=�n=z�X=,X==�x =hz=]�<��<���<\W�<��<?=8w(=nQ=�}=��=�=���=ϔ�=$�= /�=>�|=���<�Ӕ�U)����8��c����	�(���a�W���'ݮ���̿1&翳
�����8����"���[��Ϳ(T��K���b��=*��   �   vM�v��LA��A̽ȶ�Pm�;��=�sO=�%m=~�p=z�b=�qI=H*=�<	=���<t��<��{<xd\<� j<x~�<��<��=*�4=z�d=Uj�=�=1��=NA�=EX�=$�=`�{=X�<ે��i��{V4�����f龈�%���]����J���&mɿm��������Ι�W����㿖�ɿ�d��9�����^��'��   �   �]߾�	��>3�tN��Xh�� "%<)=�xI=r�]=j�W=&9?=V=|��<�ۃ<@��;��I�����P��3L�P�
��sl��e <���<�8=��S=|�=�B�=��=x�=���=ցx=�s=H�D��Κ��S'��|����۾�v���Q��������ſ�N�ؿ)����
��������q�ؿ鿿ڣ��g���S�(���   �   �ɾZZ���[�����xT�� �o<�G= �==�B=��+=�=���<��;��h��]�J�/�H�X��o�ʖr��`���8�r �Ȧg�@g�;��<��-=D2m=lT�=f��=�+�=�Kq=��=�6��\3��n�L���\�ƾ\U�n�?�l�u�s]������ �ǿH�ٿNB�L/�a"�͉ٿ6ǿ`���,r��e$v�r�@��P��   �   �%���a� ��jmn��-��Q�<Lk=�:)=��=p��<��<�C��9�<�r��g��ߠѽ�K�B(�ER�U�����O���$㌽�.����(_<4�=�9J=<�v=�܀=hd=T�=�%J;V�B��E�LW[��D������>�(�o(Y��e��a��A뱿�0¿��̿3пU\̿���������᜿�I��0Y��)������   �   ~:���n4�f�ŽV����:���<VL=*	=�>�<�1o;����EW�#�)���$��^=��#U���c�� h�J a�A]O�ة4��I��'ܽ�܏�����>�4��<��)= NQ=�eN=��= �=<|:��⪺��1�5g��f^о{��>�8��d��ǆ����O��2\��5e���)��M���񨘿k��vpc�H8�d���о�   �   �z^�\� ΅����� 'K<��<,��<4!�< �8;�DӼ���-�ؽrK�0P�;�������8�������nൾ�Y��%W��I���B�w���D�l����L�B���.� ��<NG=d&.=P�=۝<X�_����;���U_�����|��V��:A;�mt^���}� 䊿�����(��b��`�����|��|]��V:�����i�찥��   �   �p ��n����� �m:�=�<���<DX�<0�;�]�������轁1��)t���>���M,ݾh�����bp������<ھX+���~��`�i�&���ѽbU���I�@�<��=^O=���<@��:�c��ܸ�@I$���|�����9�
O�B0��xI�jk]��j�(Jn���i���\��kH��.����˕���4x��   �   y�νưB�X���,�<���<x��<�Tn<T��{\�*}ݽL�3����^����ݾp���Y�(���2�6�^2�y�'����ĉ��پ䪾�`|���+���ν.�B� ��#�<���<���<�^n<�T�Ts\�'wݽ&�3�1��⟮��	ݾ�
���7�(���2��6��Z2�D�'��������پMા�Z|���+��   �   U�جI�l"�<0�=�P= ��< 5�:xi��ḽ�L$���|����=�lQ�0��{I��n]�0j��Mn�L�i�9�\�oH��.���]��=���&:x��t ��t����� �l:|8�<���<�[�< 5�;,P���������
1��#t�{����i'ݾ������zm��O��t7ھ�&���z����i��&�`�ѽ�   �   ��.�Ę�<BL=6).=
�=X؝<`������9Y_�������d���C;�Xw^�˃}��势�����*���c��9����|��]��Y:����m�ɳ���~^�,_�U҅�d���8K<��<��<`'�< 59;d4Ӽ����ؽ�F�PP�ê�����ܶ�������۵�U���R��-�����w�c�D�(�y���ԕB��   �   p��<�*=�QQ=�gN=��=��=<$B��)���y 1��h���`о��D�8�d�KɆ�����Q��
^��g���+����������l��$sc�dJ8��e�i�о�<��r4�΍Ž8���w�:���<�L=6,	=�F�< �o;���H9W��밽�������W=�U���c���g��`�WVO�t�4�"D�	ܽ�ԏ�����>��   �   �?J=��v=ހ=�d=D�=@J;��B��H�Y[��F��������(�E*Y�g������챿#2¿-�̿�п^̿[���)���㜿�J��+2Y��)�B����'���a�:��sn���-�hN�<$k=�;)=��=���<��< �B��.�čr��_��ۗѽ�A�#��L��y��ߌ��켽�ڌ�@�.��ꁼ0�<p�=�   �   �V�= ��=�,�=�Lq=h�=B���4����8�����ƾCV���?��u�Z^������P�ǿ��ٿ�C忼0��#�2�ٿ��ǿ����:s��2&v��@��Q�Ӧɾ�[��~]�W����Z��0�o<zG=ؠ==�B=�,="=��<�,;Pqh��G�/��{X���o�؇r� `�\�8�& ��vg����;|��<�-=8m=�   �   Z�=��=p��=��x=xs=؆D��Ϛ�nT'�x}����۾Ww���Q�B������Hƿ�"�ؿ�)������������f�ؿ�鿿�ڣ�|h���S����^߾�
���?3�cP��lm��X%<�(=<yI=��]=X�W=�;?=�Y=��<P�<@��;@I�8��x�P�hL��
� 5j�@� <D�<�?=H�S=��=�D�=�   �   B�=�X�=��=��{=��<T����i���V4���Kg�Ȁ%���]��������~mɿ�m�z���&��V�������-���ɿ+e������<�^�'�GN����LA��B̽f���e�;P�=�sO=&m=L�p=��b=|sI=p*=�?	=��<���<��{<�u\<�2j<P��<���<��=��4=��d=�k�=J�=&��=�   �   ���=9�=@�=p,�=~7T= �e<� �	�佦?T�h���P��J&�V�����?��`��yZ����ʿcο��ʿHi���+���{�����W�k'�� ��S߭���c��v���l���8U<Z~=�J4=X�H=�|L=(�E=�;9=""+=��=�V=��=��=r2=��=�1=2�K=�-l=Њ�=.��=�߮=O��=���=�   �   �P�=K��=`B�=���=\�U=vx<FR�6#޽�PO��褾֓ﾍ#�yIR�rf��ϡ�����.���tǿW�ʿMuǿ$7���6��RԘ������&S�ZF$��9�$0��r.^�v:������ň��Ih<��=g4=0�F=�G=�>=(�.=�k=J�=X��<,�<�{�<`�<�=��=h91=NvS=��z=��=7T�=^n�=�;�=�   �   ��= ��=�=ۺ�=�Z=Ĥ�<� �v�ʽ2A��Ú�I�ᾟ��5G���u����v���W����������
����볿����Q����u���G��%�| 從��j�N�D(𽠹a��o;��R�<�w=�*4=DZ?= �8=t�&=9=Ȅ�<�۱<@e�<�?<�{<8U<x}7<���<@��<��=��5=vtg=�[�=�Ԣ=(�=�   �   �v�=���=,��=��=h._=���<�������f�*�^����e̾.�e�5���`�����7���w������آ���w��~Z����������`�=6�o����ξ�Վ��@6��Vͽ��0� �]����<�7=�1=�B1=�=���<Dv�<�@&< � �&�hܔ�X���\RԼh^ɼ�W����.���:p^~<���<�?=��{=�_�=�   �   �׈=��=�Н=�R�=�#c=�#�<�3�󫇽R��
;n�PU�������7SF�Sik���P钿��؝�~���~����ᅿ6k�� F��������液�nts��d��,��`����;���<Q =r�*=��=h��<Ȇ{< 88�Ո�h9	��I�ad��E����q���i�����7{��;��_ܼP�Ļ��z<HM=��Y=�   �   ��:=Fu=i+�=��=�bc=N�=�R�:��<��z߽$�A�U���i;����G(��H��e�Hu{��ڄ��A��������z�Rvd�N�G��'�e�Z�̾t��S�C�c,���^�X=:��<�<p�
=2�$=
Z=,E�<�M]< �Ȼx���\�`5��Кӽa�������Z�L����(����$l��
Wf�=޼��*:(�<�   �   T|�<�r$=�J\=:`p=҅]=�B = `R<�Լ�8��X���h�\����Aھ�	��$�w<���N���Z�:�^�ҝZ��PN�i7;�#������׾�r����d����0٠�@��p|�;��<�="=:I=l��<�	ڻX��.��4�ҽ3����2� �R��\k��z�L�~���v�׿c��3G�ӣ#�|%��#��,W3��� ��   �    �h��փ<��=�H=�O=��,=�z�<p��ּH���ҽ8�,��z�񎨾�zվ
� �n���=#���,��,0�Ҍ,��m"���������Ѿu����r���$�}�Ľ��4����t�<8h=�C,=�G=j�<@����M�|m�����>)��>]�k͇�;+��Z�����������E��&ˬ��ř�������N�Q���ɽXX��   �   |�W���G�a�<�;=��8==1=ܳ�<P�<0꼼4���:�~�3�v�v��B��e��P/޾f����t���J�����ھ�ʻ�e��Kk��'���ӽ0�W�`�G��k�<�>=x�8=�<1=���<@�<�����8��kA���3��v�F��e���3޾Q���:w�����������ھ�λ�����k�6'���ӽ�   �   *Žޡ4��N����<2f=�C,=hI=�p�<@K���E��g��,�:)�9]�ʇ�j'��0���$���O��(A��Ǭ���������N����u�ɽ*LX��h��<�=��H=гO=��,=Du�<`黪�H�`�ҽ�,��z�!����~վM� ����|@#���,��/0���,��p"�C����S�Ѿ����Ͳr���$��   �   ����ݠ���＀[�;�<B�=�"=�K=訁< �ٻ\��0����ҽ�����2���R�Vk��~z�~~���v�!�c��-G�`�#� ��@��|J3�� ����<x$=FN\=*bp="�]=�A =hRR< Լ=��l���h�����Dھ�		�H$�%<���N���Z�I�^�͠Z��SN� :;�N#�����׾hu���d��   �   @�C��0���^�(N:��7�<>�
=N�$=�[=dK�< a]<�bȻ����\�9.��g�ӽۘ�����GU������"���Ὅc��BHf�0$޼ ]-:$�<ب:=�u=�,�=<�=�bc=��=�ݒ:��<�R߽N�A�x���l;����I(�t�H�~e�&x{�g܄�:C��u�����z��xd���G��'��f���̾k���   �   ws�vf�f/����P�;��<�P =X�*=�=���<P�{< ���È��.	�|�I�D]�������i��ra����f'{���;��EܼpzĻ��z<U=,�Y=ڈ=^�=�ѝ=S�=T#c=��<��3�߮��x��>n�XW��������(UF��kk�I���꒿m��nٝ�����û���ⅿCk�R"F�S����������   �   �֎�fB6��Xͽ��0��^�x��<`7=��1=JD1=|�=8��< ��<HY&< ?���&�\Ȕ�����H;Լ�Fɼ�@��@�.��9�:X�~<���<��?="�{=�a�=fx�=Ά�=䶬=��=�-_=���<T���6��K�*�����Vg̾7/���5�y�`��	���8���x�����������x���[��� �����&�`�T>6�e��8�ξ�   �   \���|�N��)�лa��u;��P�<0w=+4= [?=��8=��&=D<=،�<��<�p�<ȫ?<��<�r<p�7<��<|��<.�=|�5=�yg=�]�=i֢=��=��=��=Z��=꺛=$Z=���<R  ��ʽ�A�Ś����|��6G�̔u�P��:���'���~½����׹���쳿=��������u���G�/&�}��   �   w0���.^��:�q���8ǈ�@Hh<��=Dg4=��F=ܼG=&>=г.=�m=��=<��<� �<���<��<f=��=�<1=�yS=��z=+�=NU�=?o�==<�=$Q�=���=�B�=u��=��U=�qx<T��$޽pQO�3餾���#�JR��f��3���}��7/��Huǿ��ʿ�uǿ�7���6���Ԙ�ͳ��0'S��F$�e:��   �   -߭�j�c���;���Ŀ���U<�~=�J4=��H=�|L=j�E=<9=r"+=H�=DW=
�=��=�2=8�=1=^�K=�-l=֊�=(��=�߮=N��=���=��=(�=,�=M,�=$7T=��e<ʰ �����?T�Bh��9Q��k&�5V������?��o���Z����ʿcο��ʿCi��}+��|{�����hW��j'�� ���   �   �/���-^��9�󏀽���Oh<�=�h4=ԦF=��G=">=´.=�n=��=���<�!�<��<��<�=��= =1=�yS=ʚz=B�=hU�=Zo�=^<�=LQ�=���=�B�=ꝝ=�U=Pyx<XQ��"޽PO�D褾i��B#�IR�8f���������g.��mtǿ��ʿ�tǿ�6��6���Ә�7���5&S��E$�(9��   �   �~��ۓN��%��a�pd;��W�<z=�-4=R]?=��8=��&=>=(��<��<Hs�<x�?<��<v<P�7<���<t��<��=��5=zg=^�=�֢=��= �=H��=���=Ȼ�=�Z=ਖ<$ ���ʽA�8Ú�A�����4G���u���ȗ��������(��5���볿ϛ�������u���G��$����   �   KԎ��>6�vSͽ��0���]���<b;=��1=nG1=b�=���<��<xb&< 0�X�&�(Ŕ�Њ��9ԼEɼ ?��؟.��K�:��~<���<x�?=��{=6b�=�x�=k��=���=4�=*1_=��<ܨ��
����*�7���
d̾-�+�5�X�`�����6���v��x��������v��cY������ ���`��;6�J����ξ�   �   6qs�b��(���}��A�;���<�U =��*=ʢ=t��<�{< �� ���>,	�H�I�P\������i���`��n񓽢&{��;�`Dܼ vĻ��z<�U=�Y=�ڈ=�=�ҝ=�T�=�'c=�+�< |3�����.��/8n�mS��������hQF�8gk����	蒿����֝����,���Z����k��F�8�����ʹ���   �   ��C�,'���^��#:��G�<��
=��$=:`=�S�<Pp]<`FȻT��ܛ\��,��6�ӽЗ��L���T�f�Փ��"����=c���Gf��"޼��-:��<�:=0	u=�-�=��=Vgc=(=��:<�<�	v߽��A�?��g;W���E(���H�;e�wr{�nل�6@��~�����z��sd���G� �'�Mc�}�̾6���   �   <���Ӡ����p��;�!�<��=R"=`P=l��<��ٻ�������ҽ�����2�m�R��Uk��~z��}~�?�v��c��-G�6�#��������I3��� ����<�y$=�P\=bep=Ί]=^H =yR<�Լ�3����X
h�����(>ھ�	��$��<���N���Z�%�^�ĚZ��MN��4;��#����J�׾�o��t�d��   �   ��ĽN�4��ޝ��<fn=J,=�N=�y�<@Ȯ��A�f����H9)�d8]��ɇ�$'����������'��A���Ƭ�����o󁾤�N�n�� �ɽZKX���h���<2�=��H=X�O=F-=܇�<��ʲH�F�ҽ�,���z������vվʊ �����:#���,��)0��,�0k"�;������Ѿ#�����r���$��   �   
�W� [G�0{�<tE=��8=C1=ܽ�<X�<�⼼Q2��9�3���v�\B����/޾/����t� ��:����~�ھ�ʻ�T��*k��'�T�ӽ@�W�|G�|o�<�A=��8=�B1=���<�<,׼�.��3�3���v�*?��S���*޾l���r�j���������ھ�ƻ����Zk��'���ӽ�   �    �h�<��<.�=،H=ƹO=-=ȃ�<��p�H�,�ҽ��,�[�z�����czվ� �P���=#���,��,0�Č,��m"���������Ѿf���Эr���$��Ľv�4����P�<�k=HI,=�O=(�< 3���:�a�����4)�3]��Ƈ�|#������������<���¬�꽙������N�{��ɽ�>X��   �   ԝ�<�$=�T\=�gp=��]=�G =PoR< ԼY7������h����@Aھ�	��$�\<���N���Z�*�^�ÝZ��PN�b7;��#������׾�r��ϋd�����ؠ���＠��;��<��=�"=&R=���<��ٻ������ҽ�����2���R�Ok��wz��v~�0�v�+�c�f'G���#�"������<3�xa ��   �   l�:=u=�/�=��=�gc=4 =���:��<��y߽��A����i;����G(���H��e�3u{��ڄ��A��������z�Lvd�H�G��'�e�Q�̾i��4�C�,���^�7:��A�<�
=R�$=Ha=�X�<�]<�Ȼ̧�*�\�<&��H�ӽ����J���O���b��W���ὄZ��l8f�$	޼ 30:�*�<�   �   ݈=��=�ӝ=2U�=�'c=�)�<��3�窇�����:n�U����� �� SF�=ik���H钿��؝�x���z����ᅿ1k�� F��������߶��Xts�fd�;,���漰)�; ��<U =�*=��=\��<�{<  �<���n"	���I��U��N���#a���X��R铽{�`�;�,*ܼ�ĻP�z<�]=~�Y=�   �   �z�=���=���=��=.1_=��< �������*�3���le̾�-�Q�5���`�����7���w������Ѣ���w��{Z����������`�=6�m����ξ�Վ��@6�SVͽ��0���]�Ė�<�:=�1=bH1=L�=x��<D��<Hx&< �� �&�����Dv��(#Լt.ɼh(��0t.����:��~< ��<h�?=��{=�d�=�   �   +�=1��=���=��=�Z=���<t ���ʽ�A��Ú�0�ᾑ��5G���u����o���O��������������볿����P����u���G��%�y 徙��\�N�(� �a��l;�8U�<^y=j-4=�]?=��8=h�&=�@=Ė�<��<<}�<P�?<�<P�<X�7<��<$��<�=��5=Dg=\`�=�آ=b�=�   �   �Q�=N �=&C�=��=B�U=�xx<�Q��"޽ePO��褾ɓﾆ#�pIR�nf��ɡ�����.���tǿW�ʿLuǿ#7���6��QԘ������&S�YF$��9�#0��m.^�i:�����4ň�8Lh<��=dh4=�F=V�G=�>=е.=p=p�=��<'�<ȉ�<��<=N�=f@1=�|S=��z=��=�V�=Np�=#=�=�   �   |]�=���=���=$ƹ=�3�=�+=@��: cZ����@[�Մ���|���<���_���N���I��	���L��Y�����QL`���<�� ��|6���fl�H�������K(�x�.���<�q�<1�<���<M�<���<��<�;�<�k�<���<Z)=�Q=�"-=}E=�\a=uN�=�H�=��=Ԟ�=
�=�8�=��=�   �   ���=���=:>�=(�=ȁ�=8�-= (;x3Q�	���<AV�=�����|1���8��[��-{�lቿ(����p�������牿BV{�^C\�cG9��8�i�ǐ����f�����é�������`	#<���<Hf�<`��<�i�<���<d��<�<���<���<Ĳ�<�=��=&b1=�M=��l=X�=�m�=~��=�t�=��=0	�=�   �   0�=�=�0�=�϶=�)�=|�5=P�;l�6�2��Z�G��,����Ծ���Խ.��\P�/n�ӂ��R��b䌿�L���͂�G6n�,�P��'/�0��+�׾������V���y���n�� �u�Uc<@��<��<<��<�I�<t��<�.�<��<��<��<PX�<�~�<[�<��<T!=̄0=.�V=�O�={��=�U�=츼=�D�=�   �   ��=���=6W�=�r�=���=�2A=��J<�,���Ľ�1��ш����c_��`;��D>�4�Y�.�o��c}�6���G}��Zo�y�Y��1>�YW�Q>����¾�{��$�=���Z�v� `��pn�;J�< ��<X��<�w�<t��<��<��I<���; c;�����)i�@�}��D��
;x�<tV�<�k�<f�&=b�[=:�=J��=��=�   �   ���=&6�=[�=GK�=٠�=tM=U�<p����K��8���+k��?���޾���G'�^�?��PS�
�_���c�(�_�Z�R��?���&�%A���ݾ�է�6#o�������l�.�@Y	�Ѐg<�>�<&4=�!=���<X�<�,(< .9�$�$��m��,����t�!��:�H����3����ڻx5<��<��,=�7m=�c�=�   �   �τ=��=��=���=퉎=��W=���<���(lh�����@���	��	뾖a���"��[3��>��A���=�A�2���!�`~��+龪7�������?�$���B��\��� ��;�{�<`�=de=�=���<(O< r޺,͏���ZN�<���w������̺�+��� ����ݑ�Z6_�F��hBK��g"<̓�<��K=�   �   ��1=p�q=QX�=4ӑ=�W�=j�]=,= �Y;��\3��Lm�LC\��%��pŽ�{E�H>��"�����������O��	�5-�!��F4���T����:U���� �� �<��=��*=t0$==�x�< ��:�C���$,�����|���x�뽵�
��Z�&;#�0$����nx����j�y�� ��7>����<�   �   ��<�!=R{^=�&}=z�|=L�\=f�=�m<`ӏ�Hm���ٽT�%�hd��`���ѱ�3�;��p��.A�����h�5!ʾ6����z����V����l���=�@��xY�<Ĺ=h==�C=��*=��<b-<��Z�B�+�ڗ��߽Q��5�6���U��am�e�{��D�v��c�v�F��V#�k����z��\x5�G/��   �   �0M�p��<��=�M=��`=>T={(=�4�<@$�������d��`%���V�vI��s���=����������ڱ�橥��4��k\x�3E���v\���1J�0M���<�=J�M=��`=�T=fz(=0�< ��l��0������N%���V�TL�������@��Ӧ��Z���dޱ�v����7��/bx�8E�,��c��<J��   �   l=� ��PO�<*�=�e==�C=��*=���<Xn-<��Z��+�x՗�~߽H��k�6���U��[m��{�����v��c���F� R#������s���l5�@"/�4�<J�!=D^=�)}=��|=n�\=�=�
m<dݏ��"m��ٽ۩%��d�uc��ձ���;!�㾱��}E��*���l��$ʾp����}���V�X��)���   �   �Y����@X�Xݳ<�=��*=�/$=�=�|�< �:�8���,�������ϩ�P�
��U�6#��*$����~s����қ��j�y�������=�0ʷ<��1=�q=�Y�=8ԑ=DX�=�]=8*=�fY;ԫ��7��2p�(G\�f(��lȽ� I�C@��$����D��ב��Q����0��#���6����T�����   �   ���\F�������l�;�u�<|�=ld=�=l��<�O<��ݺH������PN�P󅽪���]��
ĺ����뮪�֑�(_�r���K���"<���<��K=҄=��=��=r��=��=��W=���<��:rh�Y���@� �q���\c���"��]3��>�(�A���=�\�2���!����.�:��������?��   �   ��@���0�.��g	��ug<�:�<�2=�!=���<��<8(< t29��#�����p[漠"�Fy���!�4.��z��8���kڻ�\<@��<^�,=�=m= f�=y��=�7�=L�=�K�=ޠ�=�rM=dP�<H����N��T���.k�lA��9޾]��bI'�;�?��RS��_���c�1�_�H�R���?�&�&�xB���ݾ�ק��%o��   �   ի=�t��>�v�,f���[�;�F�<���<`��<x�<p��<��<@�I<0��;��;@︺�h�@N}���`:;(�<,g�<x{�<t�&=��[=�	�=���=t�=n��=���=�W�=s�=b��=�1A=�J<�0�F�Ľ�1�$ӈ�ĳ��sa���<�F>���Y�߈o��e}���8I}�p\o��Y�3>�qX� @���¾�|���   �   ��V����ѳ������v��Oc<h��<���<8��<�J�<̢�<�2�<`��<t�<��<�a�<@��<,f�<h��<�&=:�0=F�V=#R�=���=JW�=`��=
F�=�=��=1�=�϶=�)�=��5=0��;D�6�G����G��-��#�Ծ���ľ.��]P�=0n��ӂ�/S��匿rM��6΂�R7n��P��(/����(�׾m����   �   .�f�*��)ĩ����X��`#<���<�e�<d��<8j�<��<���<�<D��<P��<ķ�<ƃ=��=e1=� M=��l=��=�n�=��=�u�=���=�	�=^��=��=h>�=�=���=��-=@(;N5Q�Y���#BV��������1���8���[�=.{��ቿ����3q�����<艿�V{��C\��G9��8��i�!����   �   �fl�(�������K(�@�.���<�q�<$1�<���<pM�<��<���<h<�<�l�<���<�)=R=#-=Z}E=.]a=�N�=I�=��=۞�=�=�8�=��=x]�=���=��=ƹ=�3�="+= ��:�cZ�����c@[�����|���0<���_����$N���I��	���L��Y�����@L`���<�w ���]6���   �   ��f����©�"������#<���<�h�<p��<0m�<���<8��<��<���<P��<x��<v�=V�=�e1=!M=��l=��=�n�=���=�u�=���=�	�=���=H��=�>�=��="��=��-=@)(;b2Q�N����@V����V��61���8���[�-{�#ቿټ���p��d����牿�U{��B\��F9�:8�Wh�2����   �   2�V���������� �u�H^c<��<��<��<xP�<,��<�7�<��<� �<���<�d�<���<th�<L��<�'=��0=��V=_R�=���=�W�=���=JF�=\�= �=�1�=�ж=�*�=V�5=��;��6�c��(�G��+����ԾK���.��[P�.n��҂��Q���㌿2L��͂�!5n� �P��&/�g����׾�����   �   �=����h�v�$X�� ��;�P�<���<��<<��<\��< �<��I<���;��; ���`�h�`/}�`���N;x�<�h�<�|�<�&=(�[=7
�=���=��=���=?��=�X�=�s�=Ă�=�5A=0�J<�(��Ľ:�1��Ј������]��?:�SC>���Y���o�+b}�T���E}�$Yo��Y�f0>�V�:<���¾<z���   �   ���`�����.��E	���g<�F�<z8=�&=���<(&�<HJ(< �69��#�@����T����v���!��,�Px�����dڻ�_<���<�,=�>m=�f�=���=08�=,�=�L�=���=�wM=�]�<�w��xH����)k��=���޾���F'���?�OS���_���c��_�W�R��}?���&��?��ݾ�ӧ� o��   �   �}��>��D������;`��<<�=�j=��=<��<`!O< Nݺ䷏�z���LN���*������º� ��8����Ց�'_�����K� �"<��<��K=�҄=r�=��=���=���=�W=0��<���8dh����`�@��j����_���"��Y3�j	>���A�Y�=��2���!��|��(�
5������H�?��   �   �O�������캴�<�=��*=46$=�"=��< ��:|.�� ,�U����|���뽉�
�U�x5#�n*$�(��4s�~��d�����y�������=��˷<�1=^�q=�Z�=�Ց=%Z�=d�]=�1= Z;����-���i�?\�_#��Y½��A�G<�X �s�����N��aM����)�����1����T�h���   �   H
=�H���f�<��=�m==�#C=��*=$��< �-<�kZ���+�$ӗ�N߽J����6���U�/[m���{����v���c���F��Q#�����&s��
l5��/�<�<��!=$�^=,}=��|=��\=T�= 3m<0��m��ٽ@�%�p�c��]��dα�d�;�����<������d�`ʾ���w����V��������   �    �L�P�<��=
�M=4�`=�T=؀(=4?�<@��J��`���<��^ %���V�I������<��Ϣ��R���vڱ�ĩ��n4��9\x��2E����"\���0J�xM�@�<��=��M=�`=�T=�(=xB�<@���t��������$���V�aF�����L9��#��������ֱ�,���1��MVx��-E����#U���%J��   �   D�<T�!=P�^=�.}=.�|=�\=��= *m<Xʏ��m���ٽ_�%�� d�I`��lѱ���;���8���@��˚��h�!ʾ!����z��h�V�������=���H\�<ʻ=�j=="C=��*=��<��-<[Z���+��Η�u ߽����6���U�jUm�V�{���3�v��c��F��L#������k�� `5�X�.��   �   h�1=(�q=�\�=�֑=�Z�=p�]=�0= �Y;B���1��ll�~B\��%��Ž�-E�$>�i"�����������O��	�!-�!��44��ɋT�����T��4�����p�<4�= �*=b5$=�"=0��<�&�:�$��<,�����+w����j�
�xP��0#�N%$���Jn�a��+���<�y�����`�<�ܷ<�   �   2Մ=`�=:�=���=X��=��W=L��<X��
ih�w���@��񊾞	����ta�s�"��[3��>�ҡA���=�6�2���!�X~��+龝7�������?����B��t���p��;l�<4�=di=��=���<H)O<��ܺЭ����DN�,셽౟�	 ��a���=w��L����͑��_�����J�з"<D��<l�K=�   �   ���=�9�=8�=�M�=Ģ�=TwM=�Z�<(}���J�����_+k�C?���޾Ж��G'�G�?��PS���_���c��_�R�R��?���&�A���ݾ�է�"#o����߭����.�HU	���g< C�<67=:&=8��<h(�< S(< 0:9p�#��蠼hE漬��l�j�!�� ��`��L���ڻ��<���<x-=�Dm=i�=�   �   D��=\��=RY�=pt�=ꂒ=5A=0�J<+���Ľ��1��ш����2_��I;��D>�#�Y��o��c}�0��xG}��Zo�r�Y��1>�UW�H>����¾�{���=������v��^���v�;M�<���<|��<��<d��<��<p�I<���;@);@�@-h���|��&���;h�<�x�<��<�&=d�[=��=��=��=�   �   L�=� �=2�=�ж=�*�=�5=��;�6�����G��,����Ծ���ǽ.��\P�/n�ӂ��R��^䌿�L���͂�D6n�)�P��'/�-��%�׾������V���R��� ����u��Xc<�<���<���<�P�<h��<:�<���<�%�<��<xl�<���<�q�<<��<�,=܏0=��V=�T�=���=4Y�=��=~G�=�   �   ���=���=�>�=��=8��=�-= '(;�2Q�����AV�.�����v1��8� �[��-{�hቿ%����p�������牿AV{�]C\�aG9��8�i�Ð����f����ré�t������
#<콨<,h�<��<m�<0��<���<��<X��<��<���<R�=^�=�g1=d#M=8�l=��=�o�=���=�v�=t��=|
�=�   �   ܹ�=��=���=y�=��=cǃ=�_=P�ȻF_l�8�����L��e���aǾS����,�6H/�,�A�GM��QQ��LM���A�7~/�E���w��R�ʾG��D@_��
��Ž�|o��q�`���`j@���$��]7��W���j�pba��\2� M�����:��%<L��<�z�<�Y$=�6N=Jxw=F��=��=�;�=@q�=@��=���=L��=�   �   |��=xP�=��=�%�=@��=,J�=U=���n�c��j�"�G��N��(lþǵ���O�
	,�,>���I���M��I�>>��2,�j��Ro���ƾ�喾��Y���������d����P����G#�h
�0��PC�X@\��~Y��L2���˻ ־9��	<�2�<@4�<z�=��@=�gi=��=�՜='�=���=^��=ب�=�$�=�   �   �=���=</�=n1�=���=���=�y=@L�� ^J�&�ཌ�:�h������I��f�ў"�O�3���>�oB���>���3�B�"��7�z�꾰������4dJ����ܫ���E��#ʼ�4����@�v�PF�����0�4��E�h*6�H��`XU��BH;8�+<�M�<|��<��=HR>=g=�H�=~Ҝ=Ly�=�c�=ت�=S�=�   �   `V�=4�=ط�=V��=R]�=�І=0�!=�ٖ;zh$�v�ýw\&��mu��[����Ӿ3# �4��0�#���-��"1�}�-��o#���������Ծ���N�{��,2�cF뽀����|���n���� �H; 6X; � :�jn������0�(0I��D��w%��Dܻ�{��F|;�(2<��<$��<�$=��I=�!x=��=���=H��=��=�   �   ��=:R�=m�=��=Q�=e!�=.=E6<tp�r���N��lS�W��R���t�߾Dx��X��8��1����N���� ��W޾]B������J�T�*i�C����$N�L^���C޺H<�;S<حB<�a�;�:�:б��X�,���|�����pD�����@֭���� g�`M�����:�-A<��<��=,�P=�u�=�=pְ=�   �   
�=z�=���=$߱=6��=c�=��7=�Ώ<�'��~w�yD佴4.�B&p�a���Ż� �پ�)� ����@?��Gcﾌ
׾r���ܖ��hi�E*)�.ώ����P��c`�H�S<��<���<�۫< }s<�|�;�D9���L��7���5��nX��5���F���M�(H�B�4�x&��ȼH�&���;���<t;$=*�d=<�=�   �   t��=9��=���=懡=��=\��=D.<=�s�< rٻ�/�ܮ�- 	�;Y?�΄w�K���K��g¾�oξjҾ*�̾2���������P�j��~1��Y���`���_���˻�u<���<�q=j�=`�<�H�<��<@yg�t뒼~���D���~��㙽�D��s��V�½";����w���(�^�j����I�Pu<��<v�E=�   �   \�,=@�g=�#�=���=,�=��o=�8=��<`�;$��k}�ν8��%�=�Fhh����H��������#��Ռ��W��Ύ����W���)����gS��t!�x���<��=�i0=j>=l�4= �=�b�<c(<�����/㼴�J�d����������8��@h�j���H�M4�ѹ���c�����d�@)ἀ�H��<�   �   Lo�<�I=f�M=:�h=,�j=tcV=֌,=�B�<��;@Z�ԭ-�V����rԽ���}*��E���Z�Pg�ҍi�
a��N�|�3��K��~۽Bl������1ٻp|�<6O=��M=��h=��j=beV=ԍ,=`B�<0��;8f�Ʋ-������wԽ!�b�*�n�E���Z�KUg�/�i�U#a���N� �3��O�ʅ۽Ir����� sٻ�   �   �,�0�<0�=$f0=�f>=�4=~�=a�<�d(<`v���(��J�l���������콌��&d���BD��/������߽K���ltd�Dἀ�F�p��<0�,=�g=�%�=�=0-�=0�o=n�8=0�<��;4�r}�gν&����=��lh�����������&��ӏ���Y��e����W���)�F#���X���|!��   �   >g���˻pzu<l��<vn=��=�[�<@F�<��< kg��撼b��D���~��ޙ�"?���l��B�½�3�����y����^����x�I���<���<��E=ꫀ=:��=C��=��=��=���= .<=�p�< �ٻ� /��߮��"	�z\?�܈w�����N��"j¾�rξ�ҾZ�̾6����������~�j�2�1��_��|e���   �   S���\\�@�`���S<��<���<�֫<�us<�t�;`C9���L� 2���,��~R���5���F�`�M�*H�̵4�
��ȼ�`&� ��;H��<�B$=(�d=�>�=�=�=���=�=���=2c�=�7=�ʏ<�.���w�RH�R7.��)p�/c��YȻ��پ�,� �O��tB��Lf�L׾����"ޖ�Dli�-)��2��   �   ����P*N�(g�� �޺�<�/S< �B<R�;��:0���8,�0�|����;�������ȭ�䐘���f� ��@�:�OA<���<��=��P=�x�=h �=aذ=5�=tS�=Z�= �=��=N!�=�.=�<6<�w�#����O�*oS��X��R�����߾�y�EZ�:�y3������D� �Z޾HD��%�����T�8k��   �   I뽯���:��� o������H;�X; q :�n� %����0�H,I�H�D�(l%��%ܻ�/� �|;x@2<���<��<�*=H�I='x=n�=�=��=j	�=�W�=�=|��=���=n]�=�І=�!= ɖ;�k$���ý*^&�>pu��\��=�Ӿ6$ �X��j�#�ӷ-�$1���-��p#�Ҷ�����yԾk���n�{��.2��   �   ��iޫ�J�E�H(ʼ��4�����`�v��Q��x����4�`�E��'6� ���8U��lH;�+<U�<|��<��=nV>=#g=�J�=AԜ=�z�=�d�=��=T�=��=@��=�/�=�1�=���=|��=�x=@����`J���ޫ:��h�� �����)���"�7�3�t�>��oB�s�>�m�3��"��8���꾜������`eJ��   �   v��c��&�d����������L#��
�����RC��A\�X~Y��J2��˻ |�9
<t6�<t8�<��=ʛ@=�ii=��=�֜=�=X��=��=p��=%�=���=�P�=��=�%�=3��=�I�=>T=����:�c�l���G�3O���lþ����P��	,��>�3�I��M�n�I��>�83,�����o��t�ƾ斾p�Y��   �   �
��Ž�|o��q�슘�xk@���$�`^7��W�@�j�Haa��Z2�I�����:p�%<���<�{�<Z$=t7N=�xw=v��=6��=<�=Tq�=P��=���=V��=��=���=Ґ�=l�={�=Aǃ=j_=`�Ȼ�_l����� �L��e��bǾ�����,�HH/�9�A�%GM��QQ��LM�~�A�.~/�9���w��8�ʾG��(@_��   �   b�����J�d�����H���D#�
� ���IC�09\�vY�C2� �˻ M�9�
<�8�<�:�<��=��@=dji=P��=�֜=<�={��=6��=���=8%�=��=�P�=��=�%�=���=�J�=�U= ���6�c�j��G�TN���kþA���IO��,��>�;�I���M�x�I��>�a2,����n��b�ƾ;喾�Y��   �   ���۫�E��ʼX4�0n����v��0�����@|4�x�E��6� �� U���H;h�+< Y�<���<�=�W>=�#g=K�=�Ԝ={�=8e�==��=LT�=�=���=0�=42�=d��=���= |=����[J�9��V�:�Ug�����#�龹��"�w�3���>�nB���>���3�k�"�7�+�꾓�������bJ��   �   UC�����x�(�n� M� I;�mX; �: $n�P���x�0�8I��D��Z%� ܻ`����|;�I2<(��<�
�<�+=P�I=�'x=��=��=T��=�	�=�W�=��=��=���=�^�=7҆=N�!=���;�c$���ý�Z&��ku�,Z����Ӿ8" �����#�G�-��!1�3�-��n#��������Ծ������{�
+2��   �   ����N��T��@�ݺh!<LS<пB<p��;���:�~���d,���|��曼`1���}������8����f�`����I�:�UA<`��<��=z�P=�x�=� �=�ذ=��=T�= �=!�=���=##�=	.=�X6<�d������K��iS�ZU��G����߾�v�aW�7�e0�	������� �rU޾C@��˧��l�T��f��   �   �����C� `���S<$��<p��<��<P�s<���;��8���L�D$�� ���L���5�^�F���M�	H�X�4���ȼ�[&����;T��<�C$=��d=�>�=��=��=���=�=5��=8e�=��7=0ڏ<��	w�M?佌1.�r"p��^��Jû�;�پr&�^ �����;��`ﾞ׾ؓ���ٖ�ei�,')�#)��   �   �W��M˻�u<��<�v=��=�k�< V�<�< �f��ג�N��pD��~�]ܙ��<���j����½�2�����������^�v��h�I�P�<l��<��E=s��=���=��=#��=)�=̕�=�3<=x��<�5ٻ�/��֮��	�KU?�6�w�����H���c¾ilξҾ��̾���������̢j��z1��S���[���   �   h���<��=Xo0=\o>=��4=<�=lp�<(�(<�:��L�6�J�@�������)��t��=c�B���C�T/�$��Z�߽����hsd�|� �F�(�<&�,=$�g=]&�=#�=�.�=6�o=��8=D+�<`z;����`}�w�ͽ^����=�1ch�� ��A���c���� ������T�������W�z�)�p��mM��Fj!��   �   ���<�U=X�M=�h=�j=�jV=�,=�P�<�6�;�>� �-�/����oԽ��d|*� �E���Z�ZOg�>�i��a���N�.�3�nK�9~۽�k������+ٻ8~�<TP=&�M=��h=v�j=
iV=�,=0P�<�=�;�5�&�-����tkԽ���x*���E� �Z�WJg��i�^a���N��|3�@G��v۽�e�������ػ�   �   �,=Ϊg=8(�=��=�/�=��o=��8=�*�< a;���e}�8 ν�����=�<gh���ꮕ�@����#�������V������D�W���)�L��
S��Ts!�0���<�=�k0=hl>=��4=��=�n�<X�(<�0���㼚�J�磓�_��������f_���J?��*���q�߽�����fd�0�ༀND���<�   �   =�=���=T��=��=F��=�3<=�~�<`Gٻj/��ٮ��	� X?�Ѓw����uK���f¾~oξ3Ҿ��̾���������$�j��~1��Y���`��@_��}˻�u<D��<�s=�=xg�<$S�<�<��f��Ԓ�2���
D�H�~�ؙ��7���d��|½�+�������|���^�ʹ� cI�п<`��<��E=�   �   ��=X��=���=�=а�=}e�=l�7=�׏<$��6w�lB佾3.�\%p��`���Ż�ҘپW)�� ����?��)c�t
׾^����ۖ��hi�&*)��-�u����O켠V`�p�S<��<��<l�<P�s<0��; �8�(�L�� ������G�2�5���F���M��G���4�*�P�Ǽ`3&��H�;���<�J$=�d=tA�=�   �   D�=GU�=
!�=�!�=b��=L#�=�.=8S6<�i�����:M��kS��V�����.�߾&x��X��8��1����B���� ��W޾PB������2�T�i����z$N� ]���*޺�<BS<�B< z�;@��:����0e,�ؤ|�P㛼\+��<u��(���P}�� �f� ����I�:(uA<p�<��=��P=�{�= #�=�ڰ=�   �   Y�=r�=ƹ�=��=�^�=B҆=��!=��; f$�B�ý�[&�tmu�N[��E�Ӿ# ����#�{�-��"1�s�-��o#���������Ծ���?�{��,2�7F�L��� |���n�`t���H;�OX; t:�:n�������0��I���D��S%��ۻ ���};�\2<Ŀ�<��<X1=��I=�,x=
�=��=��=$�=�   �   ��=0��=|0�=�2�=���=���=�{=����\J�a��0�:��g������$��U�Ğ"�C�3�x�>��nB���>���3�=�"��7�s�꾩������$dJ����ܫ�L�E��"ʼ��4�Pz����v�;��X���4� �E� 6�x��@�T� �H;��+<�]�<X��<.�=�Z>=L'g=�L�=֜=�|�=xf�=P��=2U�=�   �   \��=4Q�=(�=&�=���=�J�=�U=������c�lj���G��N��lþ�����O�	,�&>���I���M��I�:>��2,�i��No���ƾ�喾��Y���������d�����ԙ���F#��
����`LC�`;\� xY��D2���˻ F�9�
<:�<$<�<��=��@=�ki=	��=zל=��=��=�=��=�%�=�   �   Z"�=�^�=�v�=O�=���=��=��q=��<�Kܻ%T�ؽ�O+��q�9霾Ny���[�����r�����D�x���z���¾���ί|�L�>�y�
�Y1Ľ-���VU���:��@��HZ�r�~��\������/���ҟ��K��"ts�]6��\�P��8 <԰�<��/=�Bm=�Z�=��=	��=&8�=�b�=���=��=�   �   ���=�^�=T��=F��=���=�0�=�r=�b�< $��M�1�ҽ��'���k�ջ��l�����۾V���je��&��e������iܾ�������v� :����y������z�J�f�0�T(6��P�F.t����񚙽ot������.���o�*`4�9ἠ�!�X� <��<�	(=X�d=�ύ=k��=P]�=�)�=���=���=,��=�   �   �t�=�;�=��=L��=��=/s�=�-r=�=�)>�N9��Yýb��(�]�h���Ӝ���5Ͼ�����������צ���}��)Ͼ2.���u����e�F,��4��XF����j�},����R���2�j�U���y�<ꊽ���!�����p`c�,�/���<G�`#�;xY�<,�=��I=��=H��=Y�=���=���=���=c�=�   �   ��=��=���=*��=��=�ߠ=��p=��= �:N���X��z3�XqG��������e���h�о��޾@�%޾�о����@ܟ������JK���ҽ���XQ6������gͼlUؼ����Y'�*eK�HIi��J{���}��Cp���S���+�x���उ���F�Ȃ1<���<T�=�ZO=�ƀ=�R�=�Э=ܩ�=A�=���=�   �   n-�=h:�=^��=�]�=���=���=�k=>�=���;�)�������i,��xb�D��������U��9žze����������"���j]��)��y��t�����J��M�P���V2��J�آ���kڼ8;��33�� K��hV�frT�xF�hn-�����G̼�rm�`_Y��	<�Ѩ<��=bn;=Dcn=m�=by�=�c�=�A�=�   �   ���=̴�=J��=��=-�=ِ=nV_=s
=H�<����B�j���ƽu���<�.�h�R����K���ޠ�?����;����eY��C{]�܄0����=b��d"_��w����E�:@��;��e;@�!��4�t���`�󼐧�΅0�@=�V�@��;�('/���&���¼`j� W�X�<�8�<R=�M=�\�=LӘ=��=�   �   ���=S��=�"�=F'�=���=���=hK=`� = <�s��@[:��ɟ��	罜����:���Y�(Tq�4��Rz��Z�z��)g���J�(�'�t �ݧ��T�f�h��P���� -<���<�Ƕ<�ԣ<��`< O�;P7��T|��(Vۼ�����1�J�J�B$]��Sh��nk�(e��3T���7���,;���~��8�
<\��<@�'=��b=���=�   �   x�q=�7�=��=��=]+�=��_=Zu,=��<�v<`Y�V����~�t��E���j���&��7�>+A���A�֥9�~�(����f���x����V�p(ɼ�XS�,�<@I�<�X=� =F�=��<4k�< (�; ���tǘ���TE7��i�zD��Ȣ��3*��6��8E��
D���♽�}���8���Լ�}����e<�p=��A=�   �   ,� =��I=��^=�>`=��O=.�/=�=�?�< aB;��e�t~�ȤP�g��gr��VQؽ�\�����.�	�T���?��^|�~:������f�+�ҍ�p��;�P�<�� =zJ=��^=�B`=Z�O=��/=*�=lD�<@zB;�e�����P�xi���u���Uؽlb�� ����	����F��;���@��i�����+��㍼`U�;�C�<�   �   <א<�>�<�S=$ =�=ԕ�<�c�<`�;���Xʘ�
���C7�hi��A��7����%���0���?��>���ܙ�\x}���8��{ԼP7����e<vw=l�A=p�q=�9�=z�=ῌ=�,�=r�_=�w,=��<`y<�Y������~������콆m���&���7�)/A���A�ߩ9�Y�(�x�����S~���V��8ɼ U��   �   �)����,<���<��<lˣ<�`<-�;�U�������Zۼ��L�1�f�J�� ]�rNh��gk�  e��*T�Ԉ7����'��06����
<@��<Ԯ'=X�b=�=���=9��=}$�=�(�=���=ǻ�=�K=� =�<(w��|^:�-̟�������:���Y�(Xq�x���|����z��-g�y�J���'�c�ସ�ҿf�Ę��   �   ��伐����:`��;�Me;�3"��4��������h����0��=���@���;�t#/�������¼��i���V��<�G�<%=&�M=s_�=�՘=��=b��=X��=���=��=.�=�ِ=ZW_=(s
=�<`ƴ�:�j���ƽw�N�<�`�h�)����M���࠾x����=�� ��M[���~]�ȇ0���lf��p)_��   �   ~�J��W� ���h2��J������tڼF?��73��K��jV��sT�|F� m-�����@̼�`m��Y��
<�ݨ<��=t;=�hn=~o�=�{�=\e�=C�=�.�=�;�=l��=^^�=���=��=�k=ܭ=��;�.��)�����k,�l{b�̇��m��䐵��W��Qž�g���³�e��������l]�&�)��}������   �    ���U6������oͼ@]ؼh���]'��hK��Li��M{���}�Ep��S���+����ԟ����F� �1<���<��=�^O=�Ȁ=�T�=dҭ=t��=vB�=��=��=Ф�=`��=À�=p�=�ߠ=z�p=�=@�:���Z���4�-sG�8�����������оU�޾��޾0о ����ݟ������LK���nҽ�   �   H��(�j��,����U���2�f�U���y�}늽�򑽦"������`c���/��漘5G��5�;�^�< �=��I=��=���=��=��=��=t��=�c�=�u�=4<�=~��=���=P��=Fs�=X-r=H�=@@>��9��[ý|����]�G���ڝ���6Ͼе�����������~�+Ͼ$/���v���e�j,��6���   �   k���p��V�J�H�0�:*6�� P� 0t���������t������E��Ro�x_4��6�0�!��� <p��<T(=�d=�Ѝ==��=^�=1*�=8��=6��=���=���=�^�=���=p��=���=�0�=<r=ta�< ,���M�?�ҽZ�'���k�[���
�����۾����e�H'�$f�s���jܾ���y���{�v��:����   �   z1Ľf����U�j�:�F@�hIZ���~��\������/��vҟ�mK��Xss�\6��Z�X���#<���<��/=XCm=�Z�=��=6��=L8�=c�=���=��=h"�=�^�=�v�=O�=���=���=N�q=`��<�Oܻ�%T�zؽ
P+��q�\霾oy���[����|�����D�u���s���¾�����|�C�>�z�
��   �   ���������J���0��'6�P�&-t�������`s��i�������o��\4��2��!��� <��<P(=�d=�Ѝ=|��=B^�=`*�=Z��=X��=���=��=�^�=���=���=��=
1�=br=�d�<����M�`�ҽ&�'�Q�k�v�������c�۾����e��&�ve�*����hܾ󽾓�����v�t
:����   �   �D��\�j��z,����P�$�2���U���y�y芽����+��P[c�ޚ/�T漀'G��L�;�c�<��=�I=��=0��=�=`��=T��=���=(d�=�u�=�<�=ظ�=��=��=t�=�/r=X�=��=�	9�Xý6����]�����ٛ���4Ͼ\�����d�������v|��(Ͼ&-��
u��5�e� ,��2���   �   b��rM6�����8aͼ�Nؼ���U'��`K�,Di�"E{�N�}�&=p���S�j�+��z����� lF�P�1<X��<��=~`O=Tɀ=lU�=�ҭ=ӫ�=�B�=h��=B�=:��=���=c��=F�=�=��p=.�=���:T���U���1�BoG�ۍ��C���Ԋ����оŉ޾k�T޾�оꊺ��ڟ�\����HK�P��ҽ�   �   Z�J�4D�ؿ� F2� �J������aڼj5�n-3�~�J�aV�jT��F�Fe-���� 5̼0Mm� �X��
<��<��=�u;=�in=p�=�{�=�e�=�C�=:/�=<�=��="_�=���=s��=�k=��=�'�;���I��?���f,��ub�������������ZS��žQc����������t���g]�e�)��u������   �   Xk� ����:�֭;��e;��!�P}4�������P���|0��u=���@�(�;�/�������T�¼X�i�`qV��<K�<v&=d�M=�_�=֘=v�=慹=��=M��=��=)/�=Nې=|[_=�x
=��<������j���ƽr�N�<�b�h�8�pI��qܠ�ޟ��A9�����\W���w]���0�����]���_��   �   �å��-<`��<Ҷ<xߣ<ب`<���;0���4l�� Dۼ����1���J��]��Fh�dak��e�&T�:�7���h#���'��x�
<���<�'=T�b=yÉ=S��=���=.%�=�)�=��=Z��=4K=�� =X3<8c���Q:�ğ�������:���Y��Oq�l���w����z�%g���J�~�'�A��l���>�f��z��   �   $�<�T�<�]= =Ȓ=��<�x�<0d�;�G��|���n���97�
i��=�������"��:.��[=��O<��Rۙ�(v}��8��xԼ`-����e<lx=\�A=l�q=}:�=+�=���=.�=|�_=�{,=��<x�<��X�`�`�~�+��B���f���&�{�7��&A�[�A�^�9�D�(� ��n�罡r���V��ɼ�wQ��   �   �� =
J=��^=�G`=��O=��/=� =hS�<�C;8}e��t���P��b���n���MؽZ�����.�	����y>��Z{ི9�� ���H�+�Ѝ�`��;\R�<�� =�J=��^=.D`=X�O=v�/=��=tN�<@�B;@�e�jt���P��`���k��Jؽ5U������	�*���7���t�k3��J���6�+������Ӭ;�^�<�   �   �q=�<�=��=R=�/�=�_=~,=���<��<��X����b�~�������Ti���&�Ҵ7�Z*A�8�A�D�9�
�(�������=x����V��&ɼ�&S���<K�<�Y=
 =�=���<�q�<�J�;�\��P���V��D97�i��;����������)��?8���6���ՙ��j}���8�peԼ 軻(f<�~=��A=�   �   T��=���=�&�=�*�=K��=f��=�K=�� =�4<�d���S:�Ɵ���*��v�:��Y�FSq�x��z��ߋz�2)g�`�J���'�: �}�����f�����򥻸-<���<�ɶ<�ף<h�`<pd�;����r���Iۼ�����1��J��]��Bh�\k��e�4T��|7����|�� ���p�
<��<@�'=̏b=�ŉ=�   �   ���=R��=���=��=0�=ܐ=�\_=Xy
=X�<t���P�j��ƽ�s���<�*�h�����TK��~ޠ����h;�����FY��{]���0�i���a���!_��v�p �@^�: ��; �e;��!���4�������󼈢�j0�>w=���@�x�;��/�D����~¼��i�`V�('<pX�<�,=�M=}b�=Tؘ=b�=�   �   �0�=:=�=���=�_�=D��=��=fk=$�=�"�; ��������h,��wb�ޅ��T������HU��žUe��u�����������i]���)��y��<���~�J��L� ��0T2���J������hڼ9��03���J��cV�TlT�F��e-�ޮ�D1̼hAm� �X�p*
<��<|�=�z;=~nn=.r�=�}�=�g�=E�=�   �   ,�= ��=���=���=��=h�=�p=&�= ��:Μ�W���2��pG�����d���*���4�оh�޾�	޾uоn���1ܟ������JK����ҽ���P6� ����fͼDTؼ����X'��cK�@Gi�,H{�
�}�|?p�t�S�d�+��z������@SF��1<���<��=�cO=ˀ=W�=\ԭ=2��=D�=t��=�   �   rv�= =�=D��=z��=8��=Vt�=�/r=L�= >�
9��Xý����]�2�������}5Ͼn�澬�������Ŧ���}��)Ͼ&.���u����e�8,��4��7F����j��|,���xR��2���U���y��銽�� ��/�� ]c��/����'G��P�;�e�<d�=��I=��=(��=�=P��=*��=~��=�d�=�   �   ^��=4_�=���=���=��=-1�=�r=�d�<���M���ҽj�'���k�����X�����۾F���de��&��e�����}iܾ�������v�:����q���t��\�J�>�0�(6��P��-t�v������t�����z���o�0^4�p4�X�!��� <���<�(=d�d=Lэ=ԉ�=�^�=�*�=���=���=��=�   �   �D�=(��=�/�=D�=���=�=v�=p�c=`��<�㈺~��߅��Nm����-��t\����A���M�������[��-���b ����a��v8��*���޽�_�������`ڍ�|l���Ͻ�����R��Z'��A4��9��4���'����|��~���Io��케������<V�<=BT�=E2�=YU�=.�=��=��=�>�=�   �   �%�=��=�8�=h!�=4��=�h�=��=��a= 0�< 7'��z�ꜽ{��2R*�D�W��W��v���T���∞��ɭ������1\��3���.�׽�����|�a��]?���IȽ����7G��#���/�v�4�4�0�H�#����!콩!���Zk��<� i��{�<��8=��=އ�=���=�]�=T5�=Z�=���=�   �   ���=��=�-�=�9�=( �=x<�=�Ж=@,\=(�< ��9b	�{ƒ�e��G����J��q�E���NX��d���b���1���p��tL���%��#�I6ý�͓��+n�:�[�l�n�cH��������޽l����� #��,(���$�Fl����޽����b�`��(�`

��Q�<ng,=��v=�P�=$�=7�=6J�=���=��=�   �   �v�=���=���=:��=E>�=0�=	��=��P=84�<@��:�w�,��tCѽ�[�&�6�bY��t�N���,3��h�����p�)fU�1�3��l��ݽ-ݢ��Cn��B9�ll(���9�p:h�sߕ��6������p�ْ�e����ڏ	������ʽJk��
;S�<�߼pd��L��<`�=`\=��=Ȏ�=�ڽ=h��=�M�=�;�=�   �   �F�=�#�=Jo�=���=���=��=���=4?==t�<@�:�^׼z�h��'����������;�?gR��Z`� d���\�N�K��3�b��]�.����5s��$�<�꼜�̼�V��1 ��b]������ʶ���ֽ_~����������v{Խ�����T��"<H�ph���Џ&<p��<�/3=��n=��=]�=�@�=��=(�=�   �   ���=�n�=�=���=�j�=���=r�`=��= �<@G��ȳɼ�zM��ߝ�]�ս:4�tC���-��8���9��{2��"�`��@��`����p��O�����(Y��ջ#�$!��b����D�q���k���e��IJǽ�˽�ĽT����/���M��ܦF����PP���]R� $p<�K�<�Q3=��i=23�=�%�=�Ѳ=9��=�   �   81�=0��=/^�=�՚=Tt�=N�e=l�/=�\�<|8<�6޻�ռ�=�Ƒ��	����ڽ������	����R3�$[�����ʽ�ߜ��XZ�H�����I��'�:80,<�PW<��$< �;p��<�¼�����V�(\��dt��~���Q(����������|��)U��)��w�P� ?`��,<\��<��=�#S=�(�=fk�=�W�=�   �   Py�=���=���=�,w=S=�+%=�'�< �X<�&ʺ�!�����?�F@{�ڟ���T����ŽcLҽD�ս^�νy4��U���|~�n/�����@+��x?><���<Ȕ�< e=��<4�<��L< d��d��V���"��L�B�k��Z��@ͅ�����<����1y�DOc�H3E����D߼�e���:�<��<҉2=p�_=I��=�   �   
�L=f:S=�H=^�.=�=�d�<��<����\���DX��4$-��U��Wx�$_��Vꔽ6���K����ѕ�I∽|i��&4��u鼈�>��F�;п�<�,=�4=B�L=�?S=P�H=Ƴ.=��=Lp�<x�< ���\����O��6!-���U� Xx�#`��>씽���ä��֕��戽�i��/4���8�>�0�;���<�&=l�4=�   �   |��<�_=`�<4(�<��L< �j�8�d��c���"�\�L�v�k��[���ͅ���������-y��Ic��,E�ʀ�,�޼��d� �:��<P�<��2=��_=���=�{�=C��=���=�1w=�S=R0%=1�<x�X<��ɺ���\���?��A{�����hW��>�Ž�Pҽ��սq�ν�9��`��� ~�2/������c���%><���<�   �   ,<�9W<��$<@�;��,�¼���� W��_��pw��
���2*���������|�,'U�)��m����� �_�x$,<���<��=")S=+�=�m�= Z�=?3�=$��=&`�=�ך=Nv�=,�e=�/=(c�<��8<)޻(�ռ�=�)���V���J�ڽ������	����6��]�
��*�ʽ$䜽�`Z������I� d�:�   �    p��1ջ�&#��-������D�����������Mǽt˽�Ľ����s0���M��n�F���I���IQ� 7p<�U�<�V3=H�i=^5�=�'�=�Ӳ=�=,��=Vp�=��=8��==l�=8��=.a=��= �<�2���ɼ�|M��᝽�ս6��E��-��8���9��~2���"�����~���p�fV�����   �   ���L�̼�a��7 �2i]����ζ�1�ֽʁ����������}Խr����T��d;H��d鼀����&<���<�33=��n=a�= �=hB�=*�=p)�=LH�=�$�=�p�=��=׊�=��=���=�@==��<��:4a׼�h��)��ޏ��k��п;��iR�t]`��d��]��L�63����a꽔����;s���$��   �   fG9�q(���9��?h�<╽�9�����\r�U������̐	����̐ʽ�k���:S���߼�T����<�=8\=:�=.��=�۽=���=�N�=�<�=�w�=���=���=��=?�=��=���=^�P=�4�<���:�z��-��`Eѽ]���6�LY�t�t���Z4�������p�4hU��3�vn��ݽ�ߢ��Hn��   �   P/n���[�@�n�rJ��7����޽������!#��-(���$��l���5�޽������`��&� �	�xU�<ti,=��v=�Q�=}%�=�=K�=X��=��=N��=d��=�.�=p:�=� �=�<�=>і=�,\=�
�< K�9�	��ǒ���R���J�dq����*Y��D���<���2��]�p�1vL�"�%��$�,8ýlϓ��   �   ����V�|�����@��@KȽ-����G��#���/���4���0���#����!�\!���Yk��:鼀<���}�< �8=Q�=���=&��=@^�=�5�=�Z�=V��=&�=p��= 9�=�!�=t��=�h�=��=��a=t/�<�b'��{��ꜽ����R*��W�*X��򋐾����`���B:�����]2\���3���C�׽����   �   n���e��ڍ�m��xϽ2����R��Z'��A4��9��4�r�'��������}��.Ho�����������<L�<=�T�=�2�=�U�=b�=6��=@��=�>�=�D�=>��=�/�=L�=���=�=�u�=,�c=���<����2����m����-��t\����T���M�������[��2���c ����a��v8��*���޽�_���   �   3d�|�$��?��yIȽ6����F�|#�\�/�ƪ4�h�0�d�#���������Wk�46�@��Ā�<@�8=��=∣=j��=x^�=6�=�Z�=z��=D&�=���=@9�=�!�=���=,i�=d�="�a=�2�< �&�\y�B霽����Q*���W�^W���������r���X\���:���0\�e�3�j�g�׽����   �   t)n�0�[�f�n�XG��˟��]�޽�����b#��+(���$��j�����޽������`�� �	��Z�<�k,=V�v=�R�=�%�=��=fK�=���=��=���=���=�.�=�:�=$!�=�=�=Җ=�.\=��< 3�9�
	��Ē�.�� ��f�J�Zq�n���lW����������0��V�p�~sL���%��"��4ýD̓��   �   @?9�i(�T�9��6h�zݕ��4����To�.�������Ӎ	�}���ʽLg��p3S���߼.�����<�=�\=�=䐧=�ܽ=��=O�==�=8x�= ��=���=���=�?�=��=���=t�P=�<�< J�:m�)��@ѽ�Y��6� Y��t�����1��-�����p�dU�I�3�.k�	ݽ�ڢ��?n��   �   (���̼N�`- ��]]����NǶ���ֽGz�t���.�����zvԽ�����O���2H��V鼐x�8�&<��<�63=��n=8�=� �=�B�=��=�)�=�H�=^%�=q�=���=���=��=��=TD==�"�<�נ:Q׼؊h��#��Y������;�QdR��W`��d���\���K�>	3���Y꽺����/s��$��   �   HD�0�Ի��"�|��|��<�D�����/���� ��7EǽZ˽i�Ľ����*��FH��
�F�P��t<�� P� Gp<�[�<JY3= �i=!6�=d(�=BԲ=x��=���=�p�=H	�=褴=m�=^��=,a=�=�'�<@V��P�ɼ�qM��ڝ���սS1�X@�[�-��8���9��x2��"����=����
p�FI���   �   pF,<fW<P�$< S;0���¼�����V�AW��o��ఝ�k"��u������H|��U�.�(��`񼨬����_�H1,<���<��=�*S=�+�=8n�=�Z�=�3�=���=�`�=�ؚ=,w�=��e=0�/=\k�<8�8<p�ݻp�ռ��=�X���=����ڽ4���:�	�����/��W�m��j�ʽcڜ��OZ�����p�I����:�   �   ���<�j=��<�?�<@M< �\���d��D�
�"�FwL���k�tT���ƅ�l��������$y�@Bc��&E��{�0�޼(�d��i:0�<t�<ڐ2=� `==��=$|�=���=���=�2w=|S=�2%=�6�<P�X<�ɺ������?��4{������N��J�Ž�Eҽ��սƳν.��`|~���.����0틻pZ><���<�   �   ��L=�DS=��H=r�.=��=4~�<��<=������:���-�j�U�JKx�yY��d唽����ȝ��ϕ��߈�`xi��#4�`q鼠�>� R�;$«<�-=ڰ4=.�L=�@S=^�H= �.=,�=Dt�<�<�f�� ����C���-���U��Lx�;Y��F䔽�������˕�0܈�Npi��4��a� �>�p��;LΫ<63=��4=�   �   '~�=�Ì={��=�6w=�S=�6%=�?�<`Y<��Ⱥ���r�҅?�25{�ٚ��lP��
�ŽIIҽ��սP�ν�2���|~�� /� ����"��C><D��<p��<�e=��< 6�<�M< ^b�عd��P� �"��|L���k�hV��;ȅ�򺆽_���l"y��>c��!E��u�D�޼P�d� :8�<"�<"�2=�`=j��=�   �   x5�=R��=fb�=8ښ=�x�=�e=��/=r�<�8<�ݻ��ռ��=����Ӈ��a�ڽ����J�	����t2�tZ����F�ʽ�ޜ�~WZ�x�����I��>�: 3,<�SW<��$<`;���h�¼���@�V��Z��:r��ȳ���$��b������*|�U��(�PZ�4��� N_�F,<���<��=�/S=�-�=>p�=Z\�=�   �   ��=7r�=�
�=H��=zn�=Š�=�a=~�=�+�<�+����ɼtrM��۝���ս�2�0B���-�"8�2�9�h{2���"�
����������p�<O�L����V�@�ԻX#���������D�����q���!���Hǽ�˽>�Ľ	����+��QI��F�����8�� \O�xTp<`c�<4]3=�i=�7�=!*�=�ղ=���=�   �   �I�=l&�=r�=���=���=� �=��=F==<%�<@�:�Q׼0�h��$��s���|����;�nfR�*Z`�yd�k�\���K��3�/�v]�䨭�65s���$�L�꼰�̼�U�b1 �<b]�[���ʶ���ֽr}���R������xԽ����!Q��p4H��W�xv��&<��<93=��n=��=$"�=HD�=��=
+�=�   �   y�=���=���=\ �=|@�=��=w��=��P=H>�< R�: n�S*��XAѽ�Z�V�6��Y�Vt�����2��C�����p��eU��3��l��ݽ ݢ��Cn��B9�l(�H�9�:h�7ߕ��6��$�佖p������X��&�	�ݢ��ʽ�h���5S�$�߼�0�����<�=�\=��=̑�=pݽ=���=�O�=�=�=�   �   ��=��=T/�=D;�=�!�=>�=�Җ=~/\=��< K�9N	�Œ��罬��J�J�}q����(X��F���J���1��ƨp��tL���%�|#�,6ý�͓��+n���[�,�n�DH��ߠ����޽N��̢�Z #��,(���$��k�
��m�޽�����`�� ���	�hZ�<�k,=��v=�R�=x&�=�=�K�=$��=\�=�   �   l&�=���=z9�="�=���=hi�=��=��a=@3�< �&�Xy�`霽����Q*��W��W��b���B���ӈ�����������1\���3����׽o����|�R��Q?���IȽ����*G��#���/�X�4��0��#����!�� ��Yk�,9鼀'��8�<��8=��=刣=~��=�^�=,6�=�Z�=���=�   �   ��=�t�=Ё�=��=��=�"�=F�=�u�=��[=.�=xU<hO���;�ʙ�Ěӽ��� ����$��k)��%�+��`��������3���{��ξ{��������w�9����@��hk����������c��w.�������ڙ��.��=Th��R9�2���H���"<����L/�<J�M=U��=A�=���=Ί�=@!�=�=�   �   ���=~%�=��=�S�=��=  �=�=���=8JW=�W=(}<xg����8�I▽�CϽl� �`t��!��E%�� ������T�ܽ����6��0�y���p��P������3<ὄ���<�n�e�xm���^��x⠾֥��9"��T����_��V�c��5�J�tD��d"7�0"���<�L=��=�յ=|��=J��=LD�=��=�   �   xu�=��=�D�=���=�8�=��=>��=�"�=�}H=8i�<�1�;P⌼P1�Q⎽Xý�*��
����]�������ܫ�Ƚ"��:̀��X�<P�8�l��2��#4̽:����-�!�U���z����
���|r��F�������|�`�U���*�z���椽=)�@$һ�q�<H'I=hC�=�k�=���=�Q�=���=��=�   �   �L�=��=�&�=.��=���=�=J�=�p=,�-=�D�<�;�����/(�m����O��nٽ���y��1�U�V.�^�̽�ȧ�U���*K�PM%��[���7�jcv��A���&�2��<�j
_��<{�{��F����������c��A������4��ξ�p���$�<�5A=��=���=� �=h��=��=4��=�   �   `#�=*��=�0�='�= ج=�Ֆ=�{=2fB=�5=xM�<�����Q����#��r��������QԽ1���zֽ�u�����}���;�b��H�ƼF����,�*.������-��j����;�]VU�[�f�a�m��Dj�x'\��(E��'����ƽ�V������;Q����< q2=
5}=F^�=6��= ��=��=�h�=�   �   ʿ�=א�=��=���==�=j�n=8*:=�\=�z�<@gG;�A�|�ۼ�s*��[d��:���~��!���𲱽_���g��>�`�\q"�`�ͼH�Y�0|���j��x���3��j"������
����>[�
+���:�dMB�J�@�*6��$�D]��\������_�����w���<��=�o^=y"�=�|�=^�=B��=�1�=�   �   ��=�Ƣ=�|�=v��=�R=�=�C�<X"5<����u���ۼ�r�F�B���e�����俊�(��矌��߂�j�c�X�4����������Rl��Y�;��]<HHw<�C2<��?:�t�����Yn��{���Y׽S��l<��z��p���@���黽� ���YG��:ἠ�8�9<8�<�s3=l1j=B��=��=L!�=��=�   �   gT�=6�=]= x.=�~�<�h<�m��z���漼+ ��D���^��)q��i{��}�&wx��j�JS�W2���HS������`!�; [�<�L�<З=(=��<h�< 1<�l컨Aڼ`�@���������Vǽ{ؽ��޽�Dڽ;�̽_��䜽�~�4�>������t���%:�̀<�{�<��/=z\=D#=���=g��=�   �   �_N=h�2=B�=p��< 5;H}n� ���A�d�u��J���*��/����f������%��f9p��&J�x��(0ݼ�yi� 9[�0�O<��<��=t�:={Q=��X=&eN=`�2=��=��<��5;pZn�ԃ�fA�>�u�dF��'�����Xd�������%��>:p��(J���H9ݼH�i���\�@�O<T��<N�=T�:=vQ=b�X=�   �   $��<|�<0<���xSڼ�@��Ĉ�����[ǽ|�ؽ;�޽�Hڽ1�̽	a��-圽�~��>����(�t���&:�ր<��<6�/=
�\=�'=�=���=�V�=܁�=��]=�~.=���<H+h< k���y�����$ �
D��^��&q�Rh{�|�}�@yx���j��NS��\2����_��������;�O�<dA�<Z�=�
=�   �   �*2< >:p�t�:���bn�ƀ��r_׽�X��J?�����������Č�e뻽�!���YG� 8�����9<d�<zw3=R5j=3��=��=>#�=��=�=!ɢ=X�="��=İR=�=PP�<8;5<��x�u�L�ۼ�o���B���e��񀽁���p�������₽�c��4�����X��� �l�P+�;��]<1w<�   �   0��DA���q"�צ��}��W��^� +���:�0PB�܍@�d
6��$��^�]^����,�_�x����w����<��=�r^=$�=�~�=��=��=j3�=���=���=��=(��=��=8�n=$/:=la=ȃ�<��G;�A�4�ۼ�s*�]d�3<�����������H���տ�������`��w"�X	μpZ�@��� ����   �   輊",��1��!���B2������;�(YU�$�f��m�4Gj��)\�R*E�d�'����ƽ2W��P���(Q�|��<2s2=x7}=�_�=vµ=k��=(�=�i�=�$�=���=J2�=��=�٬=zז=:{=�iB=�8=LR�< w��HP��l�#�t!r�2�������SԽ3�M���ֽy��<���}���;����ȿƼ�P���   �   ��7�iv��D��?*�:�>�<��_�f?{����h���������c��A�Z�R�(5��|������&�<|7A=��=���=��=h��=��=4��=�M�=��=�'�=f��=�=e�=��=�p="�-=|G�<��;�����0(�xჽDQ��wٽW������2���31��̽-˧������K��Q%��`��   �   F�l�65���6̽����.���U�k�z���������Qs���F������t�|��U���*�̷�� 椽n<)� һ|t�<�(I=&D�=�l�=���=�R�=T��=2�=*v�=8�=�E�=���=�9�=��=��=E#�=H=�j�<�2�;H㌼�1�E㎽�ýT,���
����^�ڻ���ޭ��Ƚ�#���΀���X��?P��   �   R��&���>὆���<���e�n���_���⠾F����"�������_��l�c�Ԅ5���C��:!7��,�<\�L=���=ֵ=���=���=�D�=  �=���=�%�=���=�S�=��=� �=j�=B��=�JW=�W=X|<�h��z�8��▽uDϽ� ��t��!�bF%��� �+��x�i�ܽ����7��t�y�6�p��   �   D��d���x轶��J�@�!ik�̈́��·���c��u.�������ڙ��.���Sh�"R9�����G��!<�`��2�<n�M=ѵ�=�A�=܌�=��=v!�=0�=	�=u�=��=��=��=�"�=<�=qu�=r�[=��=�S<�P����;�iʙ��ӽ҉�&����$�l)��%�B��v��C��H����3��%|���{��   �   �P��{���#<�p���<�$�e�Dm���^��⠾\����!������$_���c���5�"�[B���7��0�<��L=(��=fֵ=B��=���=�D�=& �=��=&�=���=(T�=*�=� �=��=���=�KW=Y=`�<@d����8�]ᖽ�BϽ� ��s�l!�,E%��� ���j�u�ܽ���6��l�y�>�p��   �   p�l�2��#3̽���4�-�,�U�d�z�Q���8����q�� E�����y�|�Z�U���*�����⤽�7)� �ѻpz�< +I=E�=Vm�=4��=
S�=���=z�=hv�=|�=F�=���=:�=��=���=$�=�H=�o�<PM�;�ڌ�h1�8���'	ý[(�П
����y\�������ө�KȽ� ���ˀ���X�2:P��   �   ��7�,`v��?��z$���}�<��_��:{�N������p�� ���c��A�3���0������T��(/�<�:A=��=凩=U�=���=���=���=8N�=P�=4(�=ҽ�=��=�=f�=p=��-=�N�<�0�;@�)(�A݃�hL��ٽf����
��/���5+��̽Ƨ����2K��I%��X��   �   L���,��+��/���W*��w����;��SU��f�P�m��Aj�>$\�h%E�
�'��W	ƽR���� �P����<w2=h:}=�`�=Põ=��=��=@j�=(%�=��=�2�=R �=~ڬ=@ؖ=<	{=BlB="<=[�< ����B���#�~r�m���9 ���LԽ��ʿ�^
ֽ�q�������}�F�;�^�h�Ƽ�=���   �   Xx��)��`d"�D���������X�.+���:�JB�ˇ@��6�T$��Y�>V�*�����_�l���#w��
�<��=v^=M%�=x�=��={��=�3�=���=0��=�=���=6 �=�n=T1:=<d=$��<��G;�A�P�ۼ|j*�VRd��5���y��-鯽!���'���˷��)��z�`�Tj"���ͼ��Y� S��@D���   �   pX2< %A:��t����jQn��v���T׽M��)9�������3|�?��)㻽���4NG��%ἐ�񻨲9<,�<�z3=�7j=3��=��=�#�=3�=��=�ɢ=��=���=�R=Ƨ=�T�<�F5<���h�u�\�ۼh���B��e��뀽�������������ڂ��c���4�h��� ��� �k� ��;X�]<]w<�   �   ���<��<�I<�4�p1ڼ�@�H������HPǽ�tؽ��޽�=ڽ�̽�W��Pݜ��	~��>�����t� G(:@߀<���<��/= �\=V)=���=A��=XW�=Y��=��]=�.=D��<�1h<��j���y�|��N  �bD���^�q�^{���}�lx�T{j��?S�$M2�x��A��@^���Z�;h�<XX�<P�=j=�   �   NjN=��2=��=���<�6;7n��y�N A�0�u��?��M ��7���c]��ӄ�����2-p�lJ�R��,#ݼ`ei� =Z�P�O<���<\�=ܮ:=B|Q=��X=fN=L�2=��=��<��5;�Tn� ���A��u�eD��y$��񙞽~`��#���@ ��`.p��J�d��8ݼ0Vi� +Y��O<���<��=�:=b�Q=��X=�   �   CY�=e��=*�]=��.=К�<�Kh<��h��y���� ���C�8�^��q�([{�t�}�plx�>}j��BS�ZQ2�\
�XL��0����1�;@^�<O�<�==���<�<X4<�e컘?ڼ�@�ľ�����ZUǽ�yؽ��޽Bڽ��̽[���ߜ�B~��>�D�� �t� �(:��<|��<V�/=��\=�,=\��=��=�   �   7�=eˢ=؁�=��=�R=(�=X`�< _5<�!���u�<�ۼ�c�ƌB���e��뀽^���i ��ۜ��%݂���c�h�4����(��� =l�Pb�;8�]<xKw<`F2< �?:`�t����Xn�{��FY׽ER���;�g
����V�u~���滽����PG�0'�0��x�9<\#�<^}3=�:j=���=-�=b%�=��=�   �   \��=���=��=���=6"�=@�n=�5:=�h=@��<@2H;��A��{ۼ�h*�Rd��6���z��믽��������Һ��7��p�`��o"�(�ͼ��Y�@v���e�����2��xi"�:���Y
�����[��	+�m�:��LB���@�P6��$�\��Y⽴���Z�_�8�� .w���<��=�w^=E&�=���=��=���=25�=�   �   0&�=*��=4�=�!�=
ܬ=�ٖ=�{=�oB=x?=a�< z��X?��n�#�r�S�������NԽFὋ��Qֽ�t��d
����}��;�����ƼE���輞,��-��ǫ��k-��H����;�*VU��f��m�HDj��&\��'E�'�'���ƽT����� �P����<bw2=>;}=Ca�=ĵ=���=��=:k�=�   �   �N�=�=)�=־�=��=?�=��=�p=F�-=�R�<0=�;p쒼�)(��݃�SM��lٽ;������0����-���̽5ȧ�����K��L%��[�<�7�cv��A��q&���<�T
_��<{�c��(������R�$�c��A������2������c��0-�<^:A=��=.��=��=x��=��=8��=�   �   �v�=��=�F�=���=�:�=��=p��=�$�=��H=xr�<PU�;�ٌ�j1������	ýd)�x�
����T]�~���������Ƚ�!��
̀���X��;P���l��2��4̽0����-��U���z���������mr��F������6�|���U� �*�Z����䤽R:)�0һ�w�<B*I=�D�=am�=T��=NS�=���=��=�   �   6��=8&�=���=lT�=��=$!�=�=��=�LW=�Y= �<@c����8�nᖽ�BϽ� �t��!��E%��� �v����1�ܽv���6���y���p��P�����"<�{���<�b�e�vm���^��r⠾Υ��/"��D����_��$�c���5���C��!7�����<��L=Ԧ�=2ֵ=0��=���=�D�=< �=�   �   4s�=,��=Pb�=�p�=�
�=�r�="ܷ=�d�=N�=��W=�!=H߮<@��;�S����t�1�`L_�n�{�M���h�|��|e�@LF�44(����7��<��������R��tA��F���|��Ľľ����������	�0��D4�������þ�Z����w���1��h佘^j���:� ��<�Re=��=zd�=|��=��=�G�=�   �   �=���=��=���=B��=���=k�=J��=�d�=�JO=�=�W�<`�\; �X�����l.���Y� �t�0�|�8Is��[���<�,���/����@�2�b�}����T}�9�<�H�z�����Q���O[߾D��(�!���!��C���a߾~�������r�L�-�B�޽f�b���'�8��<�f=x��=���=�]�=r�=>\�=�   �   ���=��=� �=�!�=]��=q�=�a�=���=��i=.�4=��<P�}<  �9�m�8 ��%�~J�p`�|gd�VX�ܔ?��\ ����������
>�<�\��Ƨ�V����e.�	si�a�������]�Ѿ�|�����Z2������<{Ҿ�ܴ��͓�7�c�x�"�=rν��L�Г们V�<��g=·�=�&�=���=���=$r�=�   �   j��=֍�=$��=(��=��=��=?%�=�g=\R7=�N=(��< ��;0����ڏ�(T�ة�`:5�p'B��@��/�X����Ư��R����ͼX�(��}��2OӽAD��N��Ǆ�]A���%���Ҿ'�ྺ澝��[�Ӿ&���C���Tu���M��n�̵�f�+� +��l�<��h=�U�=t{�=��=Z�=p/�=�   �   ���=+��=F��=!��=�v�=�|=N�L=n�=�P�<�x<�k�; Z���v� ����9��@p����X� �,��P.��HL���Z}��=�@�y�0=���U-���̼x�E�>䤽-?��:�,� 0a��ۊ�Ԣ�J/��d�¾��Ǿh�þ�*��Җ��T���Pg��0�-���")���� �E;�=�Vg=�Ù=���=n�=���=(3�=�   �   T5�=&�=�1�=!9�=�V=�=XU�<��P<�?�:��tڐ���ɼP4����
��&�zY�����h���ּ�阼#��q�����;H6<��;<���;�7ӻ�%ڼ�`��h���H�6�3��"a��O��d!��wS��~��������a�����Įl��f@�j��y�˽T�r�pH�����;J�	=0~`=�=E�=��= �=�-�=�   �   ��= A�=�Og= �,=p�<xG#<p;���褼���x�)��'C���P�|�S�*DM���>���)�?���ڼ(	����Q;8MV<�H�<tv�< ��<�y�<�#X<�ox� R�B�j�u���~���*��M�KPj�p�}����X���*t�q$\�<=����N�����t�:����X�-<
�=.R=�~�=$ś=Rƨ=�z�=���=�   �   @�v=��E=�=(�l<����0�Ѽ��6�Flz�]������Kΰ��s������c��������Q��Z� \ͼ�<� ]�:�%p<��<n|=ғ)=tN2=rZ'=�A=�w�< G ��]ͼ��[����+�뽒����*��;���C�ΨB�
�8�1�'����}�:R���x����h�-��3<�>�<�:=��l=[B�=��=�e�=Iы=�   �   VM&=�j�<P�;����BN.�'W��s⹽K��/�����@	��&�'�򽏃Խ:G���ш���@���h���g<���<�~=��B= �`=n�n=�dj=�kR=�S&=py�< d�;�吼�B.��P���۹��ί'��z���=	��#�D��ԽqD���ψ���@�����_<l��<`{=0�B=�`=�n=�_j=
fR=�   �   j�< P�(qͼ[��Ĭ�U��v����*�,�;�ĲC���B�c�8��'�^��[�콊T����x������-�3<�B�<B:=��l=D�=��=h�=�Ӌ=��v=<�E=R= �l<�I��X�Ѽ��6�`z�>���)�Ȱ�$o������k��������Q�"Z��]ͼ �<���:@p<x�<Rx=x�)=�I2=&U'=�;=�   �   ��x�hc�p�j�{�������*��M��Tj��}�F	���Z��6.t��'\��=�����齠!�� �:����p�-<��=N	R=��=�ƛ=�Ǩ=�|�=� �=h��=�C�=Vg=L�,=h��<�k#<��Ԥ�ڡ�|)�(C�b�P���S��?M�d�>�֋)��?���ڼ���P�@�P;@<V<�?�< m�<��<tn�<�
X<�   �   �4ڼx`�n���K���3��&a��Q���#���U�����������c������R�l��h@�ώ�F�˽D�r��I�����;n�	=�`=�=q�=��=��=y/�=J7�=j�=&4�=<�=��V=�=�d�<�	Q<�3�:���͐�L�ɼ(,����
��%��Y����8k� �ּ0񘼐##�@��� ��;856<��;<pq�; jӻ�   �   ��E�p褽*D��)�,�]3a�p݊� ֢�h1����¾��ǾT�þ`,��F������|Rg�_�0�����*�������E;Ґ=*Xg=�ę=���=��=���=�4�=D��=��=J��=k��=qy�=��|=�L=6�=\�<��x<0��;0=����v�@��� 9��4q����� �����5��`T���k}�(O��z�`c���j-���̼�   �   ����Rӽ~F���N�Ʉ�C��I'����Ҿ���z�8����ӾR���2���v���M�Vo��̵���+� %�tn�<��h=.V�=5|�=� �=�Z�=x0�=���=(��=���=ԛ�=��=��=C'�=&�g=DV7=bR=�<���;�u��xُ��T�,��h<5� *B�@���/����x$��ͯ�����lZ���ͼ��(��   �   Cɧ�q���lg.�/ui�����ô���Ѿa~�G����3��.�����{Ҿiݴ��͓���c���"�TrνR�L�P�付X�<��g=^��=y'�=d��=���=�r�=���=��=��=�"�=���=��=Kc�=�=�i=D�4=`�< �}< d�9P�m���4�%��J��`��id��XX���?��_ �|�����p���A���\��   �   ���r~���<�âz�U���0���0\߾����w���!�YD��*b߾��������r��-���޽(�b���'����<�f=��=��=^�=��=�\�=��=>��=X�=&��=���=l��=�=㈜=be�=�KO=��=\X�<��\;p�X����m.��Y���t���|��Js���[�P�<����1������2���}��   �   �����2uA��F��@}�� �ľe����������	� ��4��_��y�þ�Z����w��1�Kg�N\j���:�\��<RTe=X�=�d�=؅�=��=�G�=ds�=V��=vb�=�p�=�
�=�r�=ܷ=�d�=;�=��W=�!=\ޮ<0��;�S�����1��L_���{�����Կ|�$}e��LF��4(�Ȝ��8���<�畄��   �   ���h}�D�<�@�z�p���%���[߾��������6!�C�� a߾������)�r���-�ظ޽N�b���'����<�f=v��=f��=D^�=��=�\�=��=d��=t�=P��=��=���=C�=,��=�e�=�LO=�=`[�<��\; �X�P��@k.�,�Y�~�t���|��Gs���[�h�<�X��H/�L��$�2���}��   �   �ŧ�z���e.�Hri�߸��"�����Ѿ�{龻���1���������yҾs۴�T̓���c�z�"��nνڴL��l��^�<��g=:��="(�=��=
��=4s�=���=�=��=#�=���=�=�c�=���=��i=�4=��<�}< �90�m�p��~%�dzJ��`�dd��RX��?�4Z �<�����`�缄<���\��   �   d|��nMӽ*C���N��Ƅ�J@��5$����Ҿy���澷��n�ӾF�������s���M�@l��ǵ�(�+� ��w�<0�h=bW�=}�=L!�=~[�=�0�=���=~��=��=,��=�=0�=�'�=��g=0X7=�T=L�<��;�P��pΏ�HH����45�"B��@�L�/����(�����鋼@L��0�ͼ��(��   �   R�E��᤽+<��b�,��-a�0ڊ�yҢ�p-��\�¾t�Ǿ*�þn(������K
���Lg���0�s���5$������7F;�=\g=ƙ=���=Y�=���=5�=���=\��=���=؅�=�y�=��|=x�L=�=�`�<p�x<���;�����v�8���*���h����|� ���X"��XA���F}��+�`�y����PG-�(�̼�   �   �ڼ�	`�Me��^F���3��a��M��Z��<Q��!���(���]_������j�l��b@�މ�D�˽x�r��5����;4�	=,�`=��=��=��=:�=
0�=�7�=��=�4�=�<�=��V=N�=�g�<�Q<@��:P���Ő�\�ɼ8 ����
����P�(���`���ּ�ۘ��"� ���P��;�Z6<x�;<���;�ӻ�   �   @x�|EἮ�j��p���{���*�0�M�Lj��}����V���%t��\��=����	�齄��v:���ا-<��=�R=���=�Ǜ=�Ȩ=K}�=T�=�=dD�=
Wg=<�,=���<�p#<@⾻�Ф�T���x)�0C�r�P���S��8M�:�>���)��5���ڼ8���0��`oQ;8eV<dS�<���<���<��<�7X<�   �   $��< Q���Nͼ~�[�����غ������*���;�&�C��B�^�8���'�̺�v�K���x�r����-��*3<�N�<�
:=�l=NE�=� �=�h�=Rԋ=��v=0�E=>=��l<�A���Ѽh�6�@^z�����쨽 ǰ��l��������������Q��P��Iͼ��<�@M�:�@p<̋�<�=�)=RS2=@_'=�F=�   �   (Y&=���<���;XԐ��8.��J���Թ���ά��@��J9	�O�׾�wԽ�<���Ȉ�@�@�� ����<���<��=� C=N�`=(�n= fj=�lR=�T&=8{�<�j�;�㐼�A.�>P���ڹ�I�ό&������<	��"����|ԽA��̈�f�@���������< ��<��=C=��`=&�n=zij=xpR=�   �   ��v=�E==hm<� ��H�Ѽ�6��Rz�!����樽'���fg��&���������Q�"N��Gͼ��<��$�:�8p<؆�<=�)=�O2=�['=�B=�y�<  �t\ͼ֋[��������P����*���;�5�C�"�B�0�8�&�'�ѽ�{��N��ğx�4���-��'3<$O�<�:=|�l=ZF�=�!�=Lj�=	֋=�   �   ���=xF�=\g=&�,=<��<�#<����������,o)��C���P�J�S��2M�ھ>��)�p4�ȵڼ����`���DQ;8YV<M�<�y�<���<�{�<H'X<@dx��Pἦ�j��t��Z~���*���M�Pj�"�}����EX���)t��#\�8=�f���������z:�X��8�-<�=R=��=�ț=�ɨ=�~�=��=�   �   49�=��=�6�=�>�=2�V=��=pu�<(/Q<@w�:��������ɼl����
���$O����a�x�ּ�����#� "��0��;�M6<�;<`��;2ӻ�$ڼ.`��h��hH��3��"a��O��N!��ZS��[���d����a��������l�f@�[���˽.�r��=��p��;��	=ڃ`=��=$�=��=0�=61�=�   �   ���=���=J��=���=|�=��|=ȏL=��=l�<��x<�ג;�󸻈�v������&��Dh���� ����'��PG��`S}�8�@�y��6��HS-���̼�E�䤽�>��#�,��/a��ۊ�Ԣ�</��T�¾��ǾI�þ�*��������Pg�Q�0�n���6'���� 
F;T�=F[g=�ř=5��=��=:��=�5�=�   �   ���=l��=��=���=��=��=�)�=��g=B\7=�X=��<,�;�<�� ˏ��F�$���55��#B��@���/����X�į�X�P����ͼ��(��}��Oӽ1D��N��Ǆ�VA��z%���Ҿ�ྮ澌��?�Ӿ������u��M� n��ʵ�~�+�`��s�<�h=W�=}�=�!�=�[�=v1�=�   �   D��=��=��=�#�=���=4�=�d�=ʩ�=.�i=��4=��<p�}< ��9��m�X��(~%�{J��`�zed��TX���?��[ ����p���缴=���\��Ƨ�=����e.� si�^�������X�Ѿ�|�����U2������({Ҿ�ܴ�x͓���c��"�`qνȸL�0���Z�<��g=Ը�=�'�=��=4��=zs�=�   �   ��=���=��=���=|��=&��=��=Չ�=nf�=�MO=8�=�]�<`�\; �X�X��k.�H�Y��t�B�|�vHs�h�[��<�ܤ��/�x���2�8�}����M}�0�<�D�z�����P���M[߾C��'� ���!��C���a߾s�������r��-�غ޽��b���'�@��<�f= ��=��=^�=��=�\�=�   �   ښ�=<(�=��=�y�=*2�=���=�P�=�֠=[ێ=Vy=��S=NW.=�$	=�$�<ܘ�<��(<�ݱ;`O);�:�:`R;`v\;��V; ��8��t�ͼ��U��������U]�ğ��!Pʾ2���)m��S/���A��NM�`Q�
TM��A�dB/�W*������Ǿo��Q|N��u���\u��w�@�=���=�̯=��=��=���=�   �   ���=Ȕ�=��=�d�= d�=�|�=�^�=e��=片=��j=R�F=�j"=�0�<�n�<�8<}<ת;`�:;�(;��[;��;�ś;@��:�Jۻ�n��kK����8��>�W��<��ƾ����N{�m,�-�=�T�I��M��I�i�=���+��I�����'�þ# ����I�F���jl�pXٻ�_=H�=P��=�E�=�K�=���=�   �   D0�=F��= ��=F��=�º=��=�9�=�y�=$Pb=�?=҃=(K�<D޿<@D�<xA9<�&�;��;`a;Ċ;�9�;�<X�<��;�ȱ�h�����,��������sH��i��d��D�Q���a"��w3�m>��VB�/�>�.�3�P�"����B��R��x���R<�Y��Q��W$�R�=%�=F�=���=���=g�=�   �   >��=��=pp�=Dǰ=l��=<]�=�c=�:=��=|1�<���<ht<�"<���;��^;��;�P
;��p;@^�;h &<�]<��y<��`<p��;`P��h��U	��e��80��8z�W ��rӾ�A��a`�� #�4P-�=�0�}-��r#�h��� �D�Ӿ̍���Kv���'�S�ƽfM)� �p;��=jr�=�֭=��=���= G�=�   �   X��=VB�=ޗ�=Z�=ޑb=j-=8��<ક<�\
<�!:�g����� �,��(.����@ ӻ�u"��\&;(|<�Jj<,�<4�<��<PƎ<@�;x)}��=����?s�NmS�������?�ݾ�` �sm����:��u�����0�!s߾�b��O��[�S��������F𼨿4<��.=�4�=^��=�t�=�=��=�   �   ��=���=z�p=2=`5�<�+< =��,�h����>n(�B+�$w!�"����㼰r���/�������
<�<���<���<��=@H�<H�<@��:Aͼ�|��8ݽ �'��h�������־�P�$���������9��ؾ����ڙ��[o�g�-��'��t�p����	�<p�<=WM�=V�=lo�=0Ӻ=�,�=�   �   @��=v�O=j�=�M<�[�����`MM��ǈ��(��;8��Fl��q?����������m\�*��8��� �п�;p��<�k�<t_=^�+=6�'=�u
=���< |0����R�����f�/�e�h�ѐ���쩾nC��ڣ˾��оu;*&��G$��Z��� �u��}=��F�������&��x��t��<6F=Ѯ�=���="��=�ԥ=�=�   �   ڸ6= #�< z�:|�̼8Y��$���ؽ������]��E�������F_�E���M���:;-��b�� ��� t�<�i=83=L�N=bU=�*D=L=�|�<�:��t���������h�'�xBU���~�⏾����|��S�����ne��K9e�Z�:���Z%ǽ@�n���¼��;��<�H=�=�J�=`}�=��=�kr=�   �   |�<�s����1#����ֽ̢��{0��-K��c]�<�e�0 c�ԛV��}A���%��W��fʽ���Ȇ�$��#[<��=gB=�j=��}= y=��[=\N%=@�<�&��Jy�?����ֽ<���v0��(K��^]��e�&c�>�V��yA�)�%�EU��bʽ���`��P$�(%[<�=jeB=��j=n�}= �x=|�[=�G%=�   �   @���.�9���N���'��GU�S�~�叾������.���
���g��=e�b�:�N���(ǽ��n���¼`�;���<�H=�=L�=0�=�=dqr=ƿ6=�3�<���:�w̼lY������ؽ���{��<Y�LA��������Y����� ����6-��]��  ��ps�<Dh=
 3=^�N=p^U=&&D=nF=�n�<�   �   "��aX�������/�E�h�����𩾦F��#�˾��о�;�(���&��b���^�u�p�=�`H�,����&����<��<�6F=���=���=���=�֥=P��=.��=��O=�=��M<H.�<����?M������!��1��ue��I9��4 ��`���6g\�j��D���x����;���<�g�<�\=�+=@�'=�p
=x�<@�0��   �   H|��>ݽ��'��h���ڹ��+־T�]'������"��f<��ؾ���ܙ�C^o�'�-�6*㽺�t�H���H	�<�<=�M�=>�=�p�=�Ժ=�.�=j��=Չ�=T�p=2=�G�< ++<�娻tڙ�l~����c(��+�&o!�������4l�� �.�@���P�
<��< ��< ��<��=�?�<0��<@��:4Pͼ�   �   ���v��pS����l�����ݾTb ��n�?�����������1��t߾\d��2P���S��������@H��4<H�.=5�=��=�u�=P�=r�==��=�D�=���=t�=ܘb=�q-=���<��<@
< ,#:�)����� �,� .������һ@i"��Y&;�w<�Cj<l�<\ �<�ٹ<<��<���; A}�d�=��   �   4i�_;0��;z�7��FtӾD���a��!#��Q-���0�E~-��s#�I��� �^�Ӿ�����Lv���'��ƽ�M)� �p;F�=�r�=P׭=��=���=HH�=���=Q��=gr�=�ɰ=���=`�=��c=$�:=�==�<���<�1t<x�"<��;�_;��;�R
;��p;�S�;&<�]<�y<@�`< ��;`s軨s������   �   ���FuH�Bk�������F�D���b"��x3�j�>��WB��>�ߝ3��"�l����{R������R<�+Y佮�Q�@M$�8�=�%�=�F�=���=R��=�g�=B1�=r��=t��=���=zĺ=��=�;�=�{�=�Sb=�?=�=�P�<��<xG�<PE9<P)�;��;`a;P��; -�;`�<��<p��;�(������V�,�~����   �   �����W�r=��'ƾ����{�,���=��I�h�M�w�I���=���+��I������þ ����I������l��Mٻ�`=�H�=ֺ�=VF�=FL�=*��=���=x��=���=pe�=�d�=v}�=�_�=U��=ʊ�=��j=��F=�k"=$2�<�o�<x9<X|<Ӫ;@�:;�;��[;p�;���; _�: \ۻ�s��vnK�����   �   `��V]�H����Pʾ����lm�!T/�ÎA��NM�`Q��SM���A�+B/�*�t�����Ǿ���b{N�.t���Yu��n��=@��=kͯ=$�=x��=,��=��=r(�=�=�y�=J2�=���=�P�=�֠=Pێ=&y=��S=�V.=$	=�#�<���<��(<�ر;�F); '�:@H;�k\;��V; ��8����ͼ��U�לּ��   �   n��p�W��<��ƾ����0{�9,���=���I�o�M���I���=�$�+��H������þ-���^�I�����l�0<ٻzb=7I�=B��=�F�=�L�=X��=���=���=̾�=�e�= e�=�}�=`�=���=
��=>�j=��F=�l"=|4�<�r�<�?<H�< �;`
;;�9;��[;`!�;pʛ;@��:�Jۻ�n���kK�����   �   ����rH��i����D����Ja"� w3��~>��UB�1�>�'�3�L�"���~��P�� ��RP<�gU��Q�`
$�B�=�&�=mG�=*��=���=Lh�=�1�=���=���=��=�ĺ=�=<�=�{�=�Tb=� ?=��=\T�<,�<�L�<0Q9<�C�;�;�Ja;�ي;M�;X�<��<���; ���<�����,�.����   �   rc彼70�7z�g����pӾ"@��w_�|#�O-���0��{-��q#���� ��Ӿۋ��~Hv�8�'�؞ƽF)� �p;��=ot�=nح=��=4��=�H�=��=���=�r�=�ɰ=L��=a`�=��c=@�:=b�=l@�<Ŀ�<<t<��"<�!�;�__; .; �
;@�p;P�;8/&<�(]< �y<��`< ��;�>�Xd�����   �   �����q�WkS�a��m���O�ݾ�_ �&l�A���������>/�Up߾k`���L����S��������T5���4<t�.=�6�=z��=�v�=�=�=���=E�=횢=��=��b=�r-=���<���<��
<��#:p��x��x�,��.���0�һ`
"�@�&;Б< ^j<��<��<l�<�̎<�8�;(}�8�=��   �   |�^5ݽ��'�� h����ش���
־�M�� ��V��t��I6��ؾ����י�7Wo�|�-�L!�~t�x�����<��<=P�=��=�q�=�պ=r/�=�=N��=,�p=�2=DI�<�.+< ݨ��י�{���$a(��+�Bk!���X��l`��H�.��ĕ�h<d&�<���<���<��=�O�<��< -�:�7ͼ�   �   ����N����T�/���h�����^ꩾ�@����˾<�о;�"��!��h�یu�[y=��B�"�����&�0.����<�<F=Ʊ�=T��=Ԇ�=hץ=���=���=t�O=½=��M<�*�\����>M������ ���/��0d���7��C�������a\����l����
����; ś<�v�<Nd=��+=x�'=�y
=��<`(0��   �    �����Ǟ��xz򽻛'�>U��~�Bߏ����wy�������hb���3e�T�:�����ǽ6�n�̚¼�j�;���<֩H==�M�=M��=��=�rr=��6=�5�< ��:v̼�Y�g���ؽ4�����X��@�@������W�y���W����0-��P�� P��p��<\o=J3=�N=|fU=/D=�P=���<�   �   ���<�鐻�o�����ֽ<��^r0��#K�Y]�,�e�Uc���V�tA��%��P��Zʽ����v���#��I[<��=nlB= �j=��}=6y=.�[=�O%=,�<����x����{�ֽ���v0�p(K�B^]���e��c���V��xA�8�%�.T�w`ʽ&��r}���#��>[<��=$lB=��j=��}=py=@�[=�S%=�   �   ��6=�A�<@��:@c̼XY������ؽ�����>T�><� ������Pུ{�������)-��F�� ܛ��<�o=�3=ĮN=�dU=�,D=vM=�<�3�����^���7��@�'�PBU���~��᏾����z|�� �����e���8e�r�:����#ǽ0�n�(�¼�L�;���<ڨH=='N�=;��=.�=Fvr=�   �   ���=��O=>�=�N<�P���2M�,�������(���\���0����������X\�h��������
�
�;�ƛ<�v�<vc=N�+=b�'=w
=���<�m0�,��YR�����H�/�F�h����쩾\C��ţ˾w�оS;�%��$�����e�u� }=��E�����:�&��R��@��<&;F=���=���=|��=إ=|��=�   �   ���=k��=v�p=J2=�X�<@R+< ���(�pd����U(��*��a!������V����.��y���<�&�<X��<@��<X�=�K�<��< ��:�?ͼB|��8ݽ�'��h�z������־�P�$���������9��ؾ���<ڙ�0[o���-�=&�\�t�誇���<��<=�O�=��=2r�=gֺ=�0�=�   �   ��=�F�=���=P�=��b=hy-=���<�Ε<��
<��%:PӦ���P�,���-�ؐ��һ �!���&;h�<�\j<��<0�<L�<Ɏ< '�;�&}�~�=�����$s�8mS��������6�ݾ�` �qm����6��p�����0��r߾�b���N��ѳS���Z���(@���4<�.=F6�=F��=w�=��=��=�   �   ޟ�=΂�=.t�=�˰=j��=�b�=8�c=�:=p�=�L�<�˫<`Rt<`�"< C�; �_; U; �
;��p;��;x-&<�%]<�y<��`<��;�J��g�� 	���d彺80�t8z�Q ��rӾ�A��_`�� #�6P-�>�0�}-��r#�b��� �&�Ӿ����lKv���'�f�ƽVK)�@�p;�=�s�=ح=��=x��=TI�=�   �    2�=\��=���=%��=ƺ=��=�=�=�}�=�Xb=�$?=h�=�[�<��<R�<�Y9<�P�;@
�; Ra;�ي;�J�; �<�<���;@���|�����,�������sH��i��a��D�Q���a"��w3�m>��VB�.�>�,�3�L�"����2���Q��\��PR<��X佰�Q�`A$���=�%�=�F�=���=���=�h�=�   �   ���=֕�=(��=f�=�e�=V~�=�`�=t��=��=L�j=��F=�n"=�7�<�u�<�D<@�<��; ;;`=;��[;P!�;�ʛ; ��:0Hۻn���jK����2��:�W��<��ƾ����M{�l,�-�=�U�I��M��I�i�=���+��I������þ ����I�����l�@SٻT`=nH�=���=UF�=XL�=T��=�   �   ���=��=t�=���=`�= Ʊ=��=x�=$��=�-s=V�^=6�M=�?=�75=|�-=X�)=Ƽ(=n�)=��*=��(=��=�-=db�< �~��v�L���F��Xkf���}��,�ݨ:�*)^��}�g���m��_2��Wl��@_����}���]�L:�tD�ŵ�Ǔ��J�X�>���X����:8],=�=�=:��=0��=p��=�   �   LJ�=�=D��=f9�=��=$�=���=>!�=�zv="�^=4�J=�=;=.V/=n'=�i"=N� =.z"=x�%=�S)=�(=��=��=���<��9:����\����}���`�7r�����D�v*7�`Z�z?y��S֐�y���Qؐ�	툿�#y���Y��6�br�[;߾�)����S�3���N�`@;ƃ/=D��=��=l�=�=�   �   ^��=l�=E��=2�=�\�=)ߎ=��w=@U=��7=��=|=�=t��<�v�<���<�=�=:�=,�#=z)=L�$=��=���<M�;��ż������ �P��陾xeԾa�
�r-��QN�Bl������N���틿[Y���ρ�`l��BN���,��D
��BҾsH��iE�����e3��l�;�d8=#Փ=�'�=�n�=�{�=�   �   ���=>^�=q�=�ǒ=��t=V�C=�=���<�̕<�M<��<xl<8<�.?<H��<$��<��<V�=��=��&=_+=��=�
�<H�U<Иe���[���ݽ��7�ځ��BQ��6j���4�(�;��YW��m��{�����;{��Zm���W��)<��L�������Y󆾼�.�Ed���l	���Z<�VE=>�=�z�=�+�=���=�   �   c�=
�=�=�sB=N3=�<@g�:3;�Ҫ���ڼ�켨ἴ���Z����컀�-;�S<x�<��=(�=�#0=��.=��=4i�<�*��3�QS��]��ui�<���*%ھ�%	��$�m=�y�P�0]�քa�n[]�PQ�X�=��/%���	�x�ھ����aYg���V��좪�$�<��S=��==�=Ĳ�=���=�   �   ~��=��[=��=�vx<��л����	@��ʀ�xJ���}4�����5�����^��� �샺��6˻��<p��<b�=��/=@�<=.\0=��=�RW<�X���6q��I�-�:�ٙ��������89
��n��I0��1;��?�/�;���0��[ ��O�Nl�鶾.`��`p<��G�R+]����8��<`2a=�V�=2��=$e�=�-�=�   �   z�@=���<���:��Լf�`������߽���D��B���W�~L��� ��m׽D����h�&��`�h�:<d��<��'=t|E=�aI=�*/=H��<�;c;�� �TĞ�X�	���N��鍾PK��*�ݾ&� ����@���J��r�������E,�������Z�V�����ۧ�<����;R�=��j=a��=(�="Β=��=�   �   �[�< Fջ�!"�	c��1(�l��>���Z�ǋm��}u�Nr�B�c�<-L��-�M�O�ͽ����
��(�����<HX=x�F=�]=�U=�#,=�A�<0@���4+������>��P��刾'ۨ�y�ž �ܾ܆�q#�Y�쾷߾�Xɾ�񟎾�3]�Cv��7ν��W�()P��@�<��.=��m=�}�=N�=b�m=Ъ0=�   �   �:
�hU8�-Y���0���>�:�p�����������������2}�����L	~�n�N�jj���۽	僽�1ܼ�;4��<�i?=��i=��t=0A`=B+=�0�<�
��H8�TQ���+�l}>��p�%
������̱�� ����y�����F~�T�N�6g��{۽�ჽ0)ܼ�(�;��<>i?=��i=��t=�<`=\�*=� �<�   �   @+�ұ��6C��P��舾�ި�l�žS�ܾ+�뾶'�j��r߾�[ɾ����;���n7]��x�X;ν� X�5P��=�<��.=�m=�~�=�O�=��m=��0=�l�<��Ի4"��Z�����:�>���Z�P�m��wu�1r���c�D(L�ή-���
��ͽ�����
���$��<�X=n�F=D]=�U=,=�4�<p����   �   Uʞ�0�	���N��썾�N��	�ݾE� �3������L��t����` �8/ᾂ!��v���(�V����@ާ����� �;�=��j=[��=�)�=NВ=4�=̹@=���<��:t�Լ��`������߽��������R��G��� ��f׽�>���h������`	;<t��<`�'=�zE=�^I=�&/=���<��b;2� ��   �   P� �:�P�������H�2;
�q��K0�'4;��?�T�;���0�X] �>Q��n��궾�a��Jr<�:J�l.]���㻄��<3a=]W�=v��=�f�=,0�=t��=�[=��=h�x<�лD����?���_B��夽�,��������X�^�� ��v���˻�<���<��=��/=d�<=<Y0=x�=�<W<dg��F@q��   �   `�dyi�����(ھ{'	��$�w=���P�W]��a�d]]�Q��=��0%���	��ھз�� [g�)�����X�����<��S=��=+>�=)��=v��=��=��= �=
|B=�<=ী<�ш:X;�й����ڼX���j�p����J��P�� $.;��S<T�<��=�=�"0=v�.=��= a�<�ן�F:�X���   �   ��7�����pS���l��6���;��[W�`m��{����m={�V\m��W��*<��M��������l�.��d��*m	���Z<DWE=��=�{�=�,�=X��=���=d`�= �=�ʒ=^�t=ޥC=2 =x��<�ݕ<X*M<8�<0�<`0< D?<���<4��<��<P�=��=H�&=�]+=��=��<��U<جe�(�[���ݽ�   �   Y�P�t뙾EgԾp�
��-�SN��l����O��h�Y��wЁ�+l�sCN�&�,�%E
�3CҾ�H��6iE����pe3��r�;�e8=�Փ=p(�=do�=�|�=���=���=���=.�=_�=��=�w=vEU= �7=��=�=r�=��<�|�<h��<��=�=��=��#=� )=��$=Һ=���<�2�;@�żp���Ռ��   �   ��`�Qs����>E�H+7�?Z�Z@y�J�֐�Α���ؐ�<툿#$y���Y��6�Zr�3;߾�)��:�S�;2��b�N��(@;�/=ⴒ=���=�=��=K�=��=:��=x:�=)��=]%�=�=�"�=�}v=��^=xK=t?;=�W/=�'=�j"=�� =Pz"=N�%=pS)=>�(=��=�=���<��8:8�������~��   �   nlf����8��k,�@�:��)^�b�}�9g���m��_2��Gl��"_��5�}���]��:�D�
�� ���1�X�@<���X����:�^,=�>�=Ƈ�=���=ʂ�=���=d��=��=���=E`�=CƱ=�=��=!��=�-s=�^=ЙM=��?="75=��-=��)="�(=��)=�*=�(=�=�,=�_�< :�y�����(���   �   /�`�br����ᾂD�e*7�9Z�3?y��֐�$����א��숿#y���Y��6��q�:߾�(����S�A0��~�N��I@;��/=l��=��=R�=�=8K�=�=V��=�:�=H��=z%�=��=�"�=�}v=�^=K=$@;=�X/=� '=�k"=�� =�{"=��%=�T)=��(=�=��=L��<�|9:����ހ���}��   �   ��P��陾eԾ	�
��-�QN�sl�`���[N��%틿�X��Iρ�l��AN�~�,��C
��@Ҿ�F���fE�%���_3����;�h8=�֓=.)�=�o�=}�=���=��=8��=`�=9_�=��=��w=FU=��7=��=�=��=��<,��<`��<�=b�=�=��#=t)=��$=�=p��< S�;X�żJ���Ɋ��   �   ��7�,���PP���h���3��;�}XW�m�{����9{�Ym��W��'<�OK�G���������.��_��xe	���Z<@[E=:�=�|�=�-�=��=(��=�`�=J�=�ʒ=��t=l�C=� =��<tߕ<�.M<ض< �<�8<�M?<À<,��<H!�<��=`�="�&=�a+=� =\�<��U<H�e�Z�[��ݽ�   �   �[��si���q#ھ�$	�ʎ$��=���P�8]���a�HY]�. Q�L�=��-%���	���ھ-���^Ug����=������8�<f�S=@�=b?�=��=��=4�=V �=ƕ=�|B=N==<��<@�:��:�������ڼ���fἤ���E�����@].;x�S<���<�=��=�'0=��.=`�=�n�<�˞��/�+Q���   �   dF�מ:�P�������P徹7
�m��G0��/;�`?���;���0�uY ��M��h�
涾�]��,l<��@罌 ]�P��X��<`8a=EY�=֯�=�g�=�0�=���=�[=N�=h�x<`�лг�.�?�C��A��P䤽�+����������R�^��� �,o�� �ʻ��<$��<��=@�/=2�<=�_0=�=�aW<P��T1q��   �   r�����	���N��獾�H���ݾY� ������aH�?p����x��J(ᾑ����E�V�t���ԧ�^�� T�;��=�j=W��=
+�=Nђ=��=�@=���<�.�: �ԼD�`������߽���ȥ�Ĕ��R�rG�� �Te׽�<��,�h����8���;<���<��'=�E=�eI=�./=���<`�c;�� ��   �   -+������;��{P�8㈾*ب��žG�ܾ�������h߾�Tɾ3������� .]�tq��/ν��W�h�O�R�<�.=|�m=���=EQ�=|�m=�0=(o�<��Իf"��Z��n����>�Y�Z��m�0wu�� r�-�c��'L��-��
�!�ͽ����8
� 读���<�]=.�F=�#]=U=\(,=�K�<���   �   8�	� ?8�IK���'��x>�p�p�뎾���:���⭱���� v��&����}�\�N�b�s۽Jڃ��ܼ�y�;���<�p?=��i=�t=�C`=+=D3�<�
��G8��P���+�H}>���p�
����������۹���y������~���N�lf�%z۽�߃�� ܼPL�;x��<�n?= �i=��t=�E`=@+=�<�<�   �   �z�<p�Ի^	"�PT����X
�Һ>���Z��~m��pu�m�q��c��!L� �-���
�؃ͽ����R�	�𳯻쳕<�`=��F=�#]=U= &,=�D�< 7���3+�Z����>��P��刾ۨ�k�ž�ܾʆ�\#�>�쾒߾zXɾ��������.3]��u��5ν�W��P� I�<P�.=6�m=ŀ�=�Q�=$�m=.�0=�   �   ؿ@=���<�<�:�yԼj�`�����޽���������\M�zB�~� �$]׽�5����h�l�����0;<l��<��'=��E=LeI=J-/=���<�Pc;�� ��Þ�4�	���N��鍾CK���ݾ!� ����<���J��r������,����T�����V���ڧ�����)�;\�=\�j=&��=y+�=cҒ=$�=�   �   �=Z�[=*�=`�x<p7л��ἔ�?�ͺ���9��/ܤ��#��@���������^��~ �P]����ʻ8�<���<�=|�/=��<=0_0=��=�XW<�V���5q��I��:�͙��������69
��n��I0��1;��?�-�;���0��[ ��O�)l��趾�_���o<��F罼(]�p�����<.6a=�X�=��=�h�=D2�=�   �   ��=b"�=�=H�B=:E=���<�4�:��:�������ڼ�v��O�d���,2�� S���.;�S<P��<��=$�=r(0=Į.=��=xl�<@��R2�
S���\�tui�3���!%ھ�%	��$�l=�y�P�2]�؄a�p[]�PQ�V�=��/%���	�V�ھ}���Yg����W������4
�<��S=��=\?�=���=��=�   �   /��=(b�=,�=8͒=��t=��C=2=	�<\�<pQM< �<ذ<�V<xh?<X΀<���<�(�<��=:�=B�&=Zb+==��< �U<��e��[�E�ݽ��7�с��=Q��1j���4�(�;��YW��m��{�����;{��Zm���W�})<��L�������8�r�.��c�� k	�8�Z<�XE=��=�|�=�-�=���=�   �   t��=���=b��=��=�`�=��=<�w=,KU=�7=8 =��=�=���< ��<���<��=��=�=�#=H)=X�$=4�=���<@S�;��żr�������P��陾teԾ`�
�s-��QN�Bl������N���틿\Y���ρ�al��BN���,��D
��BҾ`H���hE�����d3�v�;&f8=�Փ=�(�=�o�=T}�=�   �   RK�=`�=ʂ�=2;�=��=l&�=+��=�#�=��v=ض^=�K=�B;=$[/= #'=�m"=�� =}"=��%=�U)=v�(=¨=X�=���< �9:���A����}���`�6r�����D�t*7�`Z�z?y��T֐�z���Qؐ�	툿�#y���Y��6�br�S;߾�)����S��2����N�@@;r�/=���=���=�=��=�   �   r�=pv�=�	�=z�=@��=5n�=��=fdu=ڃ^=�aN=�(E=��B= �E=zN=:�Y=�g=.Pu=K�=�ł=�8=�6g=�s5=t�<�Q��3h�|���/�Z��è�r�F�#��S��ꁿd���,��퍾�!ɿI�̿Tɿ�{��������Ņ��#R��"�k�P��6�N�(?ݽ�x�'�<�Z=���=~H�=xa�=�   �   3�=���=��=7	�=�ߠ=;F�=؂y=![=�>C=��2=`]*=&6)=t�.=9=`H=�?Y=t2j=�xx=��=Fo|=��f=i7=���<`s��]�WM���6U�����>�� ��3O��3�����/���P����ſ>?ɿϫſ"H��N��n}��(�~��KN�"����kޠ���I���ֽ���,Ӌ<��\=�@�=���=�k�=�   �   ^I�=�ܽ=I��=�`�=�=~{X= v.=@�
=pl�<���<di�<��<�]�<���<��=b�-= H=�g_=�o=j�s=�e=��<=���<����?�+c߽�E�����~$߾����C���q���s���籿cͻ��<��$ۻ�^�������eݎ��\q�`SC�Y��u�ܾNޖ���;�xaýp�꼨q�<�a=S=�S�=�g�=�   �   �>�=`ޠ=Sk�=��Z=��=|�<p:3< Xָ@��@�M� vZ���-�PT�� �\;8�W<t��<�]=U3=��Q=�b=>`=�&C=�
=���;����7����-�����-ɾ�	�_2���\��ɂ��政�.���]������H|���^�����傿L�\��&2�x		�SmǾ�H��pt%�k���Þ�x��< h=���=��=}�=�   �   �W�=��m=�)=���<�W;pa��#��N�F�w�~3��xd���t��(K� ����@�z��2N<�[�<>A$=J�G=8�U=�HH=B=��q<H����m�dyj�yc��}6���A���f�����i��%���`���ܘ�(���Y惿�0g��bB��L�v2�ɯ��J,g�s�	�h�x� �'=��m=,і=��=�1�=�   �   jRM=,K�<�S�;ܑ����B��>��L�˽�(��{�������.=����|�������)+�\�٨;T��<H�=<�B=DI=h,=`�<P���b�B�z`ڽ��;�$��e�ƾ����#�usC�,�_�L-v��P���ᄿ�����v�t�`��mD�/�$�ޢ�g�Ǿ���0
;�b�Խ��+��&�;<5=�p=E��=V<�=���=�   �   P��<05�����J�����ֆ�#�:�(xV�Q�h��<p��8l��T]�t E���%�������g�pOɼ��F;�U�<�8$=.�B=��<=s=HJH<����G����
���[����zѾE#�c��k�6�%�I�u�U�O'Z�q@V��nJ���7�4* �W���/Ծ{��k�_���$Ŕ����ോ<L)0=T�l=��=��l=^i6=�   �   ����=�V̹��L���C��uw�Cܒ��]��f����0������5;������6��$Q����gٽ��~�\�ż@��;4y�<:�2=�F=�2=8@�<�Dl:x��,��ҥ���h��Ş�˾C��l}������'�]�+��n(�������<�����ξ?Ԣ�Y�p�X8$�'<Ľ�_/�@�ѺT��<�@=��a=T�Z=Z+=���<�   �   �>�	JŽ�X���`�,풾|Ǵ��,Ӿm뾪?���� ��y��l���־�1�������k�|	*�R�ܽ �j��n����}<�=��G=�UN=x+=l]�<�ܻ6�>��AŽ]S���`�l钾5ô��'Ӿuh�y:��� ��t������־..���	����k��*�:�ܽ�j�(f����}<B =V�G=�RN=|�*=$O�<@�ܻ�   �   F3�������h�Hɞ�V˾�G���������'�>�+�Vq(�O���������ξ�֢�7�p�*;$�
@Ľ�d/���Ѻ��<�@=�a=~�Z=$`+=�
�<���b�=�ù�0G�b�C�Mnw�Gؒ�qY�����f,��T�S7��b���3��4Q����aٽ��~���ż �;x|�<�2=B�F=,2=�4�< Cj:h���   �   ��
��[�����}Ѿ�%����C�6�(�I���U�W*Z�UCV��qJ�/�7�9, ���`2Ծ}��V�_����ǔ�������<�)0=<�l=<�=��l=hp6=���<������"B��`�������:�IqV�:�h��5p�(2l��N]��E���%�������V�g�tAɼ`EG;T[�<�9$=r�B=��<=�n=�1H<�����M���   �   ��;��&����ƾ���k�#�vC�	�_�N0v�"R��%ㄿr�����v���`��oD�ˎ$�"��M�Ǿk���;�оԽ��+��;~5=p=���=i>�=���=�YM=�]�< ��;Dv����B��5��E�˽	��������D��N8���㽚t�������+�X�����;@�<�=~�B=I=Le,=|�<P���n�B��fڽ�   �   g}j�f���9���U�A�#�f�k���-k����������Mݘ�T���`烿x2g��cB�N�4�񰬾�-g�l�	�.j��� �^'=�m=SҖ=T�=�3�=�Z�=�n=�)=���<�	;�E����N���w�\+���\��Lt��K��	�x��� �z��HN<Lc�<�C$=H�G=�U=�FH=X=��q<@���E����p��   �   j���/ɾa�	��`2���\��ʂ��甿+0���^��Ɣ��Y}���_������傿Z�\�w'2�
	�nǾ I��u%��k���Þ����<Hh=���=C	�=1�=�@�=�=�n�=h�Z=��=���<�d3< 쿸8��ЌM�xJZ���-�P��`];�X<|��<Na=rW3=�Q=P�b=h=`=�$C=�=�f�;���;����-��   �   -���{&߾(��_�C�M�q���Z����豿Fλ��=���ۻ��������ݎ�O]q��SC����čܾsޖ�
�;�Iaý��꼸s�<0�a= ß=�T�=�h�=�J�=c޽=x­=-c�=��=ށX=�|.=p�
=�z�<���<w�<(�<�h�<h��<��=Z�-=>	H=�h_=��o=4�s=�e=�<=\��<`���!?��f߽j�E��   �   ��"@�d� ��4O�	5�����40��tQ���ſ�?ɿ)�ſcH��{���}��4�~��KN���N�!ޠ�*�I���ֽ ��l֋<�\=�A�=p��=�l�=�3�=���=	�=�
�=8�=�G�=R�y=�$[=BC=@�2=�`*=�8)=�.=9=�aH=�@Y=3j=yx=��=�n|=��f=�g7=0��<���:�]�%P���8U��   �   <Ĩ�Q���#�wS��ꁿ�d��*-�����4ɿH�̿?ɿu{�����{�������R���"�����O���N�C=ݽ�u��+�<��Z=2��=
I�=�a�=dr�=�v�=
�=�z�=��=bn�=��=�du=��^=�aN=X(E=F�B=��E=�N=��Y=\�g=tOu=�J�=ł=�7=�5g=�r5=��<�Z��6h�Y���`�Z��   �   #���>�� ��3O��3�󷖿t/���P��5�ſ�>ɿN�ſ�G������|���~��JN�D���:ݠ�ڶI���ֽz��ڋ<Z�\=B�=Õ�=m�=,4�=���=$	�=�
�=R�=�G�=~�y=�$[=NBC=��2=�`*=n9)=l�.=d�9=XbH=�AY=�3j=�yx=%�=�o|=��f=�h7=���<�z�H�]�#N��@7U��   �   g���!$߾�����C��q�[��~��Y籿�̻�<��Aڻ�v��������܎�[q��QC�&��w�ܾ�ܖ���;��]ý����z�<��a=�ß=�U�=Li�=6K�=�޽=�­=[c�=�=8�X=,}.=��
=�{�<���<`x�<�)�<�j�<���<�=څ-=�
H=�j_=V�o=P�s=(e=��<=��<���<?��b߽��E��   �   ����,ɾK�	�9^2���\��Ȃ��唿.���\��{���{���]�����䂿O�\��$2�	��jǾ�F���q%��f���������<�h=���=
�=��=TA�=l�=�n�=��Z=0�=t��<�f3< ��������M��FZ�(�-�����*]; X<���<�c=�Y3=��Q=B�b=�@`=�(C=�=���;��t6���-��   �   �wj�2b���4�����A�ܓf�����h��ܭ������ژ�³��僿<.g�I`B�K�4/�(���'(g�>�	�&^�@q �h-=�m=�Ӗ=\�=�4�=[�=�n=��)=���<�#	;�D��x�8N�0�w��*��!\���t�0K��,����bz�PSN< i�<�F$=��G=ֺU=�KH=�	=�r<(ꧼ��l��   �   \�;��"��X�ƾ���k�#�uqC���_��*v�.O��'��������v���`�kD�Ԋ$�֠��ǾR����;���Խ��+�@i�;$<=� p=R��=�?�=U��=[M=�_�< ��;�t����B�H5����˽������d������7��㽙s��U���$+��ڍ�`�; 	�<� =ĚB=	I=�k,=P�<�m��v�B�3]ڽ�   �   2�
���[�g��<wѾ�!�R���6�x�I���U�E$Z�[=V��kJ���7��' ����+Ծ�w���_�ͦ���������ǋ<�00=�l=��=�l=r6=��<@��ʮ��A����܀���:� qV��h�r5p��1l�YN]�kE�V�%����g�����g�4;ɼ |G;�b�<�=$=��B=��<=
w=p\H<����JD���   �   '�������h����˾?��{�0���'�v�+��k(���� ��I���p�ξ�Т�)�p�T3$�'4Ľ S/� Tк\��<~@=��a=Z=fb+=��< ����=�$ù�G�@�C�+nw�7ؒ�_Y���N,��6�-7��1���3���Q�@�J`ٽ�~���ż`5�;���<�2=j�F=2=�I�< �m:���   �   ��>��;ŽoO���`�`撾�����#Ӿ�c�u5��O� ��o�����Ϣ־�)�����I�k�m *��ܽF�j�`N��x&~<�(=��G=ZN=x+=�a�<p�ܻ4�>�\AŽ4S���`�]钾(ô��'Ӿih�l:��� ��t������־�-��o	��p�k�g*��ܽ�j��_���~<�$=�G=ZN=:+=�h�<�Tܻ�   �   �����=������B��C�hw��Ԓ�pU���}���'�����2��>��0���Q����Wٽڋ~�L�żn�;h��<�2=��F=�2=�E�< �l:8���+�������h��Ş�
˾�B��i}������'�W�+��n(������������ξԢ���p��7$��:Ľ]/��0Ѻ|��<@=D�a=�Z=ne+=��<�   �   `��<��ȣ��:������{���:��jV�/�h�T.p��*l��G]�E���%����}���g�(&ɼ��G;Tn�<�A$=��B=��<=Dv=SH<���iG��t�
�Ս[�����yѾ@#�_��i�6�#�I�u�U�M'Z�o@V��nJ���7�(* �G���/Ծ�z����_�����Ô���ؼ�<�-0=�l=L�=Z�l=0v6=�   �   �_M=Tm�<���;�^��x�B�[-���w˽���p�����z���2�2�㽿j������6+��ō�_�;L�<>=��B=�
I=�k,=��<@��<�B�`ڽr�;�$��X�ƾ����#�rsC�*�_�L-v��P���ᄿ�����v�q�`��mD�&�$�Т�C�Ǿᯎ��	;�s�Խ��+�P=�;�8=0p=d��=d@�=�=�   �   �\�=�	n=b�)=�Ŷ<@�	;�,����<�M�:�w��"���S��4 t��K����$��� �y��rN<du�<TK$=�G=��U=�LH=6
=�q<��]��m�Lyj�oc��t6����A���f�����i��'���a���ܘ�*���Z惿�0g��bB��L�^2ﾬ���,g��	�\f��� ��)=P�m=�Ӗ=��=�5�=�   �   �B�=6�=Eq�=��Z=z�=���<��3< ����_�X[M�xZ���-�@���@�];�>X<l��<6i=V^3=�Q=��b=BB`=�)C=�=��; ��T7����-�����-ɾ�	�_2���\��ɂ��政�.���]������K|���^�����傿J�\��&2�r		�?mǾ�H��1t%�yj��x������<�h=R��=R
�=��=�   �   �K�=�߽='ĭ=8e�=X�=��X=L�.=��
=H��<Ƞ�< ��< 8�<\x�<���<v�=f�-=�H=�m_=o=�s=te=��<=t��<����?��b߽��E�����y$߾����C���q���r�� 豿eͻ��<��%ۻ�a�������gݎ��\q�_SC�W��j�ܾ?ޖ�Ҋ;�aý|��Tt�<��a=zß=nU�=�i�=�   �   T4�=&��=�	�=x�=Q�=2I�=`�y= ([=�EC=>�2=�d*==)=�.=��9=PeH=
DY=,6j=�{x=��=q|=�f=j7=��<�oﻺ�]�@M���6U�����>�� ��3O��3�����/���P����ſ??ɿЫſ"H��Q��o}��'�~��KN�!����bޠ���I�V�ֽp��dԋ<p�\=aA�=r��=�l�=�   �   \s�=̄�=6�=i�=o��=`Pw=|�R=^Q4=��=P�=�=f�=�(=��?=�Z=w=_��=㚒=ѹ�=�Α=��=�*8=�'�<���zh;��J���m�K�%��i]����&��1�ɿNH�A/��Y�@���T����e �Brɿ|����W��Q�[�H�#�4�����v1����(�p�&=jy�=┫=1g�=�   �   �J�=e��=l8�=F�=fV�=�K[=t�3=��=�m�<<��<P<�<�N�<b�
=��$=~bC=�c=�ˀ=B��=�t�=�)�= �}=R9=̤�<��ۼ���ݧ6������徥h"�l_Y�H����3����ƿ�x����U(��v��(������E��"ƿ�������X�W�� ��&�3֓�5-�0j��p1V�L�=��=��=�޼=�   �   ��=�å=��=��q=�;=:�=D1�<��2< '�;��I: �}:�`�;X�5<4>�<T5�<�'=�yQ=h_t=S�=X��=&pv=#;=DY�<,ŭ�,:��N�(�������׾�=���M�b������:����jտ 鿉���b��g�����#mտ9���Q���킿E�L�h���ԾNt���F �;�ؔ
�p>=ȁ=��=��=�   �   ���=)�=v|I=T=�h<`�l������R�TJ)���9��G5��r�pI�p{� �|�h<�@�<�4=��\=��p=��h=�{<=(~�<��O�����q��}�¾P�
�iO;�W-p�\6��	3���'Ŀ7Dֿ���S��"�)�ֿlĿBX���1��)�o�!�:��
�Qj��̜w��S��n�@�ºf=dz}=R=l�=�   �   �_=�4=@��<`�||���i�����7ǽ�߽�����+ҽ���5Ȋ�ܒ9�L�� �K:�Z�<��=�D=��Q=L?:=d�<���r�K�_��*V�����V���$��fS����H|��A*���u����ȿ��̿�;ɿ^龿��癿�Z��g�S�w�#���	Q���}R�?��/�0k�;܌#=��q=}Q�=E�=�   �   0��< K�;��ּ�v��,Ľ8���%�;.?�dP���V�ږR��AD�,%-�|w���۽yᕽ��$�p6+�p�j<b;=��.=lM1=�=P�<����7P��]t*��"����Ⱦ��	�Q�2��9]����.#���f��올��᯿묿�󣿢ʕ������C^�g�3��5
�$Zɾ$�Z�(��孽زѼ��<�*=�^=@Xb=��==�   �   �h���&"�,˧�>0�%�6�Kh�v:���������������ƨ��U��ʳ����p�xA�_��HϿ���R��ڀ�x�D<�5�<:�=|u=XU�<h4�"<l�x���S�ݞ���ܾW��{4�QW�ӫu��󆿆ǎ��������싇�`)w��X���5��	��޾O>��0U�՜��jlh�h
�Ь�<8o+=�@=�$=�Y�<�   �   ��6�\�����;\��i��o�
оU辚���i��������_��TӾ���������e��s$�bҽ��Z���f��k<\| =��=#�<@��;�鼩<��f���l������߾���(���A��U��b�bg��\c�~W�]~C�*�kr����������p�R�� ⨽�������;\�<��#=:A=x��<�	Ȼ�   �   C����<!��Fo��R<о*l��* ���!���+�s�/�h�,���"���� �Q<Ծ��8�v�2a(��Sʽ�~;������<�=p�=�ٿ< (���%�����7!��?o��q7о�f������!�Z�+��/�-�,���"�B��@ �w8Ծ��}�v��](��Nʽ,x;��������<��=}=ο< @��.�%��   �   ���l����=�߾���=�(�6�A���U�>�b��eg�X`c��W�Q�C�O�*��t��⾃���\�p� ���娽������;p�<>�#=F=P��<`�ǻ��6�S��O��!4\��e���뱾�о�	�ڵ������+����Z�1PӾ������q�e��o$�[yҽ0�Z�0�f��k<�| =�=��<0u�;�.鼎C���   �   (�S�U���� ݾ���t�4��W�}�u�����}Ɏ�홑��������l,w���X���5�m���޾E@���2U�n����ph��
� ��<@q+=�!@=D�$= k�<����"������*���6��h�B6��-�J���	���¨��Q�������p�	A����ȿ���R�̀�x�D<�9�<��=s=�K�<��4��Fl������   �   �%��ɾ��	���2��<]����%��{h��ۚ���㯿�쬿����̕�Ů���E^��3�%7
��[ɾl��(��筽l�Ѽ`�<��*=�^=*]b=��==���< ��;��ּRyv��"ĽT��n�%�F'?�.P�\�V��R�;D�^-�tr���۽�ڕ�>�$��+�h�j<h>=�.=�L1=(�=ظ<����U��Ix*��   �   2�������	$�iS�,���}���+��`w��z�ȿW�̿}=ɿ�꾿<����虿�[��ҡS���#��R��R��@�0/� l�;4�#=n�q=rS�=�=�!_=�==��< �� m�D�i�􄢽�ǽc{߽��齚�位!ҽ4������V�9��7�� �M:Pf�<R�=~!D=4�Q=�=:=�]�<�L�^�K����.V��   �   *�¾��
�NQ;��/p��7��q4��q)Ŀ�EֿW����J$�]�ֿ�mĿY��/2��1�o��:�X 
�k����w�`T�x�n���ºRg=�|}=�Ø=,n�=*��=x�=��I=�=�/h<��k�Ц��pD��;)�6~9��95��e��1鼀F{� Ft�`<8K�<��4=��\=~�p=d�h=Lz<=�w�< �O�o����s��"}��   �   ��׾A?�1�M��b������T����kտ8鿭���s��Z������mտ����Q��4��L����K�Ծ[t���F ���8�
��?=�ȁ=M��=Z�=ؖ�=	ƥ=F�=��q=J�;=B�=�B�<��2<�q�; <L:@�:���;�	6< K�<�?�<N�'=�|Q=�at=�S�=v��=Zov=B!;=S�<lέ�q=����(�|����   �   %�徛i"��`Y�홊��4��`�ƿWy�}���(��v��(������E�#ƿ����
���6�W��� �h&��Փ��-�i���)V���=��=���=�߼=�K�=���=�9�=��=GX�=�O[=ȥ3=r�=�v�<��<�D�<V�<��
=F�$=�dC=��c=.̀=���=�t�=g)�=ޔ}=�9=h��<4�ۼò����6�Pᗾ�   �   �n�ޑ%�Kj]���m&��~�ɿ�H�p/��Y�@���T����$ ��qɿ&���yW����[���#�@��T���u1���� �p�D=:z�=���=�g�=�s�=3��=��=Xi�=���=�Pw=ҦR=�Q4=
�=4�=��=��=��(=��?=P�Z=Nw=���=r��=N��=(Α=z�=<)8=d#�<������i;��K���   �   ���h"��_Y�L����3����ƿbx�p��(�jv�P(������D�E"ƿꨨ�n8�W�#� �<%��ԓ�`-�jg��� V���=:�=^��=�߼=�K�=֧�=:�=�=]X�=�O[=�3=��=w�<���<E�<�V�<�
=��$=4eC=<�c=ỳ=蘌=u�=�)�=�}= 9=(��<(�ۼ����f�6�n����   �   s�׾�=�>�M��a��-��������iտ;�迗���T��G������kտ#~���P��	킿��L�!���Ծ�r��@D ��퐽�~
��B=�Ɂ=��=��=2��=Lƥ=|�=R�q=��;=��=,C�<��2< u�; WL:@(�: ��;�6<�L�<�A�<^�'=�}Q=�bt=qT�=S�=zqv=�#;=Z�<�ĭ�:��2�(������   �   ��¾��
��N;�@,p��5��+2���&ĿCֿw����m!⿥�ֿkĿ�V��?0����o�>�:�H
��g���w�.Q���n������k=n}=�Ę=�n�=���=��=�I=X =�1h< �k���� D�
;)��}9�95��d��/��A{� �r�$<dN�<��4=��\=�p=N�h=~<=���<�O�����\p��}��   �   o������$�eS����*{���(��t���ȿ۬̿:ɿ�羿:���4晿�Y���S�_�#�,�eN���yR��8�n/����;^�#=��q=�T�=��=�"_=�>=��<���~l���i������ǽ#{߽���7��!ҽ������Ԅ9��4���fN:�j�<��=\$D=��Q=vB:=�i�<����K� ��)V��   �   r!����ȾF�	���2�a7]��
���!���d������߯�鬿���ȕ�ҫ���@^�Ȉ3��3
��Vɾm1�(��߭���Ѽ� �<V�*=�^=�_b=X�== ��<���;�ּ�xv�["Ľ5��R�%�%'?�P�2�V���R��:D�-�r�Ƥ۽�ٕ�2�$��+��j<�A=��.=�Q1=��=X�<����LM��Yr*��   �   |S��ڞ���ܾ���B}4���V�Ĩu��񆿭Ŏ������������%w���X���5����޾�:���*U������_h���	���<w+=�%@=��$=�n�<����"�����}*�a�6��h�46���:������������Q��母�-�p��A�����ǿ�v�R��ǀ� �D<�A�<�=�y=@^�<pS4��5l�����   �   S��bl����߾Ƴ���(���A���U��b�Y^g�Yc�� W��zC���*��o������0�p�X��?ڨ�l����'�;�"�<�#=�I=���<@�ǻ��6��R��"���3\��e���뱾�о�	�̵���������pZ�PӾ�������e�ho$�Ixҽ��Z� �f��k<�� =��=�,�<���;0�8���   �   B����3!��:o��뢾}3о�a��`����!��+���/�Œ,�=�"� ��e �r3ԾX즾p�v�X(��Eʽ�i;�0����<��=��=��<���h�%�����N7!��?o��c7о�f������!�U�+��/�&�,���"�6��0 �P8Ծp��v�<](��Mʽ|u;�������<��=N�=��<@R�@�%��   �   N�6�IL�����.\�@b���籾: о��E����|��S����T��JӾ�򵾆'�e��i$��oҽd�Z�@�f���k<� =��=@,�<���;���;��,��\l����~�߾���(���A��U�}�b�bg��\c�xW�T~C���*�\r���⾿���#�p�ܙ��਽�����;��<�#=@K=���<�vǻ�   �    ņ�:"�����&��6�h�p2���뛾����L�D���.M��������p�A�������D�R�0����E<tL�<T�=*{=0]�<�]4�z:l�����~S��ܞ���ܾS��x4�OW�ӫu��󆿅ǎ��������싇�[)w�	�X�~�5��	���޾*>���/U�����ih� �	�ܵ�<xu+=B&@=��$=�x�<�   �   8��<��;�sּ�jv��Ľ��n�%�� ?� P���V��R��3D��-�>l���۽*ѕ��$��*�(	k<�G=�.=T1=��=�<�����O��)t*��"����Ⱦ��	�N�2��9]����.#���f��혬��᯿묿�󣿢ʕ������C^�^�3��5
�Zɾ ���(��䭽��Ѽ��<:�*=�^=�ab=<�==�   �   �'_=E=� �<�I�h_�n�i��{���	ǽ�p߽��齌���ҽ���[����u9���� Q:p{�<<�=()D=��Q=hD:=@k�< ����K����*V�����M��$��fS����I|��B*���u����ȿ��̿�;ɿa龿郞��癿�Z��c�S�p�#�{��P��|}R�\>��/����;֐#=X�q=2U�=9�=�   �   ,��=�=�I=�'=�Vh< +k�d���x6��,)��n9� *5�TV�|鼐{� (h�(I<�]�<��4=��\=~�p=�h=�<=<��<��O�&����p��}���¾M�
�gO;�U-p�\6��
3���'Ŀ8Dֿ���V��"�,�ֿ�lĿBX���1��&�o��:��
�?j����w��S���n��Uº�h=b~}=Ř=�o�=�   �   ��=�ǥ=T�= r=X�;=Z�=�R�<�2<н�; �N: X�:`�;�/6<�\�<�O�<|�'=��Q=gt=V�=��=�sv=p%;=�\�< í��9��2�(�������׾�=���M�b������:����jտ 鿌���e��k�����&mտ:���Q���킿B�L�c���Ծ=t��tF ���h�
�N@=UɁ=荣=4�=�   �   L�=J��=�:�=�=�Y�=�R[=��3=��=��<Я�<�N�<8`�<|�
=�$= iC=��c=�̀=#��=.v�=�*�=��}=�9=d��<��ۼ򯸽Χ6������徤h"�l_Y�I����3����ƿ�x����V(��v��(������E��"ƿ�������V�W�� ��&�+֓�-��i���.V�,�=s�=���=�߼=�   �   �Ȳ=�Ӭ=��=w�=Roc=t�4=�
=d8�<,%�<��<�f�<��<���<Tb=l3?=��g=6w�="6�=�ϙ=�J�=��w=,�= ��9�@h�����	����о@���W�����m'���\ڿm&��8��s��;&��N)��5&��[���co���hٿ#������w�U�<��I;��|����n�F�x�<ܬD=��=�=�   �   ���=��=K�=d�x=�wE=��=`�<�~<XG<P��;�;�pC<��<���<ڤ!=O=�x=�]�=��=㐏=�t=�1=���:2�^�y�
�$~�My̾���b�S�P$��j����ֿ������h��6^#��b&��_#�Һ�R���U����տ���R����Q�;����Ⱦ,w��?��~>���(<hD=t�=�u�=�   �   Tי=�r�=�f=��*=�g�< �%< ����{�T����ռ��ɼ|x��h� �O;|�<8�=��:=>�h=[��=��=��h=�>=l�;n�C�������l�# ��V�z=H�&ل�W,��R%̿���ظ���D(�B��;�(�h���l�۪˿w������6�F�Ǉ�������f�*q��;&��QP<ZvA=�d�=K��=�   �   �s=v�@=�@�<�v<�U�Ȟ���\�����䢽�=��wq��I����q�)�h/�� $��`@�<��=�cH=��_=܀S=`=�t<����۽UAR�^�������L6���r�6��S���.�ۿ�����<�����6�0���x�R��m�ۿk�����.r��M5��� ��O���UM�}�нn��Ѓ<I;=��y=>{�=�   �   d�=���<P���$!����E�ν��<����(�`B.�Li*�U}����uܽ�g����D����� ��;���<�#=(2=��=��]<"Ӽe���Ϯ0�9����و���U�c��&~��NCÿ��ܿ�������G�EN����tݿ��ÿe⦿H���d�U�y%�	�߾����A7-� 8���驼|z�<��.=J'S=z�G=�   �   ��;��м&��R�׽�L�7�E���m�ڲ�����	��+��ʚ���s�
yL�r!��b�3?���Z
�@M:�|ҟ<�I=�R=Ĩ�<��T�j����B��Vq����5���4�G;h�0r��¦���彿KqϿ$�ڿ��޿SIۿ�Hп7྿2���L(��l*i�P^5���ꃺ�%p��I	���v�@��\Y�<��=@�=(��<�   �   ��m���{��D�nӁ��䠾�˼��Ӿl������w3վ�����n������}L��9�C$�� �*�P:���w<���< ��<�md���!�e�ɽ��8��"��
�־2��q�=��Wj�c�������w�����L��������U��c��������'l��,?�����׾tǓ�^>9�)�Ƚ�J����:0޽<$"�<8�<@B���   �   �ﭽ����`�qq����ľl�E~
����m#�0
'��$�����&����{�Ⱦ�;���g��'⸽�)��ͻ�i<<;�< �<ԍ��ۏ���~�T�Y�F
���s⾯D�(�8�F�[��{�iމ�ݑ�%Ɣ�P��f���b}�>�]�/�:�~���徸�����\�O�e������L)<|ǰ<\͋<��%��a��   �   #����g��M��ܾ�
�$t&�E?�O�R��_�Vmd��`��eT��"A�F(���Ѻ߾�h����l���|-����� @a8,m�<(W�<�%�:H���5������g�OI���̢ܾ
��p&�9A?�4�R��_�$id��`��aT��A�X|(�m���߾�e��f�l���N)����� Xh8k�<|O�<@F�:x��������   �   (�Y���sx⾥G���8�2�[� {�����aߑ�sȔ�PR��s���}�q�]�ڡ:����:�/����\�RQ��g��T���hM)<lͰ<�؋<�b%�0U�_筽����`�m����ľy��z
�����i#��'�Z$�~���#����@�Ⱦ�8��Ig� ��ܸ�� )� �̻`i<�7�<0�< ���镀����   �   �%��:�־ԗ���=�a[j�x���X����y��*"������A����W��F���(����*l�/?������׾6ɓ��@9���ȽPM� ��:��<�+�<�<@���ț��c���u��D�@ρ��ߠ�NƼ��Ӿ������Y��'.վ�����j��$�����K��5�����*�p�Hx<��<ॢ< �e�� "��ɽC�8��   �   \���`����4��>h�t��ب���罿�sϿ��ڿ��޿�Kۿ�Jп⾿�����)��},i��_5�������.'p�K	�"�v�X���\�<��=&�=Ԡ�<�K�;�м��^�׽zF�ЩE�R�m�t������1���������p�r��rL�!�Z�l8��lP
�`�9�۟<�K=�Q=x��<��T�6 ��NF�n[q��   �   ������U��d�����GEÿ��ܿ������H�PP��ه�!vݿO�ÿ�㦿*�����U�r&�`�߾_���B8-�9���驼h}�<��.=�+S=��G=�=���<б�j!�jy��O�νp������(��;.��b*�Gw�x���kܽ�_���|D�����@	�;���<�#=�(2=t�=Ђ]<�.Ӽ9���P�0�����   �   ;���N6�&�r�f7��囻��ۿ����~=�����7���jy�`S��x�ۿ>���v��� r�RN5�*� �GP��]VM���н�~�pӃ<�K;=$�y=�}�=�s=p�@=8T�<��<�eU�h��"�\������ۢ�x4���h�������q��)��� ���lN�<��= gH=z�_=�S=�=�e<��#�۽�DR������   �   ��?H� ڄ�w-���&̿	����� )���L<��(�м��m�S�˿ˁ����x�F���������f��p�:&��XP<�xA=�e�=��=�ٙ=�u�=��f=��*=�y�<��%<p���pS{�y���hռ��ɼ�c�����@%P;�<��=�:=.�h=A��=��="�h=�<=PO�;��C�Ű����l����   �   �����S�%��5����ֿ����n������^#�c&�`#���t��V���տ���=����Q���F�Ⱦgw�,?��|>���(<xD=u�=�v�=⠬=���=�L�=t�x=J|E=��=�<�~<�]<p�; 5�;h�C< �<$��<��!=BO=��x=^�=�=���=Z
t=�/=�T�:��^� �
�P&~��z̾�   �   ۺ���W�����'��\]ڿ�&��b��s��;&��N)��5&��[����o���hٿ���1���U����P;�|�o���F���<ҮD=̹�=���=?ɲ=Ԭ=r��=��=pc=�4=\�
=�8�<d%�<Ԃ�<f�<��<���<�a=�2?=�g=�v�=�5�=Hϙ=AJ�=��w=&�= W�9Dh�ƃ��
����о�   �   6����S�b$��n����ֿ����ү�0���]#�Tb&�^_#�`��܈�U��#�տ.�������Q�E��5�Ⱦ�w�">��y>�p�(<�D=�u�=8w�=��=���=�L�=��x=t|E=̐=P�<p~<�^<��;�6�;h�C<��<���<�!=�O=�x=O^�=s�=#��=vt=T1=@��:��^��
��$~��y̾�   �   0�2=H��؄��+���$̿��l��r��'����:�P'�����k�˿\��������F��������f��l�N5&� gP<{A=�f�=���=�ٙ=�u�=�f=��*=z�<��%<p���pR{�xx��hռ��ɼ�b������.P;��<��=��:=*�h=ޒ�=��=,�h=�?=�n�;Z�C�������l�  ���   �   >��KL6���r�Y5��w����ۿ�����;�����5�<���w�IP����ۿߐ��u��r��K5�8� �sM��aRM�\�н|w��݃<�N;=t�y=v~�=s=8�@=TU�<@�<dU���ȴ\�����^ۢ�>4��<h�������q� )�,�� ���P�<&�=�hH=��_=��S=�=�{<�v�۽�@R������   �   J
�ԇ�{�U�b��}���Aÿ��ܿ��������E�L��у�mrݿ�ÿ�ি����ɬU�\#���߾�����3-�q2���ש����<�.=�.S=ҠG=6�=t��<@���!�.y���νX����ޒ(��;.��b*�w�C��zkܽ_��v{D�ܜ����;���<��#=\,2=&�=0�]<�Ӽl���t�0�>���   �   D������g�4�)9h��p��1����㽿AoϿ��ڿ3�޿�Fۿ}Fп�ݾ����m&��-'i��[5�{������p��E	���v����8j�<(�=2�=���<�V�;0�м����׽[F���E�9�m�f���x�����������8�r�VrL��!�ZY轤7���N
��9����<bO= W=̰�<��T�����A�	Tq��   �   � ��k�־p��5�=��Tj�����4���vu��z��읹�����ZS�����o���($l��)?�F����׾(ē�U99���Ƚ�>� ��:��<�4�< ��< ���j���c���u�lD�2ρ��ߠ�BƼ��Ӿw�����F��.վܼ��ej��������K�45������*����x<��<���<�*c���!�s�ɽ��8��   �   ��Y����+p�B�t�8��[�{�^܉��ڑ��Ô��M�����}�F�]���:�|��������^�\�NJ��]��y���t)<�ڰ<��<�2%�FS��歽ƻ��`�m����ľo��z
�����i#��'�Q$�t���#�����Ⱦf8���g�����۸���(���̻�1i<�E�<�	<(���Ƌ���{��   �   x��N�g�)F���ܾS�
��m&��=?�t�R�ظ_��dd��~`��]T��A��x(�F����߾Qa��`�l�B�� ��2�� ��8@�<|c�<���:����X��������g�@I���ܾȢ
��p&�8A?�2�R��_�!id���`��aT��A�J|(�]����߾�e���l�H�(��x�� �z88x�<0b�<@��:x���𩡽�   �   ᭽Ʒ�N`��i��L�ľa�x
�W��df#��'��$����F �����Ⱦ4���g���$Ӹ�~�(���̻�Gi<,K�<�	<��������>~��Y�3
���s⾪D�$�8�C�[��{�iމ�ݑ�$Ɣ�P��d���[}�5�]�#�:�p���徒����\��N��c��|���c)<ذ<��<��$��K��   �   ����\��Bq��D��ˁ��۠�~���xӾǒ���[��V(վ�����e��Ȧ����K�x/������*�p��3x<X�<���< Gc���!�s�ɽF�8�m"����־,��n�=��Wj�b�������w�����L��������U��a��������'l��,?�����׾LǓ��=9���ȽFG�@A�:8�<6�<Ț�< ��   �    ��;H�м���C�׽�@�>�E��}m�H������ ����(�����r��jL�F� �eN轵.��h@
� 9���<�T=�Z=���<ȢT�?���pB�OVq�����1��	�4�E;h�/r��æ���彿LqϿ&�ڿ��޿UIۿ�Hп7྿1���I(��e*i�H^5���΃���$p�NI	��v�h���d�<��=p�=`��<�   �   ο=8Ʉ<H���!�q����ν�y����Z�(��4.��[*��p�)��p`ܽaU��kD�ā��@m�;���<��#=�02=Ҧ=�]<xӼ������0�(����׈���U�c��%~��NCÿ��ܿ�������G�IN����tݿ��ÿe⦿G���`�U�p%���߾c����6-�7��t㩼h��<D�.=�/S=$�G=�   �   � s=��@=d�<��<�6U����~�\�>�ZҢ��*���^������q�x )����� A��Td�<
�=oH=^�_= �S=�=��<����۽(AR�R�������L6���r�6��T���/�ۿ�����<�����6�2���x�R��n�ۿk�����*r��M5��� ��O���UM���н:}��փ<�M;=֨y=��=�   �   �ڙ=�w�=z�f=��*= ��<��%<�\��8({��a���PռP�ɼ�K��h����P;X#�<(�=n;=��h=��=v�=Гh=�A=�{�;.�C�S�����l� ��U�{=H�&ل�V,��S%̿���ڸ���D(�D��;�(�h���l�ݪ˿w������2�F��������f��p�:&� ZP<`yA=�f�=��=�   �   V��=J��=�M�=�x=�E=��=0%�<h1~<(t<�J�;e�;��C<�(�<���<Ĭ!=�O=��x=�_�=��=B��=�t=V3=�ں:��^�f�
�$~�Ky̾���c�S�P$��j����ֿ������h��6^#��b&��_#�Һ�R���U����տ���Q����Q�:����Ⱦw��?�*~>���(<�D=u�="w�=�   �   \��=J��=��=b�[=N�%=<#�<��{<@i�; o��@�:� r���};`IK<t��<��=�SF=(�t=e��=��=慊=j�[=@`�<���춽�C�Yϩ�4D��B�_@��������ܿHe�2����0��?B���M�f R���M��B�V�0��s�����Lۿa~��?ᄿua@�jL�����^=�|��H]o�� =2Gr=�Z�=�   �   �t�=~��=ks=��==<�=T[�<���;�jȻ�-T�h:���de�H���.�:Xa[<���<|;(=�U\=���=�v�=�ׅ=��V=��<d��T`���Q>�t0��ԣ��?��݃�v����!ٿ .��S�h�-���>�J��,N��!J�b�>���-��������׿��������3�<�z� �Y��L�8��G��غ]����<�m=�=�   �   �v�=r�`=�(=��<@��;\�d�����0� VT�Xb�N�X�*�9�J��d��� l�9X�<�N=vnI=j�k=>�n=`�G=���<؎v�����8�0��������4���y��>��Iqοy���\����$���4��5?�B�B�`T?���4� �$���������Ϳ�;���w���2���������+�v`���t,���<��\=8��=�   �   �6=���<�y<8�z���)��s��~����޽Ƒ������?��1�⽋����'����=��è��u;�i�<!=��<=��,=���<'�3���V���u���V޾�*$��1d�� ������
�Pf��%��.�zE2��/�@�%����B7����&c�����c�b���"�y	ܾ�]�����;�� ͻ���<��?=^Q=�   �   T�<@.ٻ:3�������Y�.�8���S��pe��l�|�f���V���<�5�����lB���0��hC��4L<���<�4=�/�<�ǥ�T�X�����n�Vi���Y�ǜH����ui���V̿U����X�r�L�Bp�z���E����!�̿���� �� "H�	��S���Dk�������L��e��w�<P.=�=�   �   le���Cg��нл�H�S��鄾~$��T|������������G��Δ��D�K�Y�п"���۽j@|�\'Ƽ U*;�ډ<,�< �M������ʽ
�@�EꞾ���Om)�rb�� ������ծͿ�F迤b��0��d����������οƓ��O����c��)�<���\���,?���ƽ6�����:���<��<p��;�   �   >���tP��A(>���nԪ���оy��5�����	��c������V,Ծ�P���V���D��B�C+��,�����i�0��;@:�:ȗü�B���U���x�$���y	���8��2m��a�����������pӿ�߿pB㿯�߿�Կ�ÿ<g��8�����n��:�+�	�$���Qy�p �9���XŸ�@QU;�j"<�l)���ܼ�   �   ����7O�t
��#�Ǿ\������/�JoA�}WM���Q��!N���B�q1�'��P �HG˾���k&T�B�������V��`=�� L1:��D��7��A̽<�6�Ԑ��!ӾAU���:�og�ª���a��z&��&���;:��lS��?<��c������ni��<����]վ��.R8�S�ͽ�8��y<� ��:����\��'����   �   {�L������־=���T/��	Q���n�=[��;���ލ�����D��~Oq�-zS���1�nr��پA曾��O��=����������l� �Y��n���dy�@���J�L������־��Q/��Q�V�n��X���	��܍������A��hKq��vS���1�p�پx㛾��O�W8�����h���@�l��Z���Zqy�M����   �   �א�2&Ӿ5X�| ;��g�����d��0)��꺳��<��V���>�������	���qi���<����fվF��U8���ͽ8��x<�@�:����(�⼈x��x��&1O���ͥǾ���S��/�kA�SM�F�Q��N���B��1��#�bN �C˾d���!T�ۗ�����L��@2����0:x�D���7��H̽p�6��   �   	���	���8��6m�d��O��[����sӿ�߿LE�j�߿t�Կ�ÿ/i��ۏ��4�n��:���	�>&��gTy�-������Ÿ��yU;(�"< B'���ܼ�x��pE��E!>����TϪ���о�����<��h�]`�������A'ԾyL��*S���D��>��%��ؖ��@�i�p��;��:��üH���Y�My��   �   ����o)�Xub��"��3���S�Ϳ�I�}e�������:��[���>����οP��������c�u�)�@��4^���.?�@�ƽ������:X�<���<@�;�J���2g�-�н.��k�S�儾x���v��t�����H��B��@���P�����Y�p�"�'�۽�3|��Ƽ��*;�߉<$�<��N����E�ʽH�@�Eힾ�   �   �[�Z�H�v��Qk���X̿���^���������q�����F�!��s�̿#������.#H�۵�d���Ek�����4�L��2纬~�<�3=��=��<��ػ�"������⽰���8���S�Nhe���k���f���V���<�_��'��o:����0�`CC� NL<0��<6=X-�<�祻��X�����n�Ul���   �   z,$��3d�Z���ɼ������tg�:�%�F�.��F2�!/�4�%�L���7�����c��m��.�b�B�"�!
ܾ�]������@ͻP��<"�?=�cQ=v7=t��<`�<`�z�f�)��j��Ow����ݽ����n���S����Oy������=������>v;\v�<L!=֫<=�,=��<�'�ч�����w���Y޾�   �   �4�|�y��?���rο���4��l�$���4�z6?�*�B�.U?���4���$�H��~�����Ϳ�;��X�w���2�������t�+��_��Pm,���<�\=H��=!y�=��`=�"(=��<�Ԥ;��[����� �0�HT�Xb���X���9������� ��9���<�S=.rI=��k=*�n=��G=D��<X�v�?�����0�Y���f���   �   �?��ރ�M����"ٿ�.��T���-�8�>��J�j-N�Z"J���>�܉-��������׿����������<�5� ������8��F��(�]����<Bm=x��=.v�=M��=Hos=p�==��=lg�<ཋ; 5ȻhT�-��0Ke�H��@Ҥ:�r[<(�<F>(=�W\=���=�v�=�ׅ=��V=�<�
��c���S>��1��¤��   �   ۾B��@������(�ܿ�e�n��,�0��?B��M�f R���M��B� �0��s�P��4Lۿ�}�������`@��K������\=�z��xQo� =�Hr=�[�=���=̦�=b�=D�[= �%=�$�<��{< l�; [�� �:��|����};�FK<���<Ʈ=�RF=�t=ϐ�=V��=*��=��[=�[�<���`
C�GЩ��D��   �   �?�ރ������!ٿ�-��S�8�-�T�>��J�l,N�f!J�̧>��-�@��f����׿՝������<��� ����B�8��D��`�]����<:m=̀�=hv�=u��=|os=��==��=�g�<о�;p4Ȼ�T��,���Je�h���ڤ:�s[<��<�>(=�W\=���=2w�=2؅=��V=8�<��^a��hR>��0�����   �   ��4�1�y�z>���pο��������$�R�4��4?�X�B�lS?��4��$���r���C�Ϳ�:�� �w�>�2�7�����+��\��H\,����< �\=陂=�y�=`�`=#(=���<@פ;��[�4�����0��GT�
b���X�8�9�x������ ߳9��<�T=sI=��k=��n=��G=P��<h�v�򄡽9�0���������   �   *$��0d�Y���U�����,
��e��%���.�JD2��/��%�d��:6�є必a��x���b���"��ܾ�[�����������̻��<��?=xeQ=�7=��<��<Лz� �)�rj��$w����ݽW���<��������y��{��J�=����� Ov;�x�<�!=��<=أ,=���<`w'�;������(u��'V޾�   �   �X���H���^h��UU̿�����4�,����n� ���D�)���̿>���B���qH���J ��@k�������L��L�D��<�6=İ=T�<`�ػL"�������⽜���8���S�6he���k�l�f�j�V���<�,������9��v�0��=C��UL<8��<�9=�7�< �����X����n�'h���   �   ����k)�pb�]��g�����Ϳ�D�-`��ؒ���n�����a�鿆�ο����]����
c�b�)����Y��Z(?���ƽ��@��:��<��<�.�;�G���1g�ҁн��N�S�儾o���v��h�� ���6��jB��(���2���h�Y�(�"�}�۽j2|��Ƽ`�*;��<d�< �L������ʽ�@��螾�   �   ����	���8�0m�*`������i���0nӿ�߿�?�˲߿�Կ�ÿ�d��������n�]:���	� ��yKy����,���4��� �U;��"<�c&�4�ܼx���D��!>����FϪ���о����6��`�T`�������"'ԾXL��S��<D�@>��$��8����Oi�P�; �:@�üD?��vS�M�x��   �   �ѐ�cӾ-S�@�:�/�f�ר���_��
$������}7���P���9��Ͷ�����hji�b�<�����վl���L8���ͽN8��J<����:Pb��p��{w��$���0O�����Ǿ����N��/�kA�SM�@�Q��N���B��1��#�RN ��B˾<��8!T�^������xE��P�� �2:ȪD���7��<̽��6��   �   �L������־�~�N/��Q�C�n��V��G���ٍ�����>?���Fq�IrS��1��l��پ8ߛ�%�O�..�����\����l�`SY�Le���ay�P����L�o����־
��Q/��Q�V�n��X���	��܍������A��_Kq��vS���1��o��پN㛾N�O�(7��.��X���`Wl��`Y�(`��j[y������   �   ���,O������Ǿю��8�//�gA��NM�ޮQ�N�m�B���0�H � K ��=˾���^T�2��1����0��@ѵ���3:��D��7�L@̽��6��Ӑ�s!Ӿ<U���:�mg�ª���a��{&��$���;:��kS��=<��`���	���ni���<����9վ����Q8�ۢͽ�8�`<�@��:�T�� ���r���   �   kr���<���>�R��	˪���о��x��������\�:����6!Ծ.G���N��2 D��8�9���x��@�h��+�; 6�:8�üA��HU�F�x����s	���8��2m��a�����������pӿ�߿pB㿰�߿�Կ�ÿ8g��4�����n��:��	��#��Qy����d������� �U;P�"< j%��sܼ�   �   (6���$g�lyн�����S�ᄾ����q�� ��g�������<���������t�Y�t�"���۽!|�T�ż�s+;��<�$�< hL�D��9�ʽ��@�*Ꞿ���Km)�rb�� ������׮Ϳ�F迥b��2��f��������� �οÓ��L����c���)�!�ﾸ\���,?�=�ƽܸ��U�:T�<�
�<0[�;�   �   ��<0sػ����������8�.�S�D`e�L�k�-�f�o�V�<�<�p�����/�� �0�(	C�H~L<p��<�>=4>�< ���"�X�D��hn�Fi���Y�ŜH����ti���V̿W����Z�t�N�Dp�z�� F�����̿���� ���!H����6��<Dk�x�����L� ��,��<H8=��=�   �   7=���<��<�nz�V�)�Zb���m��M�ݽd{�����������⽳n������=������
w;��<\$!=��<= �,= ��<q'���� ���u���V޾�*$��1d����� ��� ���
�Pf��%��.�~E2��/�B�%����B7����&c�����^�b���"�f	ܾ�]��4��
����ͻ���<B�?=�gQ=�   �   �z�=<�`=`((=x��<��;��[�4s���0�.:T���a�L�X�T�9�j������ ,�9t�<f\=�yI=�k=��n=,�G=d��<��v�<����0���������4���y��>��Iqο{���\����$� �4��5?�D�B�bT?���4� �$���������Ϳ�;���w���2�������r�+��_���k,����<��\=i��=�   �   �v�=$��=�qs=��==��=�p�< �;�Ȼ��S����.e���� ��:��[<��<�C(=>\\=� �=�x�=�م=J�V=��< ���_���Q>�o0��ԣ��?��݃�x����!ٿ.��S�h�-���>�J��,N��!J�d�>���-��������׿��������2�<�v� �R��.�8��G��X�]�,��<"m=���=�   �   �c�= \�=�w^=�J'=��<��/<`C3�Pd\�����8���;��� r� f����<�^�<$S=�2S=Ԁ{=b�=�*y=N?6=H�H<�(�^]��p�x��Ҿ�4"�tuj��<����п�|������9�=T�nk���z��8����z���j� �S��8�����h�ο�����g�� �@�ξ]�s�k�������+u<��@=:�=�   �   �(�= �p=� B=�=0\�<�^��Q����༸���������7켤�����N��[V<H��<p�6=+e=�P{=�$n=�0=�G<�V#�����s�P�;U��6f��v��A3Ϳ@R �'��E6��5P��jf���u��{�ȫu�$[f�Z�O�R�5�pf�b���ԇ˿#���?�c�� �o�ʾRvn���P���r<T;=~�x=�   �   *�S=$�,=��<���;��z�ܮ���c��ސ�w�������ݦ��(����l��_ �`����PZ;XH�<n� =��H=$FL=X�=x�?<������C#c�7Z��F!���Y�%f���	ÿ����t���,���D�L*Y�Ng��l��>g�_Y���D���,�\	�(��W����;����W��x�J����_�Kݽ���h<Ұ(=x�V=�   �   ��<�[<��-�4 ��O���X˽x�$���%��X*��(&�?������ѽ1<��d�-��c���)<p��<.+=4"�<�'<X}���ǽ��J�-(��>$���F��Ĉ�3#�����N�������3��E�.�Q�lV���Q��F�tG4����n��/࿧~��Z���:E�v���(��QG��'½H'�0M<��=̖=�   �    �t�$P�>g��f�ڽ:c�ֆF�q'n��↾�3��S���8?����q��J�Į�n�⽨���:�@mz�X�d<̏�<0��;�ʼ�ϥ��,���A��$.��Uq�*؞�N�ǿΑ�����X��b.��v8�^-<�6�8��/�� ���cH�ȿ3Ğ���p��o-�X��"���B�)�Ж��������<|��<���<�   �   �3��:��"���_M�F0��[��n�þp[ھ%7�:�7�D4ܾ� ƾp���쉾�uR�b�.����@��&�� ^: k�9y���;��[�
�h�v��Zžҍ��L�޽��֧��P'п��'	�в����X!��v�P���
�3���][ѿcg����ZM�
r�Y�ľR0u��	��~�T���  ;`P>;`�W��   �   D}̽��&�ùt�5��1�Ӿ�S ��]��N$��.�q2��^/���%������l`׾|,��r�y�+���ҽ�c_��Ͻ��(��쏼6�A�eҽi�?�­�� ��&� �^�{�����ʿC忏���·�:;��)��a��E��Ά̿����m��	L`��w'�K��Tݜ�A�?��н�>�ஆ�0��\q��~aU��   �   �D.�lS��d������)7�B�8�#�S���h��v�|�{���w�>�j�J�U���:��_�0�����薆�g�1�P	Խ�^�T�Ӽ@ژ���	�VΓ�����Kk�Cٴ����b/��qa��h������������ɿX�Կ[ٿ\�տ('˿BT��4����ԋ���c���0�q�����l�������xN��9����ʼ0zW��KϽ�   �   ,����[���n�2�*���S�9{� ��|՜��å�r��:^���띿(k���	~��aV��-�d
�/����/���&�Mi����>�,|üD���`<��ߺ�ѕ$������V���k�v�*�I�S�4{�K���Ҝ������	��i[��N靿�h���~�^V��-�,�ߤ���-���&��e���>�T~üL����<�$纽 �$��   �   vݴ�H���e/�va�/k�����������ɿ��Կ�ٿl�տ*˿�V��p����֋���c���0�=���!��y�l������@N�,2���qʼ�mW�CϽ�>.�fO��A��A���o3��8�v�S��h���v�^�{���w���j��U���:�x\�9���)��
���`�1�
Խ�^��Ӽ�ޘ�֘	��ӓ�����Qk��   �   ���&���^���������ʿf	�����t���<��+��d������̿s����	��uN`��y'�޴�ߜ�V�?��нr>�D���`��t]�� SU�ts̽b�&���t�#
��(�Ӿ<P ��Y��J$�ʪ.�4{2�lZ/�ƌ%�m����][׾h(���y�j+��ҽD[_��ƽ���(��򏼌�A��
ҽ"�?�$����   �   7��.�L�ƿ������)п��)	����V��!�Px�ʁ��
�\���']ѿ�h��>��	M�:s���ľ>2u��	�ȅ~�$����N;��>;�jW���3��0��Ý��WM��+������þUھ�0龝��31�I.ܾ��ž����(艾DoR�q�ֹ��L�?�,�� �^: -�98����?����
�d�v�~^ž�   �   y&.��Xq�ڞ�w�ǿJ��\��<Z�vd.�tx8�/<���8��/�� ����I��ȿ!Ş�%�p��p-����⽔���)� ���D���0�<���<`�< �q��1�]��ҕڽf\� F��n��݆��.��w���둾�:����q�$�J������M��0���y�(�d<���<��;H�ʼ�ӥ��,��������   �   �F�Gƈ��$�����l�� ��V�3�~�E�ʩQ��V�(�Q�F�nH4������ 0�P�����;E����)��NQG�I'½�#�H#M<��=T�=4��<�\<�V-�����E���M˽|����%��Q*�~"&�:�����U�ѽ/4��d�-��b��*<d��<�-=#�<�'<���6�ǽ�J��*���%��   �   ��Y�Ig��Wÿ���u���,���D��+Y��g��l��?g��_Y�h�D�4�,��	��������;����W��x�B����_�| ݽ����h<~�(=$�V=��S=l�,=̪�< �;dz�����c��֐�7�������զ�/!��\�l�.T �������Z;�T�<�� =��H=@GL=Ƅ=��?<������!&c�F\���"��   �   8f��w��<4Ϳ�R ��'��F6��6P�Vkf�r�u�8{�P�u��[f���O�n�5�vf�V�����˿�����c�A ��ʾiun�i���M�0�r<;=��x=�*�=B�p=�%B=f�=�h�<�\\��B�������������*켄폼 zN��lV<���<ʦ6=�,e=pQ{=v$n=��0=��G<[#�C����s��;l��   �   Svj�g=��"�п(}���Е9�X=T��k��z��8����z�`�j���S���8����ԇ���ο�����g� �*�ξ��s������h6u<��@=�=8d�=�\�=�x^=�K'=���<��/< :3��b\������8���<�� r��k���<�\�<R=�1S=�{=��=�(y=>=6=��H<��(��_���x��Ҿh5"��   �   7f��v��\3ͿDR �'��E6��5P�&jf�&�u��{��u�ZZf���O���5��e�L�����˿Q����c�}�ϭʾ�sn�z��2K��r<,	;=J�x=�*�=��p=�%B=��=i�< U\��B����༨�����`���)�폼 vN��mV<���<*�6=-e=R{=B%n=Ƃ0=��G<fX#�B���Xs�ּ;���   �   ��Y��e���	ÿ	��Bt��,���D�h)Y�<g��l��=g��]Y���D���,�z��������:����W�Dw�6����_���ܽ
��X�h<��(=��V=� T=�,=���<��;�bz���^�c��֐���f���wզ�!����l��S �������Z;�U�<�� =��H=�HL=�=H�?<������F#c�)Z��1!��   �   7�F�lĈ��"��̗࿲�������3���E�¦Q��V�&�Q�TF�
F4�~��V��:-�
}�����8E����5&��rMG� "½<�5M<��=J�=ħ�<�\<pT-�����E���M˽i����%��Q*�b"&�������ѽ�3����-�`�b��*<���<0=t)�<��'<y���ǽ�J��'���#��   �   #.�3Tq�3מ��ǿ9�����|W�`a.�u8��+<�x�8��/�> �����E�qȿb���p�fm-��|뾂���`�)�ؐ���x���<�Ʃ<��< Qq��/�g]����ڽO\��~F��n��݆��.��j���둾�:����q���J�����������.���y���d<���<`��;��ʼ�ͥ�3
,�,������   �   ���[�L�����]����%п��&	�X������!��t��~�
�J����Xѿ"e��8��CM��o���ľ�*u��	�Tx~�L��� �; ?;aW��3�!0������WM��+������s�þUھ}0龎��"1�5.ܾv�ž����艾oR�$����@�?�h����_: D�9�n���8����
���v�2Yž�   �   K��5�&���^�����)����ʿ�忟���(���9�8(��^�����̿����-��FH`��t'�����ٜ���?���н�>�����`���U���PU��r̽$�&�X�t�
���Ӿ8P ��Y��J$�Ū.�.{2�eZ/���%�b����>[׾G(����y�+��ҽ`X_�d�����(�`�����A�f ҽ��?�ث���   �   �ִ�����_/��na��f������,�����ɿM�Կ,ٿ#�տ�#˿CQ��o���zҋ�c�c�
�0��������l��� ���(A�� ���eʼ4jW��AϽ&>.�IO��/��4���j3���8�r�S���h���v�X�{���w���j��U���:�j\������ܓ���1��Խ�^��vӼ�̘���	�'ʓ�����Gk��   �    ���kS���i���*���S��/{��	��М�н�����tX��j板f��� ~��YV�&-������)���&��\��$�>�dü$���0�;� ޺�P�$�^����V���k�r�*�F�S�4{�K���Ҝ������	��e[��K靿�h���~�	^V��-������R-��h�&��c��p�>��mü ���"�;�qں�-�$��   �   :.�jL��W��B���]0�]�8�K�S�f�h��v�;�{�r�w���j�W�U���:��X��������Ώ��Ɗ1���ӽ�^�lgӼŘ���	�̓����iKk�'ٴ�~��b/��qa��h������������ɿW�ԿZٿZ�տ%'˿@T��/����ԋ���c���0�a�������l���q ��PG��$��bʼ6dW��<Ͻ�   �   l̽q�&�
�t����Ӿ:M �8V�G$���.��v2�"V/���%����n�$U׾$#��|�y�~�*�-�ҽ�I_�������(��ڏ�F�A��ҽ��?��������&��^�{�����ʿD忐���·�:;��)��a��B��ʆ̿����h���K`��w'�(��!ݜ���?��н�	>�����@���L��HU��   �   ƀ3��(�����~QM��'��O����þOھ*���*��'ܾx�ž=���X㉾gR���䮹���?� �� �a: ��9�j��49����
���v��Zž̍��L�޽��֧��P'п��'	�в����Z!��v�P���
�0���Z[ѿ`g����QM��q�2�ľ�/u��	�N�~�����@�;`<?; GW��   �   �go��V��/�ڽ�V�
xF��n��ن�1*������,摾6���q��J�С�������@�@y��e<�< ��;��ʼ�ͥ��
,����0��$.��Uq�+؞�O�ǿϑ�����X��b.��v8�`-<�4�8��/�� ���cH�ȿ/Ğ���p��o-�=��������)���������(<ʩ<�<�   �   ��<'\<p+-�����=��D˽�� �����%� K*��&����z���ѽ+*���-���b��D*<���<�6=3�<��'<xu����ǽD�J�(��9$���F��Ĉ�5#�����N�������3��E�.�Q�nV���Q��F�tG4����n��/࿧~��X���:E�l���(���PG�2&½��p-M<4�=�=�   �   �T=~�,=���<�F�;�;z�@����c�!ϐ� �����#ͦ������l��E ������[;h�<� =��H=�ML=ʊ=��?<n�����#c�(Z��E!���Y�&f���	ÿ����t���,���D�L*Y�Pg��l��>g�
_Y���D���,�\	�(��U����;����W��x�7����_�z ݽ���X�h<(�(=��V=�   �   V+�=0�p=H(B= �=�q�<�[� 6����"�����>�����ݏ� N�h�V<ܛ�<�6=N1e=�U{=b(n=��0=ГG<�U#�����js�J�;T��6f��v��C3ͿAR �'��E6��5P��jf���u��{�ʫu�$[f�\�O�P�5�pf�c���Ӈ˿#���<�c�� �e�ʾ6vn����<O���r<�;=
�x=�   �   �t=V�b=J�5=�w�<(�L<�Ӊ�t7������l��z�*�\!�L:������ܸ�(Z4<�m�<&0=�]=r�o=�[=��=�����}�w��@H���E���<�)e���巿���(*�`S5�&4W��x��
��9 ���������z���Ix��eV��O4� �:��X0�������:��<���&�����Z�t� *W9ƍ=�z_=�   �   �7b= �I=�=(Z�<�y�:\~���r
�5@�c���o�pe��rD����?�� z��q�<^=�tD=\e]=ȖN=Z=	=����0�v�j�$���c�sY9�s���hƴ�K�꿎���2�S���s�6��`̑��M���ё�����Ts�&vR�C1�6��B�迠2��淃�_b7�́�$���?�V�n� ��8�=T.S=�   �   ��)=�q�<�R<(��jF
�:l�B֡�]�ĽRP۽����ܽ0Wǽ)[���t��m�(�:�Ƚ5<��<�$=�i(=��< ���|#e�
������A侁#/�G|������!߿�s���(��}G�*Be���zp��g�����RU�"Xe�IG�t�(���
���ݿ4y��y�y�I�-�����>�����]��;�ԕ�<<Y-=�   �   ���<�Tʺ8[���x��½H��|�"��;��K��Q�B�L�p=�"U%����DȽ����lX���g_��<,|�<�M�<�6m�2�K��� �!v�Yξ)8�hAf��y���3ͿP ��|36��P��>f��~u�8{���u���f��P��6�\ �0 �̅̿0�����d�.
��|̾;s�m���E��Z�`Z�<<k�<�   �   7���J�T�B���#@�/dr�k������z���ű��/��a���s���#v��C�3G��Ӿ�L�S�x����X:`�;�U���1��6۽,9S�!ղ�����J�QQ��o[��Ћ�r 
�Rd!��&7�&dI���U��kZ�JYV��@J��8��"��j
����K������I�e
�0���nEQ��ؽ��+� uϻP��;`.	;�   �   N6�������3�bz��P��ޤƾ�;�
� ��	��"��	����"��GAɾ�ܤ���~�-�7�?��ً����@j��s���Ჽ`-�P=��w���'+��Ym��X����Ŀ4��x�
�r��|�+�8�5��.9�6�Ĕ,����0��uU�1�ſ����+�m�+��辮���9�+��°����H�a�rT�$����   �   h��NJN�0�����žO�����V-�Kq?�b2K��~O���K�T�@�-�.�AQ�m��r�Ⱦ����Q��M�����)�d�ܼ��n�����%j�L���3�
��(B�^���Wm��srƿ��翠��־�f���~�d����|�����vȿ؉������W�B�^�
�*ź��j�F���؋�8���Լ<c$�<ߙ��   �   Z�V������vܾ(t��4��V�au�����v���S��􎿓���DSw���X��=6�*N�$^߾���(�Y�����+��26�Bm��Z�YEǽ(�.�����H־����L�{f��/e�����{�ӿ����]�y���6���J��JտCټ�
꠿o���`�M�Z
�9�׾򩎾k�/�,�ǽF!Z��t�h 3�G�������   �   �朾wf⾁�nG��ku�y���C���G��L'������6о�fK��U���t���x�+7I�'�����Di���+M�Lb������ �-�>:-�l��!��BK��✾�`�
�1G��fu�����6������#������
;�nH�����xr���x��3I����ڪ侗f��^(M�,^��S���@�-��?-�mq��w)�� HK��   �   �L־����L��h���g����ԃӿ;��ta���]:���M��Mտ�ۼ�*젿,����M�i�$�׾⫎���/�N�ǽ(!Z��p��3�Z|�����j�V���pܾ�p��	4�4{V�u�����,s��Q��8������Nw�h�X�e:6�TK��Y߾�����Y����~(�� }6��o��Z��Kǽ��.�*����   �   Ң
�R,B�z����o��Yuƿ��h�����`�����@�p�������鿚ȿ����Z���i�B�� �$Ǻ�.
j�p���؋�(���ԼX$�י�֐��BN�{���ʛži�����zR-��l?��-K��yO���K���@�=�.��M�Ig��ƕȾ����Q�/J�������)���ܼ|�������$+j�&����   �   �*+�l]m��Z��=�Ŀ#��"�
�L����+�R�5��09�6���,�~��n��}W�ѢſCÜ��m�s+����Ǫ��R�+�Wð�p����a��NT������-��X�뽂�3�"Yz�^K��ƾ�4�g� �	��?�	�v������;ɾvؤ�d�~���7�ڶ��Ӌ�t���j��s�����岽,-�)@�����   �   :�J�S��]��?���
��e!��(7�8fI��U��mZ�D[V��BJ�88��"�fk
�4��'L��Q��+�I��e
����CFQ�ؽ��+��Rϻ���; �	;�����I��踽���#@�:[r�r���6���Cu��o����*��Y��ro��v�l�C��A�F˾�ڝS�D�����:�)�;�a���1��;۽
=S��ײ����   �   �Cf�({���5Ϳ,Q �V �56�nP��@f���u�8{���u�V�f��P���6�!�� ���̿������d��
�l}̾z;s��l���E� "��d�<�y�<�ΐ< �Ⱥ�<꼎�x�T�½����"���;�l�K�h�Q��L�(i=��N%����z;Ƚ"|��PA����^����<@��<�N�<�Zm���K�&� ��
v��[ξ:��   �   [|�ʳ��^#߿rt���(�.G��Ce�D�Mq��/�������lV��Xe��IG�ք(��
���ݿhy����y�\�-���ᾩ>��B���]� s���<r^-=�*=��<�7R<a��8
���k��͡�=�Ľ�F۽����ܽ�Nǽ�S����s��b�P�:�p�5<��<"�$=&k(=ܿ�< I���(e�4��:��QD�%/��   �   ; ��\Ǵ�g��2��| 2��S���s�����̑�mN���ё�D���
Us�HvR�C1�0��!��u2������b7�.�ﾜ���>�F�n� ��8�=�1S=�;b=��I=~=�f�< [�:�n���j
�.,@�
c��o��ge�kD����3�� 	蹌y�<"=PvD="f]=��N=�;	=�����v�:�w ��re�Z9��   �   �e��4淿-��|*��S5��4W�\�x��
��M ���������W��@Ix�VeV�RO4�������/��+����:��;���%��d��x�t� Z9��=�|_=��t=��b=~�5=�y�<P�L<�̉�$6������0����*��!��:�8����主�U4<�k�<�$0=t�]=��o=� [=n�=�좺�}�ڶ�1I��G����<��   �   �����ƴ�h�꿒���2��S�\�s����	̑��M��ё������Ss�LuR�ZB1����,�迲1��!���'a7�������=�^�n� d�8�=|2S=H<b=��I=�=�f�<�`�:�n��xj
�,@��c���o�~ge��jD���x3�� ��$z�<j=�vD=�f]=X�N=6=	= ۰���v�����/d��Y9��   �   |�J���x!߿Bs�x�(�L}G�NAe����o������"����S��Ve��GG�f�(���
��ݿ�w��p�y��~-�-��=��,�B�]� �����<�_-=�*=X��<h9R<�_�l8
�p�k��͡�$�Ľ�F۽���˼ܽ�NǽYS��R�s�Hb��:� �5<X�<F�$=�l(=���<����"#e�������A�h#/��   �   �@f�y��3Ϳ�O �V��26�nP�`=f��|u�@{���u���f�,�P�~6�� ���̿����e�d�Q�.z̾7s�g��R�E����dk�<�}�<xѐ<��Ⱥ�;�"�x�%�½	����"���;�]�K�V�Q�ФL�i=��N%�d��(;Ƚ�{���?��@�^�� �<��<`U�<�m���K�,� �Tv��Xξ�7��   �   d�J��P��YZ��e�俊�	�,c!�D%7�nbI���U��iZ�"WV��>J��	8��"�i
�l��I���
��f�I�c
�1���
AQ�!ؽt�+��"ϻ �;��	;�����I�@踽���@�([r�j���,���;u��c����*��J��`o���v�;�C��A��ʾ�r�S�l����O:�J�;�0���1��4۽�7S�Բ���   �   &+��Wm�8W��
�Ŀ(��8�
������+�D�5��,9�6���,�$������R￩�ſڿ����m�Y+���辝�����+�Ļ��x��`�a� >T�L����,��ͤ�U�3��Xz�PK����ƾ�4�b� �		��7�	�l������;ɾZؤ�%�~�:�7����ҋ�r����i���s�|���ݲ�n-��;��{���   �   ��
��&B������k��Lpƿ6�� ��&������|�j�ԝ������鿉�ǿO���ܭ����B���
�&����j��}�Hы����uԼ�S$��ՙ�j���BN�f�����ž]������vR-��l?��-K��yO���K��@�0�.��M�,g����Ⱦ���H�Q��I�s���P�)�0�ܼ2��������"j�����   �   �D־����	L��d��c��m���}ӿ}��[Z�����<3��G迖Gտ&ּ�B砿	���`�M�&�G�׾6���ʗ/�n�ǽ�Z��f�d3�Qz��G��	�V���pܾ�p��	4�/{V�u�����*s��Q��5�񁇿|Nw�\�X�W:6�DK��Y߾z��
�Y����V&���v6��e�P�Z��@ǽ�.�}��   �   �ߜ�]�s��G��bu�X󐿍������ ��g����ɾ�-E������o���x��/I���,��5b���!M��S�������-�b1-�;i��S���AK�z✾�`��	�-G��fu�����5������#������;�kH�����sr���x��3I�������_f���'M�;\��[���J�-�h2-��g��$���=K��   �   fV��잾ylܾ�m�
4�wV�]u�!���cp��"N��M��#Iw�|�X�66��G��S߾����Y����g���m6��a�Z�Z��Bǽe�.�u����G־����L�zf��.e�����{�ӿ����]�y���6���J��Jտ?ټ�꠿i���R�M�J
��׾������/���ǽ~Z�2i�63��v��=���   �   ���N=N�ʝ���ž��������N-�Hh?��(K��tO��K�=�@���.��I�3`��ɏȾ,����Q�	D�B����)�X�ܼ�1�����(%j�"���)�
��(B�]���Wm��rrƿ��翠��ؾ�h���~�d����|�����qȿӉ������J�B�M�
��ĺ�j�4��ZՋ�\���sԼ�N$��Й��   �   �&��r�뽲�3��Qz��F��b�ƾ�.��� �d	�>�o�	��}��龡5ɾ�Ҥ��~��7����ʋ����x�i�`�s�$��n޲��-�=��\���'+��Ym��X����Ŀ5��x�
�r��|�+�8�5��.9�6�Ĕ,����0��sU�/�ſ����$�m�	+����j���c�+�O��������a�00T��x���   �   X��@�I��߸�6��r@�PSr�帏�)����o��Ժ���$�����Zj���v�T�C��:�տ�� �S��n�� �: ��;���� 1��4۽�8S��Բ�����J�RQ��q[��ы�t 
�Rd!��&7�&dI���U��kZ�JYV��@J��8��"��j
����K������I�e
� ����DQ��ؽx�+��-ϻ �;�D
;�   �   �ܐ<��Ǻ�$�`�x��½���h�"�̍;��K���Q�,�L��a=��G%���50Ƚqr��� ���^�T�<ĕ�<`�<��l���K�� ��v�Yξ$8�hAf��y���3ͿP ��~36��P��>f��~u�:{���u���f��P��6�Z �0 �˅̿.�����d�%
��|̾�:s��k����E�`���l�<,��<�   �   �*=x��<hUR<�;�T-
�4�k�ơ���Ľ�=۽$��U�ܽiEǽ�J��|�s�RT�m:��6<�#�<�$=r(=,��<@k��� e����v���A�#/�H|������!߿�s���(��}G�,Be���zp��g�����TU�"Xe�IG�r�(���
���ݿ3y��w�y�D�-�x�ᾬ>��E�X�]��0����<Na-=�   �   =b=��I=�=�n�<���:�b���c
�B$@�^c���o�R^e��aD�8��p#�� Q乸��<�=z{D=�j]=ؚN=R@	=�x����v�4����c�rY9�s���iƴ�L�꿎���2�S���s�6��_̑��M���ё�����Ts�&vR�C1�6��A�连2��巃�\b7�Á����?���n� آ8n=B2S=�   �   JY=�E=ʾ=ȣ<@��:,↼����:���\�Ii���^�\�=���	�ߎ��VC:���<4=yC=�W=��@=��<��N�B�����9������R�rY��=Z˿X��^%�VJ�;r��[��"���K����4��N����������nq��I��
$����&�ɿ�#��� Q�3�	��]����7��!��P7C���<�B=�   �   xE=x{*=�8�<��<��/�@*���G����o铽5����Д�����D�K�ؒ���@�8�< ��< (=�NC=$:3=<e�<��P�A5��v�5�񔦾�m�9O�ɻ����ǿā��<"��TF��Sm��E��ha�����0�����Z�����&�l��E��W!�ȫ �ʆƿ뚒��_M��9�6�����3��Û��AE����<Z�4=�   �   b�=d+�< �:�%��l�H��ř���ɽ����(�B�������i̽g̜���N���¼�Y:`��<�g=l�	=��<h�Z�팔�[Q*�͌��ԥ ���C�] ��F��hf���%���;�ԇ_������-��`��������R������W_�>R;�6���1��1���S8���vB�$B���'���(��U����O���<D�=�   �     �;(_b���1�O1��2��1�9?�AQZ���k��Kr��l��[�:;A�Zc����6���W8�Hv����;�<��%<8Ey����E������(�c2�6���������|����+��/K���i��6���f��Ď����������cj��~K��+����|(�r䭿/8��d1���羼���q��ׄ�Xun� X/<p�<�   �   �Q �bz������,'�P�_�"����r��EE��j&ž��ɾ��ž=i���쥾 .��@�b���)�_�u��~���3.��s��P|����o����K�s��ʾ�>��b�������ɿg{��ʙ��3��WL�p�a��p��!v�~3q�j�b�r=M��3�F�����n�ɿt���5za�����ɾ�gr�8����l�d���"����   �   �٬�T��LHR��������3�w������"��}������<��f��SN�����zU�
6��e��N�A�9ܼdi�H�W��=۽��I����~_���?��,���h����ٿ�{����T.���>��aJ��N���J�R�?��
/�����"��xڿWѭ�]Q����?��5�X���5I���ٽX-U�D�ۼH,ռ��<��   �   ��NLo�ݨ��#ྷ�j%)�=:B�iV�t�b�C�g��c��CW���C��*�ʆ�L�������ur�r! �Ľ�+h�X�&�V�K��������\�����Ӿ����Y�݃���4��M�ۿ�) �������|�&�f*��D'����B�����ݿ^A��/��E�Y��;�{�Ӿ@��� ��2�����I���#�&d�����   �   P?x�(L���S��iu"�D�I�F�o�񁈿C���%=���T������Y���������q��K�� $�����J2��k�z�^� �oýl�u��Q�\������L��K���G򾏢*���c�����ְ��Ͽ���]���n����V��; �i�뿹�п�@��>3��)�e��+��������L��k�q厽D]P�:is�iF��R+��   �   �����q�,�z�^�����6��m���2rǿ`ҿ1[ֿv�ҿH�ȿ�䷿Vr������4�`��{.��� �|K���Km�����5��*�l��=l��.�������k�k貾������,�у^����(������nǿw\ҿ�Wֿ��ҿ
�ȿ�᷿�o��]��`�y.��� ��H��Hm�=��4��X�l�Dl�n4��B��L�k��   �    M��*���c�M���ٰ�U Ͽ���E���p����B���< ����z�п6C��%5��)�e�D�+�˂�9�����L�6n�m厽�XP��_s��>���%��7x�G��MM��sq"���I��}o�	��-����9��wQ��y���~��������q�4�K��$������.��J�z�	� ��ký�u�\�Q�2��i��P%L��O���   �   ���UY�-����7��y�ۿ�+ ��������&��
*�G'������>�3ݿEC���0����Y�W=���Ӿ����N��������I�`�#��d��������,Do��ר�h����!)�o5B�JV�)�b���g�Бc�?W�e�C�N�*����#���󪾝or�H ��Ľ<&h�z�&�*�K����v��S����Ӿ�   �   ��?��.��%k��h�ٿh}�t��r.���>� dJ�b�N��J�X�?�t/����#��zڿ�ҭ�iR���?��6�����tI�K�ٽ�*U���ۼռ��<�QЬ���L@R�������,Ᾰ�����Z��y�����ԟ�v|�WI��
���xtU�f1�_��<�A��1ܼTj�$�W�C۽$�I�����a��   �   �b�[�����ɿ~��b���3�ZL���a���p�Z$v��5q�t�b�?M�\�3�D�t�����ɿP���m{a�°���ɾ|hr�b����l���獻���VC � q����㽈%'���_�.���~m��^?��H ž��ɾ��ž�c��y祾�)����b���)��U轔����.�@c�����z�o������s�1�ʾ�@��   �   h7��������⿶��*�+��1K���i��7��h��7Ŏ��������ej��K���+�*��M)�孿�8�e1�"������q��ք��en�(o/<��<ps�;�)b��1�7'��Kv�F*��1?�+IZ�0�k�/Cr��l�w�[�[4A�`]����
���K8���u�@,�;���<�%<�Ny����������+�&e2��   �   �!�����h���&��;�X�_������.��^���������R������W_��R;����2��l���r8��wB�B���'����(�YT���O���<�=p�==�<�g�:���d�H�����I�ɽ��ｴ#�����0��`̽Ŝ�d�N�ؕ¼�[:X��<hk=�	=��<��Z�я���S*������ ���C��   �   ������ǿb��|="��UF� Um�kF��b��g���0��c��fZ�����P�l�"�E��W!��� ���ƿ����z_M�y9�������3�F��4E� �<�4=�E=z�*=�D�<�<�t/�����G�� ��w䓽U����˔�>�����K�b����@��< ��<�!(=�OC=�93=b�<(�P��7��u�5�e����n��O��   �   �Y���Z˿����%��J�x;r�0\��M���b����4��6������s���nq�I�P
$������ɿ=#���Q���	��\��4�7�����*C����<�B=�Y=\�E=�=�ʣ<��:0������:�t�\�Ii���^���=�\�	�$Ꮌ�C:T��<�=�wC=H~W=��@=8��<�N�y����9�������R��   �   ������ǿց��<"��TF��Sm��E��a��j���/��h���Y����� �l�<E�<W!�0� �ƅƿ����^M��8�������3������,E���<�4=XE=ڀ*=<E�<p<t/������G�� ��h䓽D����˔�,���~�K�0����@��<���<r"(=BPC=�:3=�d�<��P�76��9�5�v���n��O��   �   = ��	��f���%�N�;��_�:���*-�����'���� ��Q�������U_�Q;�:��
0����67��3uB��?��&��=�(�YQ��X�O���<��=��=|>�< w�: ���H�弙�2�ɽg�ｨ#�������`̽�Ĝ���N�̔¼ 1[:��<�l=��	=
�<�Z���bQ*�Ҍ��ͥ ���C��   �   �5��c����������+��.K�$�i��5���e����Ĝ�������aj�}K���+�h��~&��⭿�5��b1���羆��[n��҄�HPn� }/<X��<`�;�%b�b�1��&��v�2*�~1?�IZ� �k�Cr�۽l�b�[�@4A�?]�G�����4J8�@�u�p9�;���<��%<�8y�ɾ�����$���'龏b2��   �   ^
b�����S�ɿ�y��Ș��3�@VL�f�a���p�<v��0q���b�D;M�2�3���G���4�ɿ����Jwa������ɾ�br������l����ō�����A �up��Q��h%'���_�$���rm��T?��? ž��ɾ��ž�c��i祾�)����b���)�LU�� ����.��@��Pr��\�o������s���ʾ�=��   �   -�?��+��dg��Ԩٿ�z�.���.���>�b_J���N�D�J���?��/�Ą�6!�vڿ ϭ�sO����?��3�����:I��ٽ U�`�ۼ�ռ�<�fϬ�Ľ�@R��������,ᾳ�����V��y������ɟ�_|�=I������-tU�
1�	^���A�,(ܼ�[�0�W��:۽��I�P��g^��   �   ���GY�W���	3���ۿl( ������b�&�0*��B'����B�����ܿ�>���,���Y��8��Ӿ������8󰽖�I�6�#�`d�>���{���Co��ר�W����	!)�i5B�DV�$�b��g�ȑc�?W�[�C�B�*�����⾮�<or�� �&Ľ~!h�"�&��K�����%������\Ӿ�   �   uD�@�*�z�c����c԰�:Ͽ�������l����P��9 ����Q�п�=���0���{e�|�+�z�������L�Qb�uݎ�$NP��Xs��<��%�?7x��F��:M��jq"���I��}o���-����9��tQ��u���y���򅉿�q�'�K��$�~���|.����z�J� �~iý�u�ĪQ�,��x��L�zI���   �   F岾������,�@�^�ױ�����.���skǿYҿ�SֿZ�ҿ|�ȿ�޷��l���뉿�|`�0u.��� ��C���@m����%+����l�T4l��+������k�A貾������,�̓^����'������nǿw\ҿ�Wֿ��ҿ�ȿ�᷿�o��W��`�y.��� �MH��lGm�8���0����l�r5l��)��h���k��   �   "2x�TC��^H��On"�¤I�syo�u|��U����6��LN��I���`��������q�o�K��$�����])���z��� ��aý��u�(�Q�1�����*L��K���G򾆢*��c�����ְ��Ͽ���\���n����T��; �e�뿵�п�@��83���e��+�b������L� i�EᎽ�PP��Vs��8���!��   �   P���=o��Ө�7ྸ��G)�1B��V��b���g�z�c��9W���C�ܷ*������ngr�� �.ĽBh���&���K����{��	�����Ӿ����Y�܃���4��L�ۿ�) �������|�&�f*��D'����@�����ݿYA��/��9�Y��;�F�Ӿ淆�ߕ�����L�I�F�#��d������   �   �Ȭ�(���9R����
���&�O����P�hu�ю������u�NC������lU��*�mT����A��ܼPἺ�W�1;۽�I����o_���?��,���h����ٿ�{����V.���>��aJ��N���J�P�?��
/�����"��xڿSѭ�YQ����?��5����VI��ٽ�$U�4�ۼ�ռ�<��   �   88 ��i���㽀'�U�_�Έ��vh���9��Nž��ɾƺž�]���᥾�$���b�A�)�LI�o����p���-�P���h��J�o������s���ʾ}>��b�������ɿj{��̙��3��WL�r�a��p��!v�~3q�j�b�r=M��3�D�����k�ɿr���-za�����ɾ�fr�0���l� �����0���   �   ���;� b���1����l�@$��*?��AZ���k��:r�l�l�7�[��,A�\V�5��t���F98�جu����;��<��%< )y��������\��o(�c2�6���������~����+��/K���i��6���f��Ď����������cj��~K��+����|(�q䭿+8��d1�x�羃���p�iՄ��Yn��/<L��<�   �   �=|I�<�j�:D�����H�����Րɽ"�ｪ�֕�ܷ���W̽J����wN��z¼��]:��<�s=`�	=��<�Z�h����P*�����ͥ ���C�^ ��H��jf���%���;�և_������-��a��������R������W_�<R;�8���1��1���R8���vB�B���'����(�'T����O���<��=�   �   2E=΂*=\K�<H<�^/������G������ߓ�T����Ɣ�6����K�t��P�@���<�	�<�'(=�TC=�>3=�k�<��P�y4��>�5�┦��m�8O�ʻ����ǿƁ��<"��TF��Sm��E��ha�����0�����Z�����$�l��E��W!�ȫ �Ɇƿ뚒��_M��9�(�����3�9Û��8E����<��4=�   �   �F=Fj1=��<@�\<P`���<ͼR�,�`�d��.������ݹ��mf�BB/�PҼ�;ѻ�V<���<�<1=gF=�h.=D��<4���!��*�L�����E��nXb�tƠ�R�ؿrr�d�0��Y��p��V^�����E=��pͿ��:�����0���%���X�J�/������׿���v'a��(�ݞ��*�K�F.��y�����<��-=�   �   Z�0=��=\^�< �;� ����$���r��-��������ԩ��AD�� wu�>�'����`> ;��<&Y=D1=�& =d��<� ���w���H������B^����!Xտh 
���-��iU����������������w��C������vɖ�t��\�T���,�N�	�#]Կg@���$]��Y�|���nsG������s��H��<"�=�   �   (o�<Pt<`��(z�Ʒt�����������#��|�H��ʺ�;���~x�n���&ϻ0�n<�f�<���<��c<�r��8���J<��A����
��dR�q���+�ʿ�j��$��I���q�k!������g���E��GȪ��מ�/-��ζq�6gI��X$�l �f'ʿ.a��~|Q�6
��t���g;��o��p���kc<P��<�   �    �ܸ�η�z�\��C��2��3-/��cS�/p��i������Z����Nq�O�T�ĺ0�1E��ҽ���`��D���B�X�<�xi;x���Ȑ����)�ә�d����?�ic��텺�o��<c�ZB8��[���}�Pލ��;������^f����L~��K[�:L8��E�O�����I���=?�x���<���)�=휽ȁ���o;� <�   �   p�'��៽��r�9��Pv�u����A���ZȾ�־"�ھ�y־�1ɾ�V��虾��x�n�;�+���2��n�*�����X�L��j��ٍ�nS��e��e�۾�X(�8�r�h�����׿��t<#��S@�hp\���t�����W���ނ��Qu�� ]�H�@��#���5�׿[|��"Or�
(�(=۾T������V����ἐ{H�Q���   �   ڈǽs����g�����nlɾ�A���H�k{��M&�-�)�ţ&�A���Z���˾H���Oj��� �f�ɽ��j�l����������y��O^�`̷�<���!N�d����}���迒}�o$���:��vM��+Z�N�^���Z�b+N�և;�%����+�ֹ��ލ�+5N��������Z�]�����������N ���g��   �   j�/��u������,�/}��|6�H*Q��:f�(�s�a�x��Ht��g��GR�J�7�{��G#��K���Ѡ��Y�1��޽(ȉ�B�M��Gu��L˽�K1��(��2;��(��Ai�י��������@��"���)���2�^06��3�h�)�Hs�"�	�t�뿥�¿@^����i�0s(���N���]1�l,˽��t�t{L�`{���ܽ�   �   D)���Nž��M_/��*Y�f����x��q��\l�������©�2���;�����ݦZ���0�I �#�ƾ<(���e2��9޽}#����{�8��������`�ð���.�7�ku�Қ��XK��\tݿ�����@�b���D��������,����޿�[��rn���5v�ѿ8�����]���na��N�Z����	{��F����ܽ�1��   �   w�¾^i
�%�:��Uo�˸��˓���Uÿr9տ���#��?6�!
ֿ�VĿ���������p���;�a7�ͽþ ���#�#�	�ɽpm��F)���ɽ<�"�8H����¾f
��:��Po�鵒�����6Rÿ�5տڼ�O�俎2῱ֿ�SĿ��������p���;�%5���þ�����#�	�ɽn���,���
ɽ�"��K���   �   ~"���7�u������N���wݿ{����B�����F��������/����޿G^��xp��9v�:�8�n���_���qa��O�^���{��A��w�ܽ�1�+%��~Iž�[/��%Y������u���m��i��`���l���*	��39���}��ƢZ�a�0����B�ƾ~%��Jb2��5޽6"��B�{�B���4�X�`��ǰ��   �   �(��Ei�wٙ�������,��H��
")�&�2��26��3�|�)�u���	���뿪�¿�_��:�i��t(�n�後O��3_1��,˽:�t�zsL��t����ܽ��/�Oq����&� y��w6�,%Q��5f���s�ĝx�)Ct�sg�5CR�C�7��������������1�T�޽)ŉ�B�M��Ku��Q˽�O1��+���?��   �   �$N�l���o���݋�N�q$��:��yM��.Z�
�^�,�Z��-N���;��%�����,鿏׹�����6N����J�����]�]��a����z�*���g��~ǽ����g�M���'fɾ�:���D�!w�I&���)�z�&�<�R����-˾� ��Ij��� ���ɽ�j�x��2��k������^��Ϸ�����   �   T�r�`����׿���,>#��U@��r\�^�t�����˶��]߂��Su��"]���@��#����r�׿F}��qPr��
(�2>۾�������U��$��0\H�x:��"�'��ן�>���9�rGv�-���<��wTȾ0�վ��ھ�s־�+ɾ}Q��u㙾͌x��;�=��\+��b�*��ꖼ��L�n��܍�<V��g����۾C[(��   �   �d���������d��C8��[��}��ߍ�=��J����g�����~�M[�M8�DF�,��_�����c>?� ��=���)�'윽�y��@p;p� < `Ƹ������\��8������%/��[S�_&p�Oe��:������zFq���T�d�0��?�ʽ�,�`�$1�� � ��< �i;����������)�)ՙ������?��   �   ������ʿzk�4�$�p�I�4�q�k"��ѻ��}���N��/ɪ�j؞��-����q��gI�Y$�� ��'ʿOa���|Q�6
�it��g;�+n��0����}c<L��<(~�<�?t<p���fl���t������彇�Z
�����v�S��ر�q���qx�����λ��n<pn�<̈�<��c<�x��;��~M<��C��P�
��fR��   �   ���;Yտ!
���-��jU���������������Ux������ ���ɖ�-t��h�T���,�<�	��\Կ1@���$]�6Y�����hrG�ӎ���l��p�<�=��0=��=�j�<��;T���$��r�m(�����e��ܤ���?���nu�N�'�P����� ;�<2[=81=D& =4��<@'���z��"�H��﴾��D^��   �   Ǡ���ؿ�r�Β0�|�Y��p���^�����_=��pͿ��:��k���/���%����X���/�Z����׿q󟿈&a�2(�ȝ����K�	,��Tr���î<��-=�F=�k1=���<��\<�V���:ͼ��,�Ąd��.����������mf�C/�|
Ҽ�EѻȗV<��<@;1=XeF=�f.=$��<�%��3$����L�������`Yb��   �   ���RXտz 
���-��iU�ޭ��������l���<w���������Ȗ��s��f�T���,���	�\Կ�?���#]�~X����� qG�$���ph��,	�<ޭ=j�0="�=Xk�< �;���$���r�^(�����X��ͤ���?���nu�"�'����� � ;��<�[=�1=<' =��<�"���x��ԀH��2�C^��   �   P�����ʿ^j�ƿ$���I���q�� ������{���>��.Ǫ��֞�0,�� �q��eI��W$�����%ʿ�_���zQ��4
��r���d;��j��𚭼p�c<���<p��<�Bt<P���l�j�t�������z�P
�����v�D�����P��*qx�l����λ��n<�p�<P��<p�c<�p���7�� K<��A����
��dR��   �   �b��L������b�zA8�V
[���}�Cݍ�u:�������d������~��I[��J8�^D�-���������;?�=��o:��)��眽$n���Pp;�� < xøt����\�}8������%/��[S�L&p�He��0�������dFq���T�E�0��?��ɽ�R�`��.�� ( ���< �i;����n����)��ҙ����8�?��   �   �r�{���A�׿<��Z;#�&R@��n\�H�t�*���䳅��܂��Nu�@]�8�@�L�#����َ׿jz��Lr��(��9۾������\P��P��HJH��4��X�'�Tן�	���9�UGv� ����;��nTȾ(�վ��ھws־�+ɾmQ��c㙾��x���;����*��v�*��䖼ȔL�8`�u׍�$R��d��(�۾�W(��   �   ( N�C���t|�����Z|��m$�ܾ:��tM�l)Z���^�ܕZ��(N�~�;�%����%(鿜ӹ��܍��1N�b��a����]���������6s�V���g��}ǽs����g�8���fɾv:���D�w�I&���)�t�&�4�I�����˾� ���Hj�^� �o�ɽ��j���������5v��^��ʷ����   �   (�!?i�fՙ�����7�꿼��V���)�f�2��-6�3��)�q�4�	��뿸�¿�[����i�p(�_�徠J���X1��#˽�vt��kL�wr��
�ܽe�/�*q������%�y��w6�$%Q�~5f���s���x�!Ct�kg�+CR�8�7������ࢹ�t���]�1���޽����M�@u��H˽I1��&���8��   �   ����7�3u�˘���H��pqݿ1����>�T��|B�z������(����޿�X���k��=1v��8�Ν�>Y��aha��I�휦���z�>��0�ܽ1��$��[Iž�	[/��%Y������u���m���h��]���h���'	��.9���}����Z�S�0�����ƾ@%���a2��3޽���"�{�̈́������`������   �   0�¾�c
��:��Lo�����׍��OÿF2տ,��y�俲.��ֿPĿ����ɞ����p�t�;��1��þ%���Ȃ#���ɽ�e��?$��eɽ8�"��G��a�¾f
��:��Po�絒�����6Rÿ�5տؼ�L�俋2῭ֿ�SĿ����������p���;�5�i�þ������#���ɽ�h���$��c�Ƚò"��E���   �   :"��}Ežt���W/��!Y�,���s���j���e�����������6���z����Z��0�%����ƾ&!���[2��+޽���J�{�҄��(����`�@ð���$�7�eu�К��WK��\tݿ�����@�b���D��������,����޿�[��ln���5v���8����U]��na�*M�������z��<��3�ܽq1��   �   ��/��m�����u �u��s6�� Q�m0f��s�!�x��=t��g�>R���7������H�������|1�3�޽5�����M��<u�FI˽~J1�8(��;��(��Ai�י��������@��$���)���2�\06��3�f�)�Fs�"�	�p�뿡�¿=^����i�s(�����M���\1��(˽�zt��jL��o��\�ܽ�   �   �vǽ���<�g�򊝾�`ɾ,4��NA�s��D&�F�)��&���C������˾����,@j��~ �=�ɽ�j�Z��j��\��v��i^� ̷�,���!N�c����}���迒}�o$���:��vM��+Z�N�^���Z�b+N�ԇ;�%����+�ֹ��ލ�5N��������s�]����7����s�r��g��   �   T�'�П�$�F�9��?v�{����6���NȾ��վ��ھ�l־+%ɾ�K��ޙ�a�x��;����� �� �*��͖��tL�dV�[֍�VR�4e��7�۾�X(�6�r�j�����׿��r<#��S@�jp\���t�����W���ނ��Qu�� ]�H�@��#���5�׿Z|��Or�
(��<۾�
�����PS����ἸAH��(���   �    ��Ԝ����\��/��k���/�9TS�5p��`������z����=q���T��0�H9�߾��j�`��� �����<�!j;����O�����)��ҙ�H����?�ic���q��<c�\B8��[���}�Pލ��;������]f����J~��K[�:L8��E�N�����H���=?�X���<���)��ꜽ8s��@[p;�!<�   �   ���<Zt<@v���a�|�t�������彈���
��'q����������`x������λ�o<��<\��<0�c<8i��|6��~J<��A����
��dR�q���,�ʿ�j��$��I���q�k!������f���E��FȪ��מ�--��ζq�6gI��X$�j �f'ʿ-a��z|Q�6
�ot��g;��m�������c<ؖ�<�   �   `�0=D�=�q�<�B ;�䛼��$�ְr��#�������v���]:���du��'�d렼@� ;L��<a=p1=.+ = Š<���w���H������B^����#Xտh 
���-��iU����������������w��C������vɖ�t��\�T���,�N�	�#]Կg@���$]��Y�l���4sG�֏���n����<��=�   �   b9==�(=�:�<�*<x���B���?���x�����?��َ��my�B�@�����
�(�*<���<�|)=d7?=��&=�֛< �ļcNŽ�U��~������i�����j߿��� @6��ba�����#���ǵ��_���
���_���õ�������()a�6�x��߿�}���\i�Q��Dj��_�U�5ƽ��ɼd<�E$=�   �   �'=��
=貚<�t������7�[ヽ�s������Ͼ������ࣽ*c��L�8�$1�� ��ʛ<��=4])=�
=��<� Ƽ���4Q�ֱ��/�B}e�#颿�ۿ�J��3��]�qօ�-l��ʡ������p���� ������e���Ņ�6�\���2���nsۿԱ��6e��
�|���mQ��r½�ʼ ��<��=�   �   ��<�OA<�>�����/�����U��2������ ������{���{[��e܅�|��X��p�C<t��<��<��8<`�˼����D���������UY�G���kѿ�h��*� �P��P{�U#��n���G������P��ͥ�	+��*N{��P���)�,K���пI����#Y�f��������D�a췽��ϼ�r0<�q�<�   �    �m�`@ڼr�m:Ƚ���$.8��x]�w{�����j���7��Ɩ{�G#^�,�8�2�B@ɽb_s��
ۼ@�f�Pq�; =/:p ܼ<��^�1��ٟ�ǅ�(VF��Ѝ��S��o��^1��>��Jc����������AҢ�����o����vkc�:�>�r1��_��N@��򿍿wAF�5���ꟾ�1�ب���߼ �9@|�;�   �   �E;��������;nC��ހ��b������jоkf޾�L�Z�޾��о|=��0�7i��/[D��n	��Ӭ���;�\���t������藽���{ڊ�����5.�߰z�N窿�Q޿����(�3G��d���~�����?��X*���~�^2e��oG���(��,�9l޿��ͼz��?.��㾪������I���TT��f������   �   {�Խ�['��r��s��O�Ѿ������(S"�p^,�B�/�>�,��"�N������ҾI*��St��)(�͹ս��}��F"�* %�����z]��g�|뾾�	�N@U��o����������*�lA�fU��lb�@7g���b�n`U���A�>S*��R��Z�ͻ������]rU�-�k#���
h�����A��B�%�HQ"���|��   �   v�8�Lk���п�E���Y�8H=�u�X��[n��6|�� p|�n�n��DY���=�T��_���e��������9��]�(Փ�`� H���^׽�9�~8�����).��Yq�����CȿkT򿶂�J��d�.���8�Va<���8�X-/��< ������_�ȿQ����q��t.�F[�v����:�_�׽ʘ���`��j��[i��   �   |2��!g;H�3�5�Ra��B��T���{ڥ����	5��w)��� ��]◿����N�a���6�4���-ξ+���״:����w������n����7���j��귾����>�֢}���ĥÿ�����t��,D�d��fd�z���X��Z忖%Ŀ`W��*F~��?��p�6b���zk����"��@ć��.���	꽱�9��   �   ��ʾط��oA�,�w� ԗ�0s����ɿI4ܿ����쿽*迩�ܿ�Lʿ�벿\D����x��B�3+��0˾8p��*�+��ֽ�ݖ�c����zս��*�<�����ʾ���kA��w�'ї��o��N�ɿl0ܿ������&� �ܿ�Iʿ�貿�A���x��B��(��-˾n����+�yֽzޖ�����#�ս��*������   �   k�ɧ>���}����ÿu�� ����lF�����f�p���Z��]�(ĿrY��sI~�(?�hr��d���}k���+�������)��{꽙�9�B.���a;pD���5�3a��?��&���ץ�%����1��%&������ߗ�����a���6�����)ξY���'�:����,���X��������;���j���   �   �,.��]q�N���Fȿ�W򿴄������.���8��c<�9��//��> ����R��u�ȿ�R��U�q��v.��]�򄙾.:���׽����	`��c���_꽴�8��f��9˿�2����T�oC=�/�X�6Vn�1|�
����j|�4�n�@Y���=������������<��g�9��W�ғ�`�-J��pc׽F�9��;������   �   �CU��q��E������:
*��nA�"U��ob�&:g�d�b��bU��A��T*��S��\�R���Ŗ��tU�1.��$��3h���@@���%��F"�@�|��ԽU'�/�r�`n��ѶѾb������N"��Y,���/�҂,�ę"�������B�Ҿ�%��tt��$(���ս�}��B"�� %�����<`���g����   �   �z�O骿=T޿$�t�(�25G���d���~�2��zA���+����~�X4e�qG��(��-�m޿����&�z��@.�6��0������4���VO��V��P���:6;��﫽$��<fC��ـ�H]�������cо�_޾F�̗޾��о�7��b.e���TD��i	�4̬�p�;����ԡ��\��뗽}���܊���Z8.��   �   :ҍ��U��Vq���2�Đ>��Lc� ��}�������Ӣ������������lc�$�>�2��`���@��b���BF�����ꟾ��1��֨��߼ �90��;@�l� #ڼ�r�T/Ƚp���&8��p]��{�P��f��83��h�{��^���8��,�T7ɽ�Qs��ڼ�!f����;�l/:�%ܼo��2�1��۟�f��eXF��   �   ����ѿzi��*�p�P��R{�d$������'H������Q���ͥ��+��O{���P�"�)�bK�#�пk���$Y�b��\����D��귽L�ϼ��0<�}�<�<@vA<������'������ �󽪄����y �o����@���yS���Յ��������C<8��<@�<��8<��˼<��@�D�����#���WY��   �   ꢿ�ۿ�K��3��]�ׅ��l������������\����Fe���Ņ�F�\���2���<sۿ�����5e�K
�ۡ���kQ�
q½�ʼ8��<��=��'=�
=���< ���D��7�Dރ�Yn��	����ɾ�����6ܣ��^���8�H%���~���Л<��=>^)=r
=���<�Ƽ����(7Q�m���+0��~e��   �   �����k߿��p@6� ca�����e��%ȵ��_���
���_���õ���������(a��6��w��߿/}��\i����$i����U��2ƽ��ɼ�ǖ<�G$=&;==�(=l=�<(*<����@���?�V�x�����=��>َ��ny��@�������*<���<{)=�5?=��&=�ћ<��ļ�PŽ��U����A��i��   �   [颿�ۿK��3��]�Vօ��k��s���j������A ��桱�^d��&Ņ�2�\���2��Qrۿ簢��4e��	�٠���jQ�No½��ʼ$��<��=&�'=��
=H��<��������7�5ރ�Mn�������ɾ�����'ܣ��^����8� %��@v��lћ<(�=�^)=h=���<0Ƽԍ���5Q�g���j/��}e��   �   #���+ѿVh�N*�t�P�P{��"������F��﫶�tO���˥��)��bL{���P���)�BJ�a�п���"Y����l�����D��緽اϼ��0<���<�!�<�yA<X����'�������󽞄����y �d����!���WS��}Յ� �������C<x��<��<��8<<~˼�
����D���������UY��   �   TЍ�HS��5n���0�*�>�tIc�������������Т���������^ic���>�0��]���>�����8?F��~�P蟾s�1�aҨ�8�߼ �9���;�l� !ڼr�/ȽP���&8�{p]�t{�F���e��.3��S�{��^�~�8��,�7ɽ�Ps���ڼ�f���;�b0:�ܼ�����1�ٟ�j���UF��   �   ��z�Z檿�P޿����(�~1G�"�d�(�~�9��f>���(��(�~��/e�^mG��(��+��i޿�񪿜�z�9=.��������������<H�xM������^4;����fC��ـ�:]�������cо�_޾F�޾��о�7��Te��{TD��i	��ˬ�z�;� ���Ę��L�T旽L���ي�P���4.��   �   �>U��n��0�������*�jA�U�Hjb�Z4g�Ɣb��]U�~�A�"Q*��P��W�A�������oU��*����[h�i��[:��<�%��A"��|���Խ�T'���r�In����ѾP���ܰ��N"��Y,���/�˂,���"���r���+�Ҿ�%��4t�L$(���ս��}��="���$������[�ŧg��龾l��   �   �'.�Wq� ���Aȿ�Q�$��l��:�.���8��^<��8��*/�x: ���A��^�ȿ�N����q��q.�iV����R:���׽���`�ya��^�4�8��f��˿�����T�fC=�'�X�0Vn��0|�����j|�+�n�
@Y���=��������ܙ����߲9�PV뽗ϓ�8
`�6D��YZ׽d�9��6��5���   �   ��u�>���}��렿:�ÿ���;�~��
B�&��(b�L���V�)W�I"Ŀ�T��dA~��?��m��]��tk����z
�����&��!����9�.��ba;dD���5�*a��?��#���ץ�#����1��!&������ߗ�����a���6�u���)ξ���f�:�7��v������䣱�85��j�跾�   �   #�ʾ#���hA�(�w��Η�m���ɿ�,ܿ�����"�@�ܿ�Eʿr岿�>���x��B�y%�o(˾j���+��ֽ�Ֆ�5���swս��*�����l�ʾp���kA�
�w�$ї��o��M�ɿk0ܿ������&��ܿIʿ�貿�A���x��B��(��-˾�m����+�(ֽTٖ�Υ��_uս^�*������   �   6+��b];�A�a�5��	a�|=��T��� ԥ�����%.���"��g��Xܗ�0�����a� �6����2$ξ᷎�N�:����Jz��/���꣱��6���j�r귾p��>�΢}���åÿ�����r��,D�b��fd�x���X��Z忑%Ŀ[W�� F~��?��p��a���yk�Q�����f����$����2�9��   �   ��8�bc���ƿ�q���dQ�C?=�m�X��Pn�g+|�$����d|���n��:Y���=����~�����������9��L��ȓ�`�aB���Z׽ڬ9�%8�����t).��Yq�����CȿiT򿶂�J��d�.���8�Va<���8�V-/��< ������\�ȿQ����q��t.�[�����:���׽���
`�g^��)X��   �   �Խ�O'��r��i��I�Ѿ����!���J"�lU,��/�7~,�M�"�b�������ҾG ��Y	t�P(�$�սL�}�3"���$�i����[�(�g�9뾾�	�F@U��o����������*�lA�dU��lb�@7g���b�l`U��A�>S*��R��Z�˻������SrU��,�&#���	h�,���<����%��="�R�|��   �   *;�n竽���_C��Հ�nX��
����]оY޾P?���޾.�о�1���蟾U`��tLD�c	�4�����;��|��d���D�:嗽z��%ڊ�g���5.�ܰz�M窿�Q޿����(�3G��d���~�����?��W*���~�^2e��oG���(��,�9l޿��ȼz��?.����T������ʛ���I�I��H쳼�   �   �Il��ڼ,�q�(&Ƚ���8��h]� {��	��Za���.��[�{�I^���8�F&��+ɽZ>s�h�ڼ`Pe�@��; �1:dܼ�����1�Nٟ����"VF��Ѝ��S��o��`1��>��Jc����������BҢ�����n����vkc�:�>�r1��_��N@��򿍿pAF�&���ꟾH�1��ը�x�߼ `�9���;�   �   )�<`�A<���F��� ���y���������t ����<���y���I��+ͅ��x��|���C<<��<"�<��8<�v˼�	��.�D���������UY�F���lѿ�h��*� �P��P{�U#��n���G������P��ͥ�	+��*N{��P���)�,K���пG����#Y�[��`��� �D��귽�ϼ��0<̄�<�   �   �'=��
=�ƚ< (缼��7�ڃ��i��گ��/ľ�@﷽�֣��Y����8���@���(ޛ<��=pc)=l=䊌<�ż�����4Q�ı��/�A}e�#颿�ۿ�J��3��]�qօ�,l��ʡ������p���� ������e���Ņ�6�\���2���nsۿӱ��6e��
�k����lQ�r½\�ʼ���<p�=�   �   xf?=FF*=���<`�3<�l�`���<��Yu�W��쒽e���N�t��;�����d
�8�<<,H�<*�-=~AC=��*= �<��i����JS�zｾ�M9h��Ǥ��3޿6��tH5�~+`�� ���4���ݴ�Up������s�����dN���&����`���5��6��޿�2����h�h���侾��T�6�Ľp�ļ;�<�s&=�   �   �)=��=�T�< tй0����5�M������b���J���ŏ���V��΁���3�H_�� �9��<�=j~-=�H=�Ǖ< )���'��*�N��*��%#�}d������ڿ���(2���[��#��᝜���������������Ȱ�����`C���5\��x2�����ۿ�c����d������\�P����|�ż4-�<�=�   �   ���<�J<�w��#�tÃ������񽰄����.�|��hZ��|�<\�����,?����V<<h�<���<8�K<�����ó��B�(L��B���X��ۙ�п����7)���O�~'z�"u��v���xq��,ʵ�j������~w���Ez��P�fr)����lпK6����X�<��-���D�������ʼ��9<t�<�   �    4F�D,ռlo��ƽF��X?7�c\���y�
U��ڑ��I����y��)\���6��i�A�Ž�m�`{м@�� V<@��:��Ѽ8褽ԫ/�����k��y1E�#���n���^������=� mb�{���a��8�����t)��SM��=l��Zgb���=�,��7�������p`����E�_��W���1�c���pڼ Zh:0��;�   �   ��8�ډ�����b�B��`���Ξ����A�ϾSjݾ�)�b[ݾO|Ͼ蹾����=���DB�ɜ�|���$g6�����Ȯo�`���������������c��?-��|y��.��\}ݿܜ
�&(��F�<4d���}�����~����x��y}�� d�<|F�2(���
�a�ݿ:f����y���-�M'㾞d��F���P���|������   �   })ӽC�&��r��룾6Ѿ�4���B���!�6�+�[/�	�+���!��,�'
��n�о�ˣ�_�q�};&�E|ҽ*x�d$�`�������� �I�e������B�-LT�@���9᾿#X�b��R�)���@��}T���a�J@f�d�a�FT���@�nz)�B���T����������T�Õ�	L����f���̟��T�"��\���y��   �   ��7�Pሾ�6��D3�������<��,X��m�t[{�x���H{�X�m��X��<�;��(��_#���҈��7��5����
[�~�����Խn8�;��ۺ�n-�h�p������ǿF��<�D��@~.�H8�L�;��+8�P.��i��T��D�ǿ[�����p�(�-��1����r�8�u�ս�ׂ�h�\�o�������   �   ؒ����̾����5�f�`�����0��	l��x��Ќ��*h��Q�����߄�Ko`�Ap5�s��X�̾������8��������{U��\8������Hi�V�������>�&�|�g���ACÿb俦� ��e����Bd����2D�P� �I%��ÿP~��k�|��>����I��?�i�[������؅�nG��Q���8��   �   ͸ɾm?���@�#Rw�ޅ�����,qɿ�ۿL�=@��1���ۿ@ɿ"񱿽h��Q5w�H�@�QJ�H�ɾ#p��N�)�k�ӽk�������=ӽ�)��E����ɾ<���@�Mw�肗�Z���mɿ1�ۿH�N<�.�yۿ�<ɿYaf��o1w�7�@�H��ɾ�m����)�N�ӽ�������uCӽ�)��I���   �   m���>���|�9����Fÿ�e俬� ��g���|f����&F�� �K(�kÿb�����|�n>�̲��K���i�X\�����Mօ�NB���罶�8�����g�̾�����5�F�`�����,���h���t��b����d���M������܄�k`��l5����[�̾ʘ��L�8���罡����V���<������Ni�� ���   �   Aq-�x�p�������ǿ���>�~����.��J8�֭;�&.8�:R.�pk�����[�ǿ���{�p���-�k4������8���ս�Ղ�P�\�ǲ��<��.�7��܈�01��4,�������<��'X�s�m��U{����'C{�"�m�X���<����~�����qψ�|�7��/����	[�������Խ�8�V>������   �   nOT�S⑿�㾿)[�,��l�)�"�@���T�|�a�*Cf��a�rHT���@�|)�����V�l������)�T���jM�� �f�T��z�����"�R���y�ӽ\y&���q�,棾�Ѿ=-���>�I�!���+��/���+���!��(������оWǣ���q�j6&�2uҽXx�P ����T ��L� �Ӽe�����AE��   �   �y��0���ݿT�
��'(�H�F��6d���}��������z��t{}��d��}F�T (���
���ݿ-g��*�y���-�c(�%e��}���<��P�{������x8����>��h�B��[��:ɞ������Ͼ�cݾ�"��Tݾ6vϾ�⹾����9��>B��������\6�8��x�o����������������-g�ZB-��   �   ����p���`��H����=�ob�U|��c���9��S
���*��mN��m���hb���=�г�"��������`��?�E����W���1��a��Dhڼ �i:�4�;�}E�ռ�Yo��ƽ����77��Z\���y�kP��<����D��@�y�R"\��6�0d�^�Ž0tm�gм`�� e<���:ЫѼb뤽��/�Ŏ�����3E��   �   �ܙ��п����8)�@�O�F)z�-v�������r��=˵�k��S���x���Fz�FP��r)���Qlпp6��¢X�<��-��D�$���4�ʼ�9<��<$��<h�J<�H�d�+���D콽���'�i��)���RU��s�DT������^4�X���/V<�o�<@��<�K<�����Ƴ���B�N������
X��   �   �����ڿ����)2���[��$������c°�c��-���K��cȰ�Ͱ��{C���5\��x2����ۿ�c���d����u��L�P����t�żL4�<�=��)=R�=�a�< �̹8��� �4��G������ﷵ�䑼�����R���Ɂ�x�3��S�� N9���<�=h-=`H=�ĕ<�/���*��R�N�X,��A$��d��   �   ?Ȥ�84޿����H5��+`�+��.5��#޴�op�����s�����$N���&���`�6�5�:6�A�޿L2����h�����㾾�T���Ľ��ļ\@�<v&=Jh?=�G*=���<��3<h�@���<�0Yu�-��쒽�����t�ش;�����i
��<<LE�<��-=�?C=x�*=��<�������tLS�����B:h��   �   P���ڿ ���(2���[��#������Z���I�����1��Xǰ�䯜��B���4\��w2����ۿ�b��	�d�ݮ�q����P������żX7�<t=F�)=��=hb�< �̹Э����4��G������ڷ��ؑ������R���Ɂ�^�3�8S�� �9H��<8=�-=DI=�Ǖ<H+���(����N�T+���#��d��   �   wۙ��п���x7)�J�O��&z��t�������p��ɵ��h��e���qv���Cz�LP�Fq)�����jп5����X��:��+��~D�ׂ����ʼ@�9<X�<���<��J<0F�������콽����\���(����DU�}s�#T�������3�(���2V<Dr�<���<�K<4����ó��B�0L��:���X��   �   ���7n���]��L���=��kb�7z���`���6��~���'���K���j��Deb�(�=�ұ����'����^��r�E���GU��1�I]��`\ڼ��j:I�;�cE��ռ�Xo���ƽ����77��Z\���y�bP��2����D��.�y�<"\���6�d��Žtsm��dм f� o< J�:�Ѽ�椽"�/�������0E��   �   {y��-��|ݿ�
��$(���F�D2d�<�}���������w��v}�b�c�zF�j(�@�
��ݿ;d����y�3�-��#��a��L������ ����{�ġ���v8��~����8�B��[��'ɞ������Ͼ�cݾ�"��Tݾ*vϾs⹾�����8���=B����^����Z6�dy����o�����b���R��ѵ��}b�?-��   �   {JT�ߑ��߾�,V�"����)���@��{T��a�h=f�~~a�\CT�(�@�Tx)�x���Q�\������5�T�D��XH��J�f�ʸ�����6�"�M�|�y��ӽy&�x�q�棾�Ѿ(-���>�B�!���+��/���+���!��(������о@ǣ�I�q�6&�2tҽ2	x�Z�*��t����� ���e�䮽��A��   �   ?l-��}p�j�����ǿ���,;�d��|.��E8���;�2)8��M.�Xg��٠�G�ǿב���p��-�$-�x����8���ս�ς�x�\�?�����车�7��܈�1��,�������<��'X�k�m��U{���� C{��m�X���<����j�����Hψ���7�(.�[��T[�����v�Խ�
8�C9��<���   �   ���T�=���|�O����@ÿ_��� ��c����b����
B�J� ��!俜ÿz{����|�>���	E����i��U��ﯽ�Ѕ��>�������8�f���>�̾}����5�;�`�����,���h���t��^����d���M������܄�k`��l5����5�̾������8�I������)Q���3��<��#Ei������   �   E�ɾ�9���@�Iw��������Xjɿ��ۿSD�]8�#*翝{ۿ49ɿ 뱿fc��P,w���@��D���ɾ�i����)���ӽ��������9ӽ�)��E����ɾ<���@�Mw�゗�W���mɿ/�ۿH�K<�.�uۿ�<ɿV]f��g1w�.�@��G���ɾ�m����)��ӽٞ��$����7ӽ��)�nC���   �   ����B�̾���$}5��`���*���e��Wq��񅱿ea���J������ل��e`�rh5�+����̾W���~�8���������N���3������Gi����r���>��|�b���=Cÿb俥� ��e����Bd����2D�N� �F%��ÿL~��c�|��>���@I��_�i��Y�����х�K=�����J�8��   �   �7�fو��,��r&��-����<��"X�5�m�P{�d��\={�~m���W��<����Y�����ʈ�:�7�e$轲��*�Z�ĸ���Խ?8��:�����n-�_�p������ǿB��<�B��@~.�H8�J�;��+8�P.��i��Q��C�ǿY�����p��-��1����D�8���ս�т�|�\�4���Ǎ��   �   �ӽ�s&���q��᣾1Ѿ�&���:�#�!�8�+�5/��+�#�!��$�&���j�о����x�q�'/&��iҽ��w���������� �\�e�B����B�#LT�?���8᾿ X�b��R�)���@��}T���a�J@f�d�a�FT���@�nz)�B���T��������v�T�����K����f����8�����"�I���y��   �   �l8�tw�������B��W��`Ğ�L�����Ͼ]ݾ��Nݾ�oϾdܹ�8���54���5B�������"K6�b�� so�����K������V����c��?-��|y��.��[}ݿܜ
�&(��F�<4d���}�����~����x��y}�� d�<|F�2(���
�b�ݿ:f����y���-�'�Hd��0���������{������   �   ��D�t�Լ(Ko�˰ƽ��017�(S\�_�y��K�������?��C�y��\�}�6��]���Ž$am��Gм�����<��:ȗѼ�夽�/�U���\��s1E�!���n���^������=� mb�{���a��8�����s)��QM��=l��Zgb���=�,��9�������o`����E�P�|W���1��`���aڼ k:Pf�;�   �   ��<��J<�$�$
�R���'佽e��z���R#�H���O�%i�J�����%�����YV<���<��<@�K<����³���B�L��9���X��ۙ�п����7)���O�~'z�!u��u���yq��,ʵ�j������~w���Ez��P�fr)����lпM6����X�<��-��D�������ʼ��9<��<�   �   6�)=��=�h�< Yʹ<�����4��C��壡�����y���,����L���ā��3�PB�� �9��<�=��-=PM=�Ε<<$���&����N��*��!#�|d������ڿ���(2���[��#��������������������Ȱ�����`C���5\��x2�����ۿ�c����d�������P������ż�3�<*=�   �   HL=f�7=lX=�Qx<�4������$�&�Z�C}��`����{��>X�j� ��N��@=C���<j�	=Z�==@�R=,;=�q�<���4���F������q.^�����wտ�E
�:�-��*V�l`��j����}�����h�����������1��
���d�V�ά.�`���ֿ�
����_�"�����>I��D���Ù��t�<�3=�   �   n!7=$=Ȏ�<���;Č�d��6vi�J���#-��/�������߼��� f��������0��;8{�<�!=��==��,=@��<Ո�Tu��T�A�p~����@4Z��^����ѿT
�V�*��7R��x}�P���Л��QU��ĸ�S�������ʔ��~���R�Ψ+�^���$ӿO��z�[�KF�Kb���E�֚�������߬<��%=�   �   �o�<�d�<0 ��l���hl��i������4������>��V��޽08��8�g�����E2���<���<�|=��<8�������6����3�W�N�����6�ǿ��Ѓ"��G���n�7�������L��g���7��nw��5��N�n��kG�R#�>���ȿ)[����O��	��ϧ���8��X���L���-~<ȁ�<�   �    ��:D*��~U�����a�jk,��-P��ll�u~�%A��^�}���k��O�� +�v��6��T�O�XΝ�`�G;��U<��;�S��&Z���#����;�����<�uH���𷿸��֙��,6�b�X���z�Y%���<����f�����dRz��qX��A6�������ٖ���⇿�=���������|&�<����]��0°;��<<�   �   �������Ǫ��ji7�-bs����o4��J�žUӾ��׾��ҾsRž�u���0��z�q���5�[����ᘽ����q�����ļF1�������=j׾/�%�L!o�d~���տ�p��!���>��dZ�,$r����3��D����q���Y��1>���!�$q�]տWۣ���o��R&�S�ؾ�E���,��Ո���Ѽ��)�(߃��   �   �½(G�.e�>�����Ǿ1�����j]$�ƍ'�#$�4t��n�����ƾ�
����c����X���6Z�������D�q��$��OX�5��΢��XK����n������l��B#��]9�ֶK���W��\���W��K�B�8�`�"�&��8�g����4��H�K�I �O-���Z��[��w�"�
�"����^��   �   =-��ہ�&H����jM�5��vO��$d��Dq�w�u�|�p���c��N�JP4�ƙ�/�ﾻZ��+$���+�S�ս������>��5f�+ý8�,��A��2��Q�%���f��q���a�����"����f�'��1��(4���0�RS'���d��kM��꿿�<��=�f��&�.⾦א�0�-�PBŽ�0j�r�B�2����v׽�   �   aP��6þF���
.���W���?l��%���ѧ�k���@��������㐿�~��V�O-��M��|¾�ԅ�R'-�G�ս���d�m�0R��X�[)\�.��v�T6��r�9{��`���(ܿ9d���J��]�*��������f���>ۿAc��}����^r�O�5�6s��(���\���m��&�o����� �ֽ�-��   �   �8��n	�K�8���m�|Ǒ�Ʉ���¿B�ӿ��޿1s��g޿�ӿ&U��w̪�.����l��g8�ի�῾�~�R���j½�Ӆ�Hυ�Ug½c��\~�4��7��:�8�Ԗm��đ�����a¿��ӿ.�޿ho�&d޿_ӿR���ɪ��+����l��d8�����ݿ��~�����h½{ԅ�v҅�im½8��c~��   �   @���6���r��}������,ܿh���L� `�L�������Gj��oAۿ�e��� ���ar���5��t�!+����\�\��m��X�o����� �ֽ2�-�RL���0þ���W.���W����-i���!��nΧ�����������ᐿ-�~���V��K-�K��x¾�х��#-�L�ս�����m�%V���	��.\�<
���   �   Z�%���f�`t���d��)��$�Լ���'�1�P+4�B�0�^U'�� ����O��쿿->����f��&�p0�ِ���-��BŽ4-j���B��}��Om׽��,�Gׁ��B����_I�r5�zqO�kd��>q��u��p���c���N�OL4�l�����V��!����+���ս������>�r9f��ýG�,��D������   �   \K����ᦷ����|n��D#��_9�b�K���W��\��W�K��8��"�Z��:�⛷�6����K�_!��.���Z�w\�J}w���
��v�>�^���½}@�}%e�����m�Ǿ������Y$�a�'��$�:p�&k�����}ƾ}���c�.���Q��,.Z������N�q��)�5TX�f8��#���   �   [$o�O���� տ*r���!���>�\gZ��&r�;!���������q���Y�N3>��!��q�\^տCܣ��o��S&�^�ؾ0F��-��Ԉ�̤ѼXp)��ȃ��������-����a7�Ys�y����.���ž�Ӿ�׾_�Ҿ�Lž@p���+����q�D�5������ژ� v��|q�����ļ,4��\����m׾��%��   �   �I������� ��X.6�P�X���z��&��B>��ę�������Tz��rX��B6�r����{���ㇿx�=�%���R����|&�����U����; �<<@\�:����U�T򶽐[�.d,��%P�,dl�'l~��<����}���k��O��+�* �;.���xO�����`DH;��U<p��;�X��5]����#��
��T�����<��   �   (�����ǿ�����"��G�T�n� 8������M��h���8��.x���5���n�0lG��#�t�5�ȿN[����O��	��ϧ��8�wW��lE��(@~<���<�~�<�w�<𣄻��Xl�{`����|����Y��;9� R�,�޽�0��R�g��n鼀�1�t�<��< ~=��<,��������6�o����*�N��   �   h_����ѿ�
��*��8R�z}�����{����U���ĸ�uS��榧��ʔ��~���R�Ȩ+�N���$ӿ�N���[��E��a���E�
���Ȍ����<��%=�%7=X)=H��< /�;����@��^li���'������
��]����f�Ґ�$�����;���<!=��==��,=��<�ۈ�x��f�A������5Z��   �   ]��axտ,F
���-�8+V��`������"~��+���h������}���Q1��˶����V�h�.����ֿ2
����_�h����X=I��B��(����y�< �3=!L=�7=�Y= Wx<�*������ $�z�Z��B}��`��,�{�N?X�2� ��P��@PC�$�<��	=ؚ==��R=0;=�l�<����r��F�������^/^��   �   �^����ѿf
�`�*��7R��x}���������T��{ø�cR��饧��ɔ��~���R��+�����#ӿ3N���[�4E��`��fE�V���`�����<��%=�&7=�)= ��<p1�; �����0li�	��'��슬���O���nf����䪃���;��<r!=R�==t�,=ؐ�<(׈�Yv���A��~��S��4Z��   �   ێ����ǿ��~�"�G��n�y6��A����K���e���6��\v�� 4����n�RjG�<#�^�~�ȿ�Y����O��	��ͧ���8�BT��=��0K~<L��<@��<0y�<𞄻 ��HXl�O`����n����H��.9��Q��޽]0���g��m� �1���<l��<�=��<���`��� 6����.�;�N��   �   	H��,����<���+6�2�X��z�R$���;��`���	��6��Pz��oX�&@6����|�����=ᇿ=�Q�������ly&�����(J����;(�<<���:����U���h[�
d,��%P�dl�l~��<����}�r�k�vO��+� ��-��LxO�����`]H;(�U<���;�M���X��j�#��������<��   �   �o�y}��Vտ�o�ع!�J�>�"cZ��!r�{���������q�`�Y��/>�F�!��o��Zտg٣���o�xP&���ؾC���(�Eψ�ܖѼ ^)���������������a7��Xs�g����.����ž�Ӿ�׾R�Ҿ�Lž3p���+����q� �5�:���ژ�Vt��qq����L�ļ�.��S�
��i׾I�%��   �   YWK��������,�濒k�JA#��[9���K�j�W�.\�؊W�LK���8�b�"�p��5�򗷿�2���K����)��ZZ��S��qw�f�
�r���^���½@�6%e�����P�Ǿ��������X$�X�'��$�3p�k����}ƾh��͆c�����P��(+Z�ޡ�����q�-!MX��3������   �   ��%�#�f�Yp���_��Q�z!���X�'�Z1��&4���0�Q'���|��J�迿&:��I�f��&�l)�.Ԑ���-��9Ž�!j��B�@{���k׽2�,�ׁ�zB����PI�f5�pqO�bd��>q�ޡu��p���c���N�FL4�b�����eV��� ��(�+� �ս"���0�>��-f�ý�,�@������   �   �}��6���r�5y�����&ܿ�`���H��[��������c���:ۿ`�������Yr���5�Yp��$��h�\����d��<�o�����Ŭֽn�-�L��s0þ���G.���W�t��(i���!��iΧ����	�������ᐿ$�~��V��K-��J��x¾�х�#-��ս*����m��M�����%\�����   �   �0�����8�8��m�M��~��G¿�ӿ��޿�k�S`޿��ҿ�N���ƪ��(���l��`8�W���ؿ�~���v_½A̅�6ʅ�d½V�\~��3��#��*�8�Ȗm��đ�����]¿��ӿ*�޿do�$d޿[ӿR���ɪ��+����l��d8�����ݿ�~�����e½�υ��ʅ�b½�	��W~��   �   ^I���,þ2���.�~�W����of�����4˧�ŭ�����������ݐ���~��V�G-��G�ws¾�ͅ�2-��ս%����m��M����o(\����`�B6���r�3{��Y���(ܿ5d��~J��]�(��������f���>ۿ>c��}����^r�E�5�"s��(���\�����h���o�ǟ��ֽۨ��-��   �   ��,��Ӂ�>>��B��E�i5��lO�Wd��9q�N�u���p�!�c�p�N��G4�[������P�������+��xս����<�>�j*f�|ý�,�zA�����@�%���f��q���a�����"����d�'��1��(4���0�PS'���b��jM��꿿�<��9�f��&��-�Pא�
�-��>Ž�%j��B�Yx��f׽�   �   #�½:;��e����Ǿ����������T$��'�[$��k�'g�z��twƾ*��Q~c�2���F��nZ�ȗ�Vy�Z�q��!��NX��4������XK����k������l��B#��]9�ԶK���W��\���W��K�B�8�`�"�(��8�h����4��A�K�8 �-���Z�Y��vw��
�Bn���^��   �   ���қ������>[7�Qs�����7)���ž�Ӿ��׾׾ҾGFž^j���&��z�q�m�5�����И�e��Dq���l�ļ�-�������j׾$�%�F!o�c~���տ�p��!���>��dZ�*$r����2��C����q���Y��1>���!�$q�]տYۣ���o��R&�'�ؾ\E���+�D҈�H�Ѽ�U)�𶃼�   �    e�:�����T�c鶽V��],��P�\l�wc~�68����}��k�x�N�]+����B#���fO�@��� I;x�U<��;PE���W��R�#�W�������<�sH���𷿸��֙��,6�b�X���z�X%���<����g�����dRz��qX��A6�������ږ���⇿�=�p���ކ��*|&�Ѥ��XO����;`�<<�   �   l��<Ą�<p^�� ��jKl��X��zགྷ��`������3��L��޽R'��yg��R� 1��&�<\��<ą=0��<В�������6�l��+�R�N�����7�ǿ��Ѓ"��G���n�7�������L��g���7��ow��5��N�n��kG�R#�@���ȿ+[����O��	��ϧ�"�8�LW��C���H~<h��<�   �   z'7=�+=X��<�T�;����8��di��쒽�"�������y�� ����f���������X�;���<�!===H�,=䗼<\Ј��t���A�`~����>4Z��^����ѿT
�V�*��7R��x}�O���ϛ��RU��ĸ�S�������ʔ��~���R�Ψ+�^���$ӿO��y�[�FF�;b��~E���� ���T�<p�%=�   �   L�a=�eN=!=,�<0��;0�[�d����*���J�>U���H�$�&�� ���>�@��;��<��'=�X=yl=8UV=V$=@�ƻ�?���7/�N����R�g�L��,��Mƿ�k ��!�H&E��Il������!ئ�I����ަ�";���&��.$m�1F� "��h��ǿ���a�N���P����3�^������ ��<��J=�   �   ��M=��3=���<��F<0�8�B�8�4Iq��m���#��r=��H�l���2��FӼ ^��80k<:h=��==:�X=�I=X8�<�z˻�����`+�.��������H�꬏���¿<����h���A���g���������������}��e���S*���eh���B��^�F����iĿ��� �J��i��S����/�8����J����<��==�   �   �X=���<���;d����;��l��4�����S;��jd������y�_ҽ�i����2�dM�����;���<f�=�
 =��< ��Jф�<\ ���������>��d���f��k������7�*�Z���}�����P�����A6��؍�x�}��[�HK8�@u�o&򿤬���}��P�?� ���s��z$�닽$��ں<�=�   �   �= <6�P�%�I~����潨���	:�@T���d�mZj�Xd���R��8��p�5���o��p�������H<�ΰ<P��<���Ԅo�!��l#��qLᾥ@-���y�����	޿� �D�(��G�*ye��M��q��W���?��$�~�p e��LG�n�(��M�s�޿ti��u�{�ֱ.���j=���?��:|��@��Z<p8�<�   �   �,��뀽��ܽ�#���Z������:L��6����ľg����S��Qԟ�.T���X��9 ��'׽d�w���Լ,�� �i:`�Y�2�S������Ni��	ľ�����\�r����ſ)7���;�p0��2I��^��l���p���k�"I]�<kH���/�`��+��SGƿ�痿�]������ž~�l�H���؂^�8񀼀+�� �߻�   �   �w���	�P�M��n��:��$�ݾ@a �_;�������e�����۾n0�� Ë�(�J��!�T⠽��&�\쩼�ӯ��[=�f8̽˹@�	h��ڝ��X>;� ����p���kֿ��>��(�+�b3<� �F�<�J��|F�B_;���*�<��z>���տ]R��گ��]�;�Nl �����&C���н��E�/��T,��L�.��   �   .A�j��䥾�ܾl���&��e?���R���^�<�b�W^�x�Q��7>�{�%���	��ھ�<��log�������M� E��63�yf��P"������;�l�w�T��<������ؿ�x��r�����
:$�.�&���#��-��'�������׿|��ߌ���T�G��icξ^Ƃ�ߣ��l��J39�&Q�GT������   �   NBr�ݱ�2e���7 ��G�Ήl�ͼ������/���TH��mF��]蒿�셿��j��E�M��f��愰�^Xp����(�����]�n�:��Z���+彠�D�f蝾���'���`��7���ˮ�Q�̿W?�����0q�����������]�˿z���'s���_�J'���z坾�$E��j�m҄��>�jNa�$�������   �   �����3���b*�h�[����s>��e��'�Ŀe)Ͽ��ҿo�ο��ÿ�K��)��*��R0Z�d)������8����c�ԑ�"��pW� �W��~�������d�����-���^*�̘[�C��k;���a����Ŀ�%Ͽ�ҿ�ο��ÿ�H���&���'���,Z�_a)������5����c����8 ��&qW��W���������d��   �   ���'�"�`��:���ή���̿�B�����*s������������˿Ÿ��u����_��'�A�쾠睾>'E��l�x҄� >�Ea��������:r�ر��^���3 ��G���l�칆�ꍓ����9E��mC���咿�酿��j��E�;�����R���NSp�?~�v���Z�]���:�p^��I2���D�-읾�   �   �o��T�=?��ʿ��2�ؿ9|��f����8<$�X�&���#��/��)�m���,�׿`��������T����eξ�ǂ�-��Um��09��I� ;T�����;��j��ߥ���ܾ��
���&��`?�r�R���^��b��Q^�ķQ��3>�Ƈ%���	���ھ�8���ig��������M�D�n:3��j��&�}����;�   �   EA;������r��Knֿ�����8�+��5<�d G���J��~F�:a;���*�����?�`�տ�S��氁���;�Rm �ج��V'C�x�н6�E��#��T��p�.�n����	�\�M��i��g���t�ݾ�] �h7�z����������Z���۾�+������J�8��۠���&��䩼Lԯ��`=�I=̽ڽ@�k��0����   �   ��\��s��- ƿ�9��=��q0��4I��^�rl�
�p�ؚk� K]��lH�,�/�`���,��Hƿ�藿��]�o����žp�l�����̀^��瀼@?��0{߻ 輆‽�{ܽ�
#��Z���T��bF��*z���~ľ��N��eϟ��O����W��3 ��׽�w�X�Լ������j:X�Y���S������Ri��ľ����   �   �y�#����޿����(���G�.{e��O�s�������@���~��e��MG�6�(��N�H�޿j��D�{�Y�.���㾢=���?��8|���?�X5Z<DH�<Pg <��5���%�8t�������5:�8T���d�$Rj�Zd�D�R��8��j�U���g���������H<Tհ<���<���r�o����`%��OOᾣB-��   �   �e��9h��	�����7���Z�8�}������Q�����7���؍�v�}��	[��K8��u��&�⬺��}��k�?������r���y$��鋽X�#���<4"=�_=\��<`��;�����;�|d���*�����1��M_�����p�ʽ��a����2��9��p�;x�<��=, =��<���Ԅ��^ �����2����>��   �   ������¿l����i�̭A���g�p���+���/��`����������*���eh���B��^�'����iĿ������J�~i�mS����/�����p=�X��<��==4�M=��3=t��<�G<8� ����8�x?q��h������8����l�j�2�:Ӽ�3���@k<:k=��==(�X=�I=D5�<p�˻J����b+���������H��   �   c-���ƿ�k �P!��&E�HJl�7����7ئ�J����ަ��:��q&���#m��0F��"�2h�z�ǿ������N��M�����3�7������$��<��J=�a=hgN=�"=��<���;��[����D�*�F�J�>U��H���&�\���>��|�;,�<D�'=x�X=twl=XSV=�!=�ƻ�A��9/�P���PS�B�L��   �   �����¿b����h��A���g�����N���:��c���
��˸���)���dh�̑B�,^�����hĿ;�����J��h��R��s�/�����(5���<��==��M=��3=,��<�G<@� �� ���8�T?q��h������8����l�J�2��9Ӽ�2���Ak<�k=J�==��X=�I=8�<p�˻����Va+��������H��   �   cd���f����F��n�7�|�Z���}�`���O�����K5��׍���}��[�J8�Bt��$�F���h|����?�f���,q��Bw$��拽`�#���<�#=�`=0��<��;|��(�;�Id���*������0��>_�����dp� ʽ��a��|�2�9��@"�;��<��=� =� �<p�� ф�>\ ����������>��   �   ��y�����:޿6 ���(��~G��we��K��p��-~���>��ܹ~�f�d��JG���(��L�u�޿�g��Ѓ{�ϯ.���6;���<�40|�p�?�0DZ<4M�<n <��5���%��s����潼��:��7T���d�Rj�Bd�/�R��8��j�%�Ὑg��&��X����H<�ٰ<x��<���J�o�|���"���K�!@-��   �   y�\�0q����ſ�5���:��n0�21I��^��l��p�
�k��F]�iH��/����u(��Eƿ旿��]�h����ž��l������v^��ڀ������c߻��ွZ{ܽW
#���Z�ֽ��?��PF��z���~ľ��N��Yϟ��O����W��3 �Z׽άw���Լ@ꓻ��k:��Y���S�i���Mi��ľ����   �   �<;����-o���iֻֿ�޴�z�+�f1<���F�ږJ�8zF��\;���*�h���<���տP������d�;�j �E���$!C�1�нJ�E�������@�.��l��M�	��M��i��I���V�ݾ}] �^7�p���������J���۾{+������ξJ���۠��&��۩�TƯ��U=�!5̽��@��f�������   �   /k�,�T�x;��0�����ؿ�u���������7$� �&���#��+��%������׿����܌�ԽT�d��_ξ!Â����d���$9�hB�"6T�@����:��j�zߥ�q�ܾ��
�t�&��`?�f�R���^���b��Q^���Q��3>���%�~�	��ھ�8��Eig��E���z�M��<��/3��b�������D�;�   �   /	�9�'��~`�6��_ɮ���̿2<�|���Jo������4���I��	�˿�����p����_��'����s᝾�E�$a�ʄ�|�=�>a�\���I��;:r��ױ��^���3 ��G�~�l�幆�䍓�	���4E��jC���咿�酿��j��E�3�����2����Rp��}�L�����]�j�:��V���&�8�D�松�   �   �񮾏)��\*�;�[����8���^��s�Ŀb"Ͽu}ҿs�ο�ÿ�E���#��=%��3(Z��])������0����c���b���aW�t�W��{�����F�d������-���^*���[�;��e;���a����Ŀ�%Ͽ�ҿ�ο��ÿ�H���&���'���,Z�Ua)�����q5��V�c����%���gW���W��y��F��q�d��   �   65r�SԱ��Y���0 �G��l�X���������B��K@���Ⓙ煿L�j�}�E�J��!�-|��UKp�x�ǈ��*�]�ʾ:��V���(彼�D�蝾Z�s�'�ρ`��7���ˮ�K�̿Q?�����,q������������Z�˿x���$s����_�A'���>坾�#E��g�[΄��=��;a��������   �   z6��j��ۥ�_�ܾt�
���&�{\?���R���^���b��L^���Q��.>�q�%���	���ھj3��9ag��u�`�M�z5�8,3��b��,!�=��i�;�l�h�T��<�����
�ؿ�x��n�����:$�,�&���#��-��'�������׿{��
ߌ���T�<��;cξƂ�Ȣ�}i���(9��A��0T�����   �   �f��Ū	��M��e��f�����ݾ$Z ��3�y�����נ��������d�۾�%������J����Ѡ��q&��ȩ�����xS=��5̽�@��g������L>;�����p���kֿ��:��$�+�^3<���F�<�J��|F�@_;���*�:��{>���տ[R��ٯ��W�;�>l �^���@%C�:�н.�E������n�.��   �   ���ۀ�Hrܽ�#���Z�����P���@��At���xľy쿾:H���ɟ��J�� �W��, ��׽0�w�T�Լ�����hm:X�Y���S�����Ni��	ľ�����\�	r����ſ$7���;�p0��2I��^��l���p���k�"I]�<kH���/�`��+��UGƿ�痿}�]������ž�l�<���X|^��݀��t��08߻�   �   �� <`�5�Z�%��k�������V�9��0T���d��Ij��d�3�R�@�7��c�]�Ὕ]�����y���H<��<���<���*�o�b��0#��PLᾝ@-��y�����޿� �B�(��G�*ye��M��q��W���?��"�~�p e��LG�l�(� N�s�޿ui��v�{�ұ.����6=��&?�6|�8�?� FZ<�S�<�   �   Td=���<�>�;�&�;�!]��Q"�����'��$Z�[���}f㽺���FY����2����Px�;��<��=\ =h)�<`���τ��[ ���������>��d���f��i������7�(�Z���}�����P�����A6��؍�v�}��[�JK8�@u�p&򿦬���}��P�?�����r���y$��鋽�#���<`%=�   �   ��M=ܟ3=��<HG<�� ����N�8��6q�-d������3���l��2��(Ӽ ���@\k<Pq=D�==��X=I=t>�<Pi˻���b`+���������H�꬏���¿>����h���A���g���������������}��e���S*���eh���B��^�G����iĿ�����J��i��S��i�/�{����A����<P�==�   �   t�|=@jk=lp?=zU=�o�< �����r�4ռX/���ĕ���Ǽ�|L� �;��<��=��O=��|=G|�=H�z=L�1= �<�KP����$��=�[�4�2���`����濚c�2�/�JiP�@�p�����jC��ڹ���I��_����[q��>Q�N�0����迍9�����w^7�>J�r�������	f���G;�>=�'h=�   �   V�j=�R=�$ =4��<0��;��Z��B�V*�.J�V�S�FUF��Z#�T�ۼx[*�`�<�\�<:�0=�+d=��|=&�n=�
+=HM <vzJ��D��&���}�1����^r��;�⿈���,���L��l��������t����'ǃ��wl�BOM�j�-�������+���f��3�3�@�����P(�8�_��'C;�=�&\=�   �   >�3=J%=t;�<�=̻ /����Y���񷽚�̽2ӽu�ʽ!3��������L�4~ؼ ��@�<"
=T"E=��H=γ=PV�;�1:��k�ˈ���پ��'���r�奿q*ؿp[��4$�l�A��^�n�w��D���@���,��2\w�ʴ^�j+B�<�$����ٿKJ���+u���)�_�ܾ)�������$N� a%;��=�=7=�   �   �<���:lμ�zh�5.��Co��� ���3�oB��%G��LA��|1�48�����%����qX�J��P3�;�:�<\S=�$�< ��;\	#�����f��Mľ���a^��k��;ǿ�����5���1���J��/`��n�L�s��5n���_��lJ���1�N�wc��_ȿm_����_�bb�mEǾ��k���@�4�@��:T��<�h�<�   �   �nf�^!:�j�����9�R�j�%P���~��_��.ાB���24��������f���5�.U�Փ��*��+(��b<0�e<�w�::�
�
�Ľ�sE����l����C�����r��߿&�����T53���D�aP��LT�0�O�p�C�p2�fe����C�޿����񙇿��D�ذ��W��y�I���̽���`�(��?*<���;�   �   ��{��Yὖ .�Bns��0�������T�1/��/��������ȅ��<&߾�E��춛�ŵn���)�Duٽ~�m��¼����ֻ�6ƞ�U$!�㌾r�߾.{%� �f�8n��us���@�^J�����#(�"T1�Z4���0�O'���p��4迉翿�H��h�f�_&�z2�ka���)$��ɤ�@ �����Y��Wݼ�   �   +���oG��������э���J�'y)��:���E��[I�D2E�_�9��(����ߏ�	M���_���C�o���n��|�8���ݼtv������^�A.���%�Y�<���{��
����¿r�㿀� ���TQ�6������A�]U���F�H���:����z���<��3�?���
�_��A���l~�������O���   �   r�N�y^��"׾^�{0�xUR��+p�w������4_�������􂿀Gn��[P�<�.����n�Ծ�����K�֯��9���@��L��*�;�F���<%�2���aϾ���zZG�֊��~��1۷���Ͽ/k�1�-��!`�!�YFο�a���E��x�}��0F�h:�\�ξ���L�%�����LE?��>���J����	���   �   �����Aܾ�~���B���p��\��y���{����߹�`༿[N��삯�\������n�
EA�3>���ھ����(�@�$�⽤�v��&����xx�Ɛ�TB�����%<ܾ{���B��p��Y��y���P���Zܹ�+ݼ�BK��	����Y�����n��AA��;���ھ�����@���:�v��'�t��R�x�ߘ� ZB��   �   �fϾ���V^G�{������9޷���Ͽ�n�� ��c��$�*IοHd���G����}��3F�m<�@�ξq����%�(���VE?�|6��.B�����(����N��Y��X׾�Z��v0��PR�S&p�������a\��������Bn��WP�֤.�����Ծ�|��p�K�֩��݊����t���;�L���A%�h5���   �   D(���<� �{�����¿���@� ���@S���d���C�EX��uI�f����;��]�z���<�5�8���r�_�>D���m~��
�W�� ���hG�㨏�Z������G��t)�l�:��E�WI��-E�"�9��(�/��C��H��k\����C�	���9i��n�l���<�ݼ|v�i���'^��1���   �   �}%���f�Mp���u���C��K�R��v%(�*V1�\4���0��P'�����6�(鿿AJ��T�f��&�O4ᾈb��+$� ʤ������6�\>ݼ��{�KN�k�-�oes�n+������6N�(��|���}�~� ��; ߾�@��������n��)�mٽ�{m���¼pd��@ֻd?�˞��'!��匾Z�߾�   �   �C�;���t��_߿���8��73���D�,cP��NT��O��C�tq2��f������޿��������´D�����X��Q�I���̽"��@(��Z*<�ֳ;h:f�z:��⯽��d�9�w�j�>K���y���Y���ڪ����M/��J�����f�|�5��O�������)��	(�8w<��e<�K�:�
���Ľ|wE�N��Z���   �   �^�Dm���<ǿ�����6���1�z�J��1`���n�2�s�v7n��_��mJ���1��N�d��"ȿ�_����_��b��EǾ�k�؇�V�4����:���<Pw�<(1�<@
�:8�ͼjhh�}#��c������3��gB�.G��EA��u1�"2�,x��A���JcX�p3�� v�;�E�<~V=$&�<Pw�;�#�]�轡�f�Pľo���   �   ��r�@楿�+ؿL\��5$���A�N�^��w��E��WA��e-��F]w���^� ,B���$��m�ٿ�J��/,u��)�\�ܾ���2���"N���%;΍=C7=��3=\-=\O�<��˻���|Y��疽�跽U�̽�ӽ��ʽ�*��������L�Thؼ``����<=z%E=$�H=P�=�A�; 7:��m�^���,پ�'��   �   ��Es��H��$�h�,�l�L��l��������t��_��cǃ��wl�jOM�x�-�����俧+���f����3���꾕���o'�&�_�@WC;�=V*\=N�j=�S= * =���<0Ǔ;��Z� 2�HM*�4�I���S��LF�S#���ۼPD*���< d�<�0=�-d=��|=�n=�	+=B <�~J��F�6(��L�M�1��   �   �2���a��C���c���/��iP���p�⌆�}C��ڹ���I��>���`[q�D>Q���0��~�^��9�������]7�Iﾇ���(���f��H;�@=�)h= }=�kk=�q?=�V=�q�< �����r��2ռ/� �������ǼpL���;��<z�=P�O=l�|=�{�=��z=�1=`�<\OP�����$��t�#�4��   �   ����r��Y�⿎���,�x�L��l�N���,��%t������ƃ��vl�lNM���-�������*���e����3�k�꾿���N&�(�_��vC;6=B+\=��j=(S=`* =h��<�ɓ;ȥZ��1�$M*��I�d�S��LF��R#�\�ۼ�C*��<xd�<2�0= .d=T�|=��n=�
+=�I <*|J�pE�d'��~�r1��   �   n�r��䥿*ؿ.[�j4$���A� �^�\�w�BD���?���+���Zw�^�^�0*B�4�$�����ٿI���)u�X�)��ܾr������N�@�%;`�=�D7=��3=R.=�P�<��˻����{Y�Q疽跽-�̽�ӽv�ʽ�*��`�����L��gؼ Z����<�=r&E=��H=��=�^�;�1:��k�Έ���پz�'��   �   � ^�Dk��\:ǿ�����4���1���J�R.`�4�n�b�s��3n���_��jJ�(�1��L�Ua���ȿ�]��q�_��`��BǾ��k�����4����:ԧ�<|�<�4�< 3�:L�ͼ�gh�#���b������3�vgB�G��EA��u1�2��w������bX�82�� }�;�H�<�X=�,�<���;#����T�f��Lľ+���   �   g�C�����q���߿H������33��D�4_P��JT��O�t�C�Dn2��c�N����޿z���H����D�خ��T���I���̽ر��(��k*<@�;�2f��:�,⯽ԓ�)�9�D�j�'K��}y���Y���ڪ�󧦾@/��<�����f�\�5��O�G�����)��(��<f< �:"�
���ĽWrE��������   �   �y%�9�f��l���q���>�$I����!(�<R1�X4���0�*M'��	�Ѓ�41�忿�F����f��&�h.�e^��n%$�h¤���P���$�(8ݼ`�{�xM��-�%es�J+��o���N��'��p���}��}���, ߾�@��w�����n��)�}lٽ.zm�$�¼�B����ջ�+Þ�j"!��ጾ��߾�   �   5$�F�<�%�{������¿���� �J��O�L����� @��Q���C�p����7��~�z�:�<��0�M���'�_��8��P^~�xj��嫼\ �������hG�����1���߆��
G��t)�^�:��E��VI��-E��9��(�&��1��jH��S\��h�C�(����g��2�\���Xyݼ�lv�0����^�,���   �   �^Ͼp���WG�^���|���ط���Ͽh����\�:�Cο�^���B��λ}� -F�I7���ξ���Ɓ%�[����6?��"���;����������N��Y��.׾sZ��v0��PR�B&p�������\\��ܕ����Bn��WP�Τ.����	�Ծe|���K�����و��Ξ�l��v{;�]A���9%��/���   �   ����G8ܾ�x�_�B�"�p��W��Б��a~��8ٹ��ټ�H���|���V�����@�n��=A�C8�a�ھω��*�@���
�v�j����rx����rSB�^����;ܾ	{���B��p��Y��q���I���Sܹ�%ݼ�>K������Y��}���n��AA��;�ǉھ㍖��@�:�⽎�v��@���ox�Ȋ�PB��   �   ��N��V���׾�W�ss0��LR��!p����\����Y�����B�=n�*SP���.�@��H�Ծ�w��:�K����� ���.�����F{;�bC���;%��1���aϾp��hZG�Ċ��~��*۷���Ͽ)k�-�)��`�!�VFο�a���E��s�}��0F�]:�;�ξJ����%������=?��'���9�]��������   �   ����bG�1�������<����C��p)��:���E�FRI��(E���9�b(�H��q��B���W��&�C�.����_��&�������rݼ|mv�m���=^�.���%�I�<���{��
����¿k��|� ���RQ�4������A�[U���F�G���:����z���<�}3����l�_��?���f~��q�|䫼������   �   �{�MEὖ�-�^s��&��0���H�D!����� z�Hz��w���߾�:��D���¥n�)�>aٽim��k¼����@�ջ '�Ğ�v#!��⌾D�߾{%��f�1n��os���@�ZJ�����#(� T1�Z4���0�O'���n��4迉翿�H��g�f�Y&�\2�1a��))$� Ǥ�h����(�*ݼ�   �   `f��:�گ������9���j��F���t��QT��@ժ�����*��_����f���5�TI�������)���'���<8 f< ��:*�
��Ľ"sE�\��\��{�C�����r��߿"�����P53���D�aP��LT�.�O�n�C�p2�fe����D�޿����񙇿��D�ϰ��W���I�ȯ̽����4(�0r*<P�;�   �   �?�<@:�:��ͼ,Yh�A��,X�����3�H`B��G�4>A��n1�Z+��k��jz���PX�(��`޶;�[�<�_=�6�< ��;#�l�转�f�bMľ���Z^��k��;ǿ�����5���1���J��/`��n�J�s��5n���_��lJ���1�N�yc��aȿm_����_�]b�TEǾF�k������4�@T�:���<���<�   �   �3=3=0^�<��˻�����nY��ߖ�?෽W�̽�ӽE�ʽ�!������8�L��Lؼ@��x�<�=�,E=��H=��=�w�;*/:�8k������پ��'���r�奿o*ؿp[��4$�j�A��^�j�w��D���@���,��2\w�ȴ^�j+B�<�$����ٿLJ���+u���)�R�ܾ���5��4"N� �%;��=�E7=�   �   � k=�S=- =���<@�;��Z�$＄E*���I���S��CF�J#�čۼ�$*���<�p�<��0=�2d=.�|=�n=�+=pU <yJ��D��&��~}�1����]r��:�⿈���,���L��l�����~���t����'ǃ��wl�BOM�l�-�������+���f��1�3�;�����(�ܿ_�`HC;�=�*\=�   �   ���=��=(Kc=��.=���<@�j<���: ���Hg_�H5y�x�I����� ��;H-�<�==J�H=N�=�ܓ=t�=e�=�e=�m�<��߼)ڽ�)c��ľt(���^��	��Cȿ���
��ʩ2�0GL��(b�"q�@nv��%q�>Xb���L��\3��������ɿ9К�' b�4����Ⱦ"�k�������u�<:�E=3u�=�   �   츄=Wt=��G=�=���< �E;@�/��B��X�伌���ټ8��;廠�;`��<��&=
�c=��=��=g��=�!_=���<��ռ�<Խ�^�����D��Z�Yt���Ŀ[����g���/���H���]�nEl�gq��Bl��]�L�H�40��/�����ƿ�����]���تľeAf�/�㽦.	��/�<l}@=�k|=�   �   * Y=̅2=d��<�@<�d?��w�@�K�KD��o蓽6������y�<�0�ݼ�[Ȼ��x<�=�O=�;v=�~y=�L=\�<<ݹ�7Bý�%O�񍴾����bO��뎿�M��e�4L���&��>�4�Q�Ԩ^��Ac��^�N`Q��>��.'�����[�Ӭ���E����Q�� �������V���ѽ\����<V�/=z$\=�   �   >=� �<P-�����T��N¾����D���6�����}�
��s�d���V�q��＀���J�<d] =^�>=6�+= �<x�������+<8�ܓ���� �J=�H���a����ؿ�>����<.�b>?�p�J�HkN�4AJ���>��-�xz�jW��mٿB6��z���@)?�O�������>��(��0gż�}<�=R�#=�   �   �%;��ϼ��x��Ͻ%y��=���c������������m2���5~��V_�4�8����ýԅ_��$����<Ȯ�<� �<Q�<@�R��V��D��j51ྏ/&�r�g��+���`���g꿊	���I)�¬2�2�5� I2���(��<�^��>��Y���w��Ѩh�D`'�f��|}��`� ��Δ�8{��8�L<"�<P�<�   �   �� �r_���(	�A�E�d��S,�����Ҿ�߾���[�޾�'о�����1���s~�Y'?�u�����v�
��d}�X�A<x�4<0]�`-S�|���3Xe�+���� ���D�	��Op��eʿk��\��B���R����n�����X���k�uɿ�𥿏���P$E�W��8��I�h�p � c���V���;���;����   �   �9����W�k�ߓ���T;V���������T(�ub+�a�'�����!��P����ɾz@��*�e���Z����,��F�  �5 
�������p�1�i��؎�t � �W��ۉ�������ſ�K߿qB�}���N����t����ݿ�:Ŀ�X��T��h�V�d ���=���Jn3�h,���� �p�)� �Z����l�=��   �   �&%���}�����0|�'��a3��}M�S�a�x�n���r�X�m�]`�u�K�sM1�}������ư��y�D5!����j=0�L&��@�8�Ƽ��~�* ���]�{��������)���Z�^����㞿����gĿ��ο��ѿοN<ÿ1����}��ُ��V%Y�jz(�0��0𫾂,]��� �L‽��мX�3�8O���:�%y���   �   ��x�C��JI����%��N�O�t�)@��h������J�����rs�����K-r�'�K��$��v��g���	v�x&������\�p+{�x"�rb������'���x����TC��(�%��N�t�t��=��6e��ԣ��?G��"���p�����C)r���K��$�ir��(��� v�i#�)����Y��.{�x5�~k������,��   �   �¬�i�����)���Z��Æ�k枿���kĿհο��ѿ�ο?ÿ����(�������W(Y��|(�������/]��� �2䀽�м��3�d@��:�:��p��� %���}�����v���\3�5yM�t�a�x�n���r���m��X`�k�K��I1�������"ð�y�N1!�p���v70��"�����Ƽ|�~�@� ���]��   �   E���v ���W�މ�1���v�ſ�N߿�E��������8��M��M�ݿ�<ĿwZ�������V�0 �w��󡔾`p3�w.��F� ���)��xZ�\���p�=��/��j�I�k�玠�O;����ԫ����P(�Y^+�h�'�C��m�K����ɾ�<�� ~e�R��מ����,� �F�  �5 !����Ĺ���1�����   �   ���D�� ��|r���gʿ:�������T�@����R�����n��vɿ򥿭����%E�����9��8�h�j �� c��V�P$�;P�;����� ��U���"	��zE��_��'��B����Ҿ�߾^��&�޾0"оe���:-��l~�,!?����֛��X�
���|���A<p�4< l�5S�Ԥ���\e������   �   �1&�Q�g�e-���b��j��	�����J)�j�2���5��J2�ت(��=�P�����;Z���x��5�h�?a'����?~��� �ϔ��w��P�L< .�<x0�<��;��ϼX�x��~Ͻqr�e�=�p�c�&�����&��-��J-~�O_���8�q���	ýxw_�h����<ȷ�<�<�N�<`�R��Z��~�������4��   �   L=�����c����ؿ�?�4���=.��??��J��lN��BJ� �>���-�:{�X�nٿ�6�������)?���������>�q(���cż��}<� =��#=�	=�<�����}�RK�����������D0�9	�<����
�i�+���ȭq�0�}���X�<nb =0�>=��+=T�<t�������<?8����&� ��   �   �dO��쎿�N����M���&��>�`�Q�
�^��Bc��^�&aQ��>�F/'����=\�$���0F����Q�!�����^�V��ѽ�򼸭�<�/=)\=�Y=��2=Л�<�i<�4?��i�p�K�i<��P���+���S��2�y��;���ݼPȻ�y<�=�"O=�>v=8�y=��L=���<湼�Eý�(O�援�����   �   \�Z�%u���Ŀj����h���/�@�H�J�]�$Fl��gq�rCl�b�]���H�$40��/����یƿ�����]�3��P�ľ�@f�����+	�L5�<L�@=�n|=���=D[t=h�G=��=(	�<@F;��/�83���������ټ�噼��p/�;���<�&=f�c=��=�=J��=� _=���<t�ռ�?Խ�^�3��F��   �   ��^�
���ȿ����R���2�tGL��(b�@q�@nv�t%q�
Xb�L�L��\3����U���?�ɿ�Ϛ�P�a����x�Ⱦ��k���Z���z�<Z�E=v�=u��=��=RLc=��.=���<��j<���:p��� f_�5y�H�I�P��� ��;�+�<�<=L�H=<�=5ܓ=��=��=� e=�h�<P�߼V+ڽK+c��ľ#)��   �   X�Z�~t��5�Ŀf����g�ء/�R�H�2�]��Dl�tfq�8Bl�D�]���H�Z30�/������ƿ�����]�n��<�ľ?f����>)	��8�<��@=�o|= ��=�[t=��G=��=�	�<�#F;��/��2��,�似��p�ټt噼�
廐0�;��<&�&=��c=��==�=���=�!_=��<��ռ�=Խ�^�&��EE��   �   �bO��뎿TM�����K�X�&��>�b�Q�ҧ^��@c�ւ^�_Q��>��-'����;Z쿃����D����Q���������V�1�ѽ��򼀴�<b�/=�*\=BY=�2=P��<�l< 2?��i���K�0<��"�������-���y���;���ݼ�Ȼ0y<��=�#O=�?v=��y=��L=0�<�ܹ�7Bý�%O�却�l���   �   iI=����Ja����ؿ2>�B���;.�8=?��J��iN��?J�\�>���-�>y�VV��kٿ�4��&���#'?������)�>�9#���Uż��}<�#=�#=V=��<0����|��J��?������҄�"0�	� ����
��h�����d�q�<���j���Z�<�c =�>=��+=$�<(�������v;8�T���,� ��   �   �.&��g��*���_��+f꿘	�����G)�:�2���5�vG2��(�;�������V��&v���h��]'����z���� ��Ȕ�g���L<�5�<6�<`�;��ϼ�x�*~Ͻ,r�+�=�<�c���������-��--~��N_�h�8�N���	ý�v_�h��س<L��<�<HY�<x�R��T������틾�/��   �   ���H�D�����n��ScʿJ����Ԡ�BQ�������B�����i뿇rɿx����I!E����o4����h�r �Jc�P�V�pV�;�?�;����� ��T��["	�BzE�]_���&��!����Ҿf�߾G���޾"оT���*-���k~�!?�t��L�����
� �|��B<��4<�H��'S�����Ue�x����   �   /��Cr ���W�aډ����l�ſSI߿�?�[���������9�񿴶ݿ�7ĿV��%����V�r �W��ɜ��i3�m$���{ ���)� Z�p灼^�=��.�����k������N;i���ë�����P(�L^+�^�'�;��d��J����ɾs<���}e���	����,�x�F�  �6���j������²1�����   �   ѻ��q���3�)���Z�����ឿ6��,eĿ��ο��ѿ� ο>9ÿK���O{��v���<!Y�w(�����뫾&]��� ��ڀ��mмȳ3�4�� �:�o��f %�P�}�|����u�k���\3�$yM�e�a�j�n���r���m��X`�c�K��I1�}�����ð��y��0!�B����30� ��`��@�Ƽ��~�g| �&�]��   �   ��x�4
���>��P�%�N�X�t�);���b�����bD��A��n���	��j$r�t�K�1$�dl��^�����u���B0K���z�`��\�����'�N�x�d��,C���%�|N�e�t�z=��/e��ͣ��9G�����p�����>)r���K��$�Yr������v��"�|����T�H{�@�4Z�X���$��   �   �%���}�ó��q�s��CY3�uM���a���n���r���m��S`�ԆK��E1�����������y��*!������'0���������Ƽ��~�R~ �e�]�E��������)���Z�S����㞿����gĿ��ο��ѿ�οK<ÿ/����}��֏��R%Y�dz(����,]�ʟ ����<zм��3��0��z�:�j���   �   �(��u��~k�ˊ���I;����h��>���L(�,Z+�@�'�?����8D����ɾ�7���ue����d�����,�(mF� �`7�����������1�-�����t ��W��ۉ�������ſ�K߿jB�w���L����p�񿿹ݿ�:Ŀ�X��Q��d�V�\ �Й�����m3��*��� �p�)��
Z�L߁�J�=��   �   ظ ��M���	� tE��[��j"��悼��Ҿ0�߾��㾪�޾�о���'���b~�e?�<��n�����
� $|�(B<(
5<P@�|(S�ٜ���We������ ���D���Hp��eʿb��Z��>���R����n�����V���k�uɿ�𥿎���N$E�O���7��ڿh�� �nc���V��Q�;U�;(���   �    q;��ϼ��x�uϽ�l�|�=���c�ʭ��]��^)��$~��F_�ę8����8�½,d_����<���<L�<(a�<�zR��T�����91ྃ/&�h�g��+���`���g꿆	���I)���2�0�5� I2�~�(��<�\��?�� Y���w��Шh�@`'�R��T}���� �͔�Tp��(�L<�8�<t>�<�   �   *='�<`l��^p�)C������|��~��)������H�
�8]�[�����q�l�� �p�<&l =��>=h�+=���<\~��S����;8������� �J=�C���a����ؿ�>�����<.�`>?�n�J�FkN�2AJ���>��-�xz�jW��mٿC6��z���>)?�J����R�>�`'��X_ż��}<$=��#=�   �   �	Y=$�2=��<x�<X?�4^� ~K�5��lؓ���+��J~y��;� �ݼ@�ǻh:y<D�=�*O=jEv=(�y=Z�L=��< ع�eAý�%O�ۍ��y���bO��뎿�M��b�2L���&��>�2�Q�Ҩ^��Ac��^�N`Q��>��.'�����[�Ӭ���E����Q�� �����b�V��ѽL�򼜯�<��/=�+\=�   �   G��=(]t=�G="�=��<�sF; �/��%����伌�� �ټ֙�0��g�;l��<��&=l�c=��=��=-��=z$_=L��<�ռl<Խ�^�����D��Z�Wt���ĿY����g��/���H���]�nEl�gq��Bl��]�L�H�40��/�����ƿ�����]�}��ѪľOAf����r-	��3�<�@=:o|=�   �   ῗ=FJ�=�4�=��V=ܡ&=D��<��<@�9<P��;@�;x�<�/}<D��<�=��M=�ց=��=��='��=�٪=y��=�m.=����|��<�*�1ɚ�܃��D�6���}�T��
uҿ����DD��U)���9��E�^�H�8E�|:��)�n��., ��Կ�¨�Lo�� �9�����)���5��N���G[�Y�< i=� �=�   �   ��=�3�=k=�:=�j= $�<p< ���(��0һ`}W��Pz;(�j<�<r+=6Yf=(��=4�=<��=��=(��=�-= Ku��)��&�&�:w��!��!e3��Gy�`V���Ͽ�������h{&��6�TzA�<GE�zA��6�R�&�4G����9�п�ڥ�%C|��96�������l�0��Ԟ���F�L��<��d=Y��=�   �   ��y=��X=�~#=���<���;�]$���ʼ֤���/�ޑ6�t_'�R7�W���I�L��<ȍ=�CR=��=S��=�E�=_̃=��*= ��:B v�^'�<֍�����)�ll��8��l%ſ���2��"I��Z-��O7�x�:�>77�VA-��L�<�Z��/ƿ�g����n�s,�!Q龱���P�#�F)��h���G�<l.W=\�|=�   �   ��2=|,�<�<o^�����3}�������ʽU߽��K2۽�½a�����^���@�q�Т�<>e&=Xaa=PR{=�kj=R0#= ��;�lK���}�P�ξ*_�T6X�=o��*���aܿ�� � ��1�^�'���*���'�����p�-� �͐ܿ
���*����Y��3��hҾ��BQ���n��p�X��<�p>=f�M=�   �   ��<0h����������ֽ���z:.�ӾF��V��Z�U�S�&�B�$R(��l���ŽH~u��3ϼ���;&�<Ƣ/=��==�{=(�<���U�޽��W��Ȳ�q���W>���}��l����Ŀu濺��4���@�,��J���=� r�^�7(ĿIm����~��G?�c�qy����]����B5����:���<T�=4c=�   �   t����3W���Ž|��\J��}�#���(���Ʋ�B��C���.Z������g;v���A����x����2��"����<<��<�v�<��O<�ü�U����-��{������ �YbX�Y���"���ƿWN࿱��� ����U �Hr�A߿�rſVb��	���K)X�H'!���� ��.�1��γ�Ԅ�0o�;��<�s�<p�<�   �   D�}���齝25�W�|��ڣ�44Ⱦ5�,� ���i��=��`��*�Lľ�����jt���,��]ڽlW`��j|���#<��<�^<N<���k���� mf��A��F8���0�$�c����������̿z�ֿ�3ڿ�"ֿ��ʿĿ���棿�!��.b��0�>��h5���jg������v�X}v�(�<�u<�a�;����   �   �.�=D��]��f�������L�`R(�"�9�pcD���G�O�C�T 8�q&�b1����k�������,�=�����h�$ǈ��'�;o=< ���Ԓ
��5��RI(�Z��{�Ⱦ�
�ʱ3��^��惿�������mӬ�ڧ��I��O���Ɣ�V���Hw\�N�1������ƾm
��t8'���\���,B�x�<`�@;���{��   �   L�?�ё�5�̾<����(�KI��Jf��|�Wi��p���B�*{��%d�4G�F�&�t�ŊɾdF����;�W�ٽJJ��F�0��;���;�p[�d�R�a�߽^�?��͑�2�̾+��R�(�-{I�^Ff�D�|��f��������	{��!d��0G�b�&���ɾ�C����;�"�ٽ&J���F����;0u�;p�[�\�R���߽�   �   �����Ⱦ�
�@�3�&�^��胿u������֬������K������Ȕ�2���kz\���1������ƾ���H;'�.�������-B���<@�@;�ݩ���{��$�7D��Y��;������OI�N(��9�1_D�m�G�=�C��8��m&�h.����`���Z���u�=�����h����� 5�;�h=< !��ƛ
��<��DN(��   �   DE���:���0���c�� ��I��T���̿F�ֿQ6ڿi%ֿf�ʿ�����裿_#��Łb��0�����7���mg����T�v��v� �<�!u<���; ���"�}�[���+5��|��գ��.Ⱦ�x��� �����e��:��Z��x$�=Gľ⧟�dt���,��UڽjL`��M|�H�#<D�<X�^<�e<���k�ʼ�irf��   �   ��ᾕ� �weX��Z��%��A�ƿ�P�l���S� �z��HW ��t�Z ߿Vtſ�c��C�2+X��(!����x����1��г�<��@|�;���<Ȁ�<ȥ< v��6#W��Ž�u�UJ�N�}�E������������<�����UU��<����3v�^�A�����p����2� ��	�<|��<lv�<�O<�*üJ[����-��~���   �   W��oZ>�� ~��n����Ŀ�����~��$B�z����� ?�s��_忇)ĿUn��/�~��H?�7��z����]��뽸5���:���<d�=rj=0��<�����������ֽh��T3.�(�F��V�(�Z���S� �B��K(�>g�#�Ž�nu�tϼ0Ϡ;�2�<��/=:�==�z=��<R��é޽��W��˲��   �   �`��8X��p�������bܿ�� ���82���'���*���'�����q��� �̑ܿ�
��L+����Y�:4��iҾ9Â��Q���n�@�o����<�t>=ЕM=*�2=�>�<0"<�8^����!}�w��L�ʽJ߽��佶'۽.�½n����^��� �p�ܳ�<�k&=�ea=�T{=$lj=�.#=���;XsK�����}��ξ�   �   c�)��ml�:���&ſ	 �����I��[-��P7�R�:�87��A-�`M������{/ƿ�g��L�n��,�CQ龮����#��(�����L�<�1W=L�|=��y=��X=0�#=���<��;x/$��vʼr��أ/�>�6�LR'�+��@�� �����<p�=IR=��=���=QF�=2̃=��*= b�:`&v��)��׍�Ȝ��   �   ?f3�NIy�-W���Ͽ����L���{&���6��zA��GE�tzA�V�6�~�&�LG����4�п�ڥ��B|�N96����3�����0�?Ӟ��F����<(�d=���=�=�5�=>k=>:=8p=0�<h�< ����򮻀�ѻ�W��z;x�j<�$�<+=\f=)�=��=���=x�=���=Л-=�'v�>,���&��x��߭��   �   ��6�q�}�����uҿ-���~D��U)���9��E�`�H�"E�V:��)�4���+ �Կ|¨��n��I�9�����(����5��L���;[��]�<�i=��=���=�J�=e5�=��V=΢&=���<D�<8�9<���; �;��<(.}<,��<f�=�M=qց=Z�=0�=���=�ت=���=�k.=����u����*�ʚ�����   �   be3�.Hy�wV��Ͽ�������<{&���6��yA��FE��yA�~�6�·&��F����Oп!ڥ��A|�j86�R��J���l�0��ў���F�4��<J�d=#��=b�=�5�=�k=�:=�p=�0�<��< ������ѻ W���z;0�j< %�<<+=@\f=I�=��=�=��=��=@�-= �u��*��̃&��w������   �   ��)��kl��8��%ſ������H�*Z-�O7���:�T67�l@-��K�n�����-ƿdf���n��,��N�򀒾��#�Z%��8���R�<�3W=�|=��y=��X=�#=D��<��; -$�tuʼ���b�/�փ6��Q'��*�H@�����@��<ڔ=�IR=�=���=�F�=̓=^�*= ��:, v�Z'�.֍�b���   �   �^��5X��n��k���`ܿ� �<��*0�T�'���*�x�'�����o�*� ���ܿ���X)����Y��1�$fҾ����;N���n� �o�l��<�w>="�M=��2=�A�<@'<@4^���� }��v����ʽ�I߽���x'۽��½=�����^�,�＠�p����<Vl&=�fa=^V{=�nj=�2#=P��;�jK�m��}���ξ�   �   ����V>�0�}��k��9�Ŀ��������?��������<��p��[�)&Ŀ}k����~�E?�n�zv��>�]�0����4�@��:d��<8�=@m=���<@���x��b����ֽ"��3.��F��V���Z���S�ߙB��K(�g��Ž$nu�$ϼ�֠;�5�<��/=P�==0=x�<����޽T�W��ǲ��   �   ��ᾥ� �o`X��W��e!��~ƿ9L�L}���� �����T ��o�߿pſ*`��&&X��$!��������1�ȳ�tn���;0�<��<(�<<q��P!W�8�Ž@u��TJ���}�"���у�������<������@U��*����3v�:�A����&p����2�� �<�<T��<���<��O<ü�R����-�Ez���   �   M?���6�x�0���c�����������j̿һֿ�0ڿ�ֿ6�ʿ)���e䣿���q{b��0�����1��eg������v�(Ov��<�9u<0Ņ;������}�\��r+5���|��գ�Z.Ⱦ�x辽� �����e��:��Z��f$�+Gľϧ���ct���,�XUڽ�J`��D|�8�#<��<��^<87<���k�����if��   �   ��h�Ⱦ�
�2�3��^��䃿��������Ь�.���VF���	��YĔ����5s\���1����7�ƾ����2'�V鲽����rA� �< BA;�թ���{��#�6D�ZY��
������9I�mN(��9�"_D�`�G�1�C�~8��m&�_.�t��M���D���8�=�=���h�T���P]�;�=<������
��0��F(��   �   �?��ʑ�n�̾���[�(��wI�ZBf�Ա|��d������t{�d�s,G���&���ɾ�?��j�;�W|ٽ��I��nF�P��;`Ѹ;�[[���R��߽ۖ?�_͑��̾��<�(�{I�LFf�3�|��f���������	{��!d��0G�\�&���ɾ�C��n�;�+�ٽ(	J��F�0��;�Ǹ;�S[��R�!�߽�   �   �2D�@V��������?F��J(�"�9�[D�&�G���C�b8��i&��*�U��"��������=�%����g�d���`��;�=<����8�
�4���H(�"��L�Ⱦ�
���3��^��惿�������gӬ�ԧ��I��K���Ɣ�T���Dw\�H�1������ƾL
��
8'�t�T����A��<`TA;�̩�@�{��   �   0|}����Z&5��|�tѣ�x)Ⱦ s辜� �5��b�7��S��"征Aľߢ���[t���,��Jڽn:`�|�x$<�(�<p�^<�7<���k�N���lf�_A��28�r�0��c�u���������̿t�ֿ�3ڿ�"ֿ��ʿ¿���棿�!��(b��0�7��N5���jg�r��p�v��hv��< :u<p߅;�과�   �   �`��xW�J�Ž p�RNJ�f�}�Þ���~��Z���;7������P��R����*v���A����e����2��� ��!�<���<@��<��O<�ü]T��/�-��{������ �JbX�Y���"���ƿON࿩��� ����U �Gr�>߿�rſTb�����F)X�B'!��������1��ͳ��|� ��;��<(��<��<�   �   x��<�������ĭ����ֽ����,.�ЯF��U��Z���S�>�B�qD(��`���Ž�Zu�4�μ =�;�I�<>�/=��==��=��< ��&�޽~�W��Ȳ�c���W>���}��l���Ŀm濸��0���@�,��H���=� r�^�8(ĿJm����~��G?�]�^y��]�]����$ 5��t�:���<6�=�p=�   �   � 3=�M�<�G<
^���2}��m���ʽF?߽��体۽f�½Y�����^�X����o��˦<�u&=0na=\{=�rj=�5#=p��;*jK�����}�6�ξ_�J6X�8o��&���	aܿ�� ����1�\�'���*���'�����p�-� �̐ܿ
���*����Y��3��hҾ���P���n�`�o�d��<�w>= �M=�   �   �y=f�X=��#=��<�M�;$��_ʼ؊�b�/�Rv6�dD'�~�L'������́<��=QR=8�=y��=�H�=�΃=�*= '�:�v�'�#֍�y���)�ll��8��g%ſ���2�� I��Z-��O7�x�:�>77�VA-��L�<�Z��/ƿ�g����n�q,�Q龡����#��(������N�<3W=��|=�   �   ��=x6�=�k=R:=�s=9�<X�< �}������ѻ��V� {; �j<�0�<�+=�`f=]�=��=D��=&
�=S��=��-=� u�E)���&�/w����e3��Gy�_V���Ͽ�������h{&��6�TzA�:GE�zA��6�R�&�4G����9�п�ڥ�%C|��96�������U�0�AԞ��F����< �d=쨋=�   �   �F�=�9�=�ŉ=�@r=��M=�+=n=��<`��<Dr�<�<�G=�6=��a=���=��=0��=/��=6��=�@�=YK�=�+y=�3�<fx���V&d��z��"��!5I����������ο�c�	�D��*7�~"!�(?����NR	�_(��ϿP���V��EL�V����þXqq����G��X�;T '=f9~=��=�   �   ��=Z�=�R�=��Z=42=l�
=|��<�P�<ͅ<Lׅ<�<���<(=T�@= t=(��=D�=w��=b��=@�=h��=^Dx=���<l1���5߽z�^�撹�$�a�E�z���d@���˿x��<_����lb�0���n�����zx̿�^���5H����Yv��:�k�����t�=��=�;��'=8B{=�͑=�   �   A��=^q=��F=T=P��< �<�X���� �p�m�H�v�`�8�@�Y�(4<0�<=�[=猋=�5�=�n�=�f�=�ʡ=$u=���<�L̼Kq˽3dO�;���4���:���y���������㿸^ ��0����\|� ��#��e ��b�lT¿�ϟ�N�{��/=�|���v��([�~��"��F <8)=
�q=ǋ�=�   �   �#T=x.$=�%�<K�;X�c�B@�B�G���z����s����:����a���"��F�� ��9�0�<Ԡ,=�Cr=�Ƒ=Fr�=2
�=J�m=$��<����Y쬽\7�0����� g*���d����G��>0ѿ���F�$��[
����� �9쿥ѿps���f��m�e�=�+�4J�/ɠ��7A���ý�;�m<�t)=>�_=��j=�   �   PU=�I<��E���!��d���ý�.��ξ�yt�.�� ������㽻9��~�`���ɼ���;�
�<�4G=�Qx=롁=:�_=�2=�Eۻ`ۆ���h��1о�?���I�A��i��XF����ҿ�	��F�)[������o�x,ҿʹ��+��fG��K	J�� �ˀҾ/��2� ��U���:��L(�<�J%=*C=~34=�   �   @�y;d�Ҽ�|�B�ϽrO��V;��_���{��̆��^��Zd���hv�ʇW�� 1�)������yB���8���<Z =~�L=�_H=�U= �t;l�9�n���Y�b�������~�*�TH\�룇�$	��4w��e/ƿ?�п:ԿFRп�rſg���&C�����M�[��n*�����)���.o]�2~��ЕT��T���i�<\0=L�=�C�<�   �   ��o8���3��;�R0w�yƘ����@�ƾ�Ӿ1�׾�RҾ�@ľHˮ�����+<l��8/���ց�l����9<n�=��$=:(=��Z<�D̼�7��� &��҇�<�ȾX^
��4�7_�J���y����������/y������ۣ�5���;V���]���2�Q�	�a�Ǿȕ����&�Zǭ���꼀�<��<Z�=0z�< ��9�   �   eϟ�h��UST����,B��-j����d���L�����������޾�M���ˌ�	RJ���^��`	���<���<��=ԧ�<P�ƻ\�N��?�<�H�y�����վ�����/���Q���o�Pd��S���y��L��������m�f�O���-�Z��Ӿ�p���E��R佤L� �q�< c�<�ù<��3;����   �   S
��9Y��B��zѾ{����� 6�t�H��%T�g�W��^S��G��/4��c������̾fS���;R�2�ك�\��� ]I<��<�<�<�m$<X*��d������3Y��>���Ѿ�������6���H��!T�`�W��ZS�G��,4��`�L���̾lP��7R���ԃ�����eI<0��<X6�<8U$<�=��Z����   �   ��H������վ���8�/�{�Q�Ӆo�}f���������;N������1�m�z�O�q�-�q
��
Ӿ�r��4�E�2W�\L� !Ỹp�<�g�<�͹<@d4;4���dǟ����LT��ۑ�6=��zd�ф�}�kI�<������B����޾vI���Ȍ��LJ�����������(
<���<b�=П�<0�ƻz�N��G��   �   �Շ�+�Ⱦ�`
� "4��:_�L���{��˦������z{���!���ݣ�����W����]���2���	���Ǿ����,�&�Pʭ����8�<L�<T�=P��< a�9���/��.��:�U(w�����������ƾ:�Ӿ��׾�MҾ�;ľ�Ʈ��򓾄5l�B3/� 꽼ρ�y��H�9<��=��$=N&=ȯZ<U̼�=��%&��   �   ����Ȟ���*�hK\�����#��[y���1ƿ��п�<ԿhTп�tſ%����D�����S�[�op*���̩��`q]������T�`Z��4l�<v3=x�=�R�< 2z;��Ҽ�|�ڴϽFI�zO;�*�_�N�{��Ȇ�,Z��"`���`v���W���0��#� ���XlB��8� '�<�^ =��L=�_H=\S=`dt;  :��t�r�Y��   �   Eо�A��I��B���j��7H���ҿ��I�>]�����q�.ҿd˹�
-��FH���
J��!�%�Ҿ�/��B� ��V��p;��<*�<M%=*C=V94=.]=p=I<p�E���!�i[��n�ý#�����n��|��{�F���㽃0����`���ɼ�܆;�<�9G=Ux=���=|�_=�/=�qۻ�߆�������   �   ڝ��h*��d�Q���~H���1ѿ���.���\
����~� �J:쿯ѿEt��cg��b�e���+�K�ɠ�)8A�1�ýx;��m<�v)=Z�_=�j=z)T=�5$=\8�< ��;��c��1��G�l�z��v������;2����a�4�"��,�� 1:�B�<�,=>Ir=yȑ=Ks�=g
�=�m=��<X�����_7�M����   �   6��:�s�y����������h_ ��1�r��}�����#��e �Zc��T¿П���{�%0=�����v��([�1��ƙ"��L <�9)=��q=b��=J�=&cq=��F=�=0��< �<@��g �H�m�X�v��8��[Y��X< (�<�=��[=��=�7�=�o�=�f�=�ʡ=~�t=l��<tV̼ u˽�fO��<���   �   %���E�$���#A���˿�x����_����b�x��4o���￉x̿�^���5H�����u��~�k�����V�=��M�;z�'=@D{=�Α=��=��=jT�=��Z=�2=^�
=�	�<�[�<T؅<@�<h��<,��<D,=��@=#t=R��=��=���=���=,�=���=�Bx=��<�9��9߽��^�P����   �   ����5I� ��@��?�οd�@	�b��87�~"!�?����&R	�(�W�Ͽ�O��XV��� L����Øþ�oq����xG��m�;V'=;~=��=TG�=H:�=7Ɖ=�Ar=l�M=�+==��<���<hr�<��<\G=��6= �a=a��=1�=¥�=���=���=8@�=�J�=�)y=�.�<�{� ��'d��{���   �   R$���E�����j@���˿�w�r��_�l��b�ȋ��n�^�￧w̿�]��o턿�4H�
���t����k�����b�=�p^�;�'=hE{=jϑ=Q�='��=�T�=D�Z=62=��
=�
�<`\�<�؅<��<؉�<���<z,=�@=>#t=o��=9��= ��=���=v�=X��=�Cx=���<|4��7߽&�^�J����   �   �4�K�:�.�y�b���p����T^ �R0�,���{�l��L"��d �ia�7S¿�Ο�n�{�O.=�=���t��L[�*���"��\ <�<)=��q=A��=��=ddq=
�F=�=��<H�<�����d � �m���v�p�8��UY� Z<�(�<6�=�[=I��=�7�=�o�=}g�=Pˡ=�u=h��<L̼6q˽dO��:���   �   ��Tf*���d�a���3F��;/ѿ쿌�R��Z
�0���� �C7��ѿ�q��ie��&�e�_�+�AG��Ơ�34A���ý�+�03m<{)=r�_=r�j=�+T=�7$=p;�<P��;`c�j0��G���z�6v��0����1���a�ȵ"��+�� M:�C�<��,=Jr= ɑ=t�=��=R�m=���<����B묽B[7������   �   �о�>�S�I�>@��h��E��p�ҿ��E�Y�����m�m*ҿ+ȹ�9*���E���J����}Ҿ�,���� ��O���(���7�<R%=�C=H<4=�_=�EI<P�E�L�!��Z��ßý~"��T���m��|��{������D0��L�`�ȡɼ�;��<8;G=�Vx=壁=|�_=�5=�+ۻoن�L�q���   �   ����V����*�IF\��������ru��j-ƿ�п<8Կ�Oп�pſ9���"A�����(�[�@l*�����椭�5j]��v���T����{�<�8=��=lY�<�\z; �Ҽ�|��Ͻ�H�O;�֜_��{�qȆ�Z��	`���`v���W�`�0��#�Ǯ���kB� �8� *�<�` =��L=�cH=�Y=@�t;<�9��j�m�Y��   �   ч���Ⱦ�\
��4�V4_��H���w��w���x����v��]���٣�	���9T����]���2�Ń	�I�Ǿ������&�迭�L�꼈<|"�<��=؏�< �9���.���-���:��'w�����Ψ����ƾ�Ӿq�׾mMҾ�;ľ�Ʈ���Z5l�3/����9ρ�0v����9<Ȉ="�$=�,=�Z<�8̼�3���%��   �   |�H�𥘾��վ���D�/���Q�~o�Rb��.���@���I��p�����m���O���-�}�Ӿ�l���yE�tI�tL� ��@��<�v�<�ع<`�4;����Ɵ����LT��ۑ��<��Jd㾻���|�[I�.����}�8����޾bI���Ȍ��LJ���(��������<@�<Թ=̲�< Sƻ"�N�:��   �   ���.Y��;���Ѿ����6�ڃH��T�Q�W��VS�G��(4��]�P��ٷ̾CL��h0R�����̃��s��ȑI<��<lJ�<�$<�"������3Y��>��MѾp������6�s�H��!T�T�W��ZS�G��,4��`�D��ڼ̾ZP���6R����Ӄ������uI<��<�G�<x�$<8������   �   ������GT�gؑ��8��x_����y�F���3������޾hD��PČ��EJ�P����ݽ�H9<��<��= ��<�bƻ�N�J>轺�H�A�����վ�����/���Q���o�Hd��K���t��L��������m�a�O���-�U��Ӿ|p���E��Q�HL�p�ໄ{�<�r�<�ٹ<@�4;�����   �   ���(���)�_�:�X!w�ý��D�����ƾ��Ӿ͘׾�GҾ6ľ����KR-l�N,/����\Ɓ��Z����9<�=��$=j/=��Z<D=̼16��< &��҇��ȾC^
��4��6_�J���y��}�������)y������ۣ�2���9V���]���2�K�	�M�Ǿ������&�iƭ����8<�<��=���<�O :�   �   ��z;8�Ҽ��{���Ͻ�C��H;�ȕ_�,�{�>Ć��U���[��Xv��xW�B�0�m�9���ZB��e8��?�<�h =��L=�gH=�[=��t;b�9��l�n�Y�8�������m�*�BH\�㣇�	��,w��^/ƿ9�п{:ԿCRп�rſe���#C�����H�[��n*���������n]�q}��t�T�`8���t�<8=��= a�<�   �   :d=paI<PcE��!�S����ý������g�$v�/u�����㽪%����`��ɼpL�;X1�<�CG=^]x=:��=��_=J7=0+ۻ6چ�6�>��о�?���I�A��i��RF����ҿ�	��F�&[������o�v,ҿʹ��+��fG��I	J�� ���Ҿ /��� ��T��5���0�<�P%=~C=�>4=�   �   �.T=V<$=|H�<0�;hUc��#���G���z��m��V���)����a���"�,����:�Z�<(�,=�Qr=&̑=~v�=W�=�m=��<����~묽�[7�������f*���d������F��90ѿ���C�"��[
����� �	9쿥ѿqs���f��l�e�;�+�*J�!ɠ�^7A��ý�7�X$m<2y)=F�_=��j=�   �   ��=gq=��F=�=Ш�<�<�ڻ� = ���m� �v��`8���X�x�<�;�<ʎ=v \=u��=�:�=r�=@i�=�̡=u=��<pI̼�p˽ dO��:���4���:���y���������㿷^ ��0����\|��� #��e ��b�lT¿�ϟ�M�{��/=�z���v��[��彊�"�xN <�:)=��q=s��=�   �   h�=���=fU�=T�Z=�2=,�
=��<te�<��<L�<���<`��<�1=��@=�'t=l��=���=���="��=��=f��=�Ex=���<�/���5߽`�^�ܒ��$�\�E�y���b@���˿x��<_����nb�0���n�����{x̿�^���5H����Vv��,�k������=�PE�;��'=2D{=-ϑ=�   �   <}�=M�=���=��u=�a_=R�J=ܲ:=v�0=�F/=��6=PG=��`=ɀ=�=v��=ü=~g�=�.�=X�=���=��=�P�=:�C=`�&;�{�	��ܱ���tӾ����,M������a���콿�6׿e7�M��8���?'���_��׿oz��'%��쓄�>rO������پ{I��W�*�����e����<p�8=
�y=��=�   �   hэ=f��=(}=�c=$�I=.�1=T>=��=��=�)=�&=��@=:�c=���=7՜=Ψ�=�= �=tF�=$>�=l��=�˟=�F=��;�lq�.��«��y0Ͼ� ��xI�V�������ź���ӿV�s��o\��s���o翟�ӿ>���U��
6��~�K�����?վ� ��R]&�ǣ��۫��!�<L:=��x=��=�   �   �x�=��p=|cQ=��,=8=���< <NK<@�(<�|:<��<@��<
6	=z>;=�q=�=O��=&-�=8��=4w�=N��=/ �=*L=��<�6S�e����w��¾���s�>��Vu���������Yɿ/ܿ���,�远ܿUiɿcֱ�-*���v�`i@�4��uȾ�{�� ��&z����x����<�r>=�t=�F�=�   �   ,�\=,G7=4n=D#�<���;�K�����dO�����0�\��|2��pB�� w5<��<�>=���=�o�=&x�=��=Fg�=�8�=��S=�Rj<J�$��Q��e\�'x���.��d�-��f`��4��S&��<(���oʿ$uտ�0ٿlLտ�3ʿ�������r\�� a��.�*�"���fNg�X��1j�`�л��<<-C=L�j=�hp=�   �   �� =�B�<pӦ;����r��r�k��%���q���*Ž��ǽ�뻽V����N}��#� ��H�<0=VV=i.�=��=���=�m�=�[=���<@�Լ������9�����޾L�W�E�`t����l��	볿�½������������� ���M���
t�ۯE����"�߾�ę�n�A��kӽ2�"�P��;z�=,�E=$rY=z�J=�   �   �ř<p晻���w݁�o�½|g �"��0�0��P=�NV@�X99�$y(�����M�s���BD-� �����<`�/=8�s=��=Հ�=^�^=���<��+��Ӊ�(� w�ٯ��2����>'���O���v�ż���;��?Ȣ�����B|��ϸ��s!���u���N���&�4l��︾iTy�����1�������L�<�=�GB=ܒ==m=�   �   �u	��E-������ ��)/���[�h�����P����N��LИ�������x��UN���R�ݽ���������y1<�3=�X=��p= �[=��= %�;�*�(cֽ}`>�#��{�;���ѣ)��J�f�g��`~��c��S������T2}��f�0�H�R(�3C��r˾�����=���׽.6� 	P���<�K,= W6=R =xǔ<�   �   �A/�Ô��P���lQ�y���P§�`Kþ��ؾ�b�t�꾍�來�վD���c�������B�(��������<��	=��D=:�O=�(=�˙<Ȑ��+��$����Y�/̜�q�ѾnT�$��
�6��I���T�_�X�T��G��4�[���;���;� ��HHS�\��}΂��=��t�<2]=�5=�W=�3�<�Q���   �   ���BV���`�`q���1ľ
��n>	�W���� �
�#�' ��C�U?�m���Ѿ��ғ�|U�F��D�� PҼp]/<�|=D�9=��3=`3�<0Q�;��
�>���eQ�D�`��m��c-ľä�;	�9���� �٪#� ��@��<����Hξ��ϓ�UwU����f?��BҼ�n/<�~=&�9=v�3= *�<��;��
��   �   \��z�Y��Ϝ�ԭѾW���O�6�I�$�T��X�uT�5�G���4����>��;|��LS���C҂��F���ܑ<�\=T5=�[=�?�<�	��85/�������xfQ�����⽧�tFþG�ؾx]�~�N�侣�վൾ��������\�B������ ��@�<p�	=�D=��O=��(=l��<𡌼11���   �    e>� &��_�;[����)��J��g��d~�ce��,���]���5}��f���H�k(��D�>u˾뱐��=�\�׽�26���P��<�L,=�Y6=.%=�Ք<hM	��8-������ �l#/���[�q������昚�J��̘��|��j�x�SON�����ݽ�{���q��`�1<�8=�X=��p=��[=�=��;Z*��iֽ�   �   �w����8���OA'���O�%�v������=��ʢ�u����}��g����"��|�u���N���&��n�����Vy�����3������8K�<��=�IB=��==�r=Tՙ<Г��̶�lՁ�ܢ½�a �����0��I=�wO@��29��r(���D�%����6-���D�<F�/=�s=��=���=v�^=���<�,��؉����   �   D���<޾N���E��bt������m���쳿HĽ�c��7���b�������N��it�B�E������߾�ř���A��mӽ$�"�@��;��=ċE=uY=��J=v� =TR�< #�;�s��*}��k����!h��� Žjǽ�ỽ#�=}�\�#������<h=�$V=�0�=q��=4��=Fm�=D[=̷�< �Լκ��&�9��   �   \z���1��(�-��h`�6���'���)��qʿ�vտ2ٿ�Mտ5ʿ�������]�� a���.��*�ը��HOg����2j�@�лT��<�.C=��j=�kp=��\=�L7=Vu=�4�< ؚ;(�����4漴���"���༸���䠻H�5<���<>=f�=�q�=�y�=��=wg�=!8�=@�S=�Aj<ڐ$�pV�i\��   �   ��¾ا��>��Xu���������)ZɿIܿ���-���fܿ�iɿ�ֱ��*����v��i@�k���Ⱦ�{�����y��@�x����<t>=rt=�G�=z�=��p=>hQ=R�,=�=��<�ҍ<qK<P)<��:<��<p��<l=	=�D;=��q=N�=��=p.�=��=�w�=3��=���=�L=��<�<S�y��v�w��   �   �1Ͼ��zI��V��H���dƺ�W�ӿ�V����\�����p���ӿ5>��V��6��c�K����N?վ� ���\&�#ƣ�`ث��$�<|M:=�x=��=bҍ=���=�}=4�c=��I=�1=�B==�=.=&&=V�@=��c=��=m֜=©�=��=t�=�F�=>�=��=�ʟ=<F=p΂;rqq�ڊ�ܬ���   �   ~uӾ��u-M�I���Bb��	��6׿�7�e��=���)'���_�Ҍ׿'z���$�������qO�%����پ�H��-�*�����`��T��<�8=\�y={�=�}�=��=(��=X�u=�b_=��J=`�:=��0=2G/=��6=@G=n�`=�Ȁ=��=&��=�¼=$g�=\.�=�W�=6��=q��=�O�=.�C=`�&;��{�4�������   �   �0Ͼ�yI�V�������ź�q�ӿ�U����[�����o���ӿb=��PU��l5��i�K�Շ�&>վ�����[&�cģ�(ӫ��(�<�N:=X�x=�=�ҍ=�=�}=��c=R�I=��1=C=�=`�=f.=j&=��@=��c=2��=�֜=ݩ�=��=��=�F�=L>�=f��=p˟=�F=�߂;8nq��������   �   ��¾l���>�OVu�K������pXɿiܿ���+���翁ܿ<hɿVձ�3)��Y�v��g@����|Ⱦ;z������v����x�軹<�v>=�
t=�H�=�z�=&�p=�iQ=��,== 
�<tԍ<tK<0)< �:<��<P��<�=	=>E;=�q=��=E��=�.�=f��=x�=䆾=� �=�L=��<�6S�F��^�w��   �   gw���-����-��e`�54���%��A'��znʿ�sտO/ٿ�Jտo2ʿ���y��9[���a�=�.��(�˥���Jg����)j��Sл���<�2C=ؕj=�np=]=O7=Vw=T8�<p�;8�P����1漾��"����|���࠻X�5<|��<�>=��=9r�="z�=|�=th�=�9�=D�S=�Yj<T�$�RP��d\��   �   �����޾K��E�V^t�����j���鳿 ������?������
L���t�t�E�߾���߾`���A��eӽ��"�p��;>�=��E=yY=4�J=p� =�W�<�5�;8o��{�D�k����tg�� Ž�~ǽgỽ�2=}���#�����<=n%V=/1�=B��=Z��=�n�=6[=$Ʊ<p�Լy����9��   �   ;�v�򭸾����;='���O���v�Y���7:���Ƣ�Ϛ��dz�����������u���N�{�&�h���븾2Oy�����+�� ���t]�<��=<OB=�==rv=�ۙ<�|��$��3ԁ���½za ����A�0��I=�2O@�~29��r(�����C�ѭ���5-���4�<��/=��s=�=���=�^=|��<��+��Љ�)���   �   t]>�!��Ɗ;?����)�S�J�q�g��]~��a��v�������.}�\f���H�s(��@��n˾�����=���׽�!6� �M��(�<T,=\_6=�)=tݔ<H@	��5-�>��� ��"/�V�[�:�����������I���˘�~|��8�x�(ON�R�a�ݽm{���o����1<�:=bX=|�p=2�[=4�=@O�;	*��^ֽ�   �   ����Y��ɜ��ѾTR����)�6�kI�$�T�̌X�wT���G���4�T��L9�3�;0���HBS����ǂ��%�� ��<�e=J5=�`=|H�<�쩻2/�1���r���eQ�Z�������>Fþ�ؾP]��}�1�侊�վɵ������q��0�B���i�����H�<�	=��D=�O=Ή(=�֙<����j&���   �   W����M�H�`�^j���)ľ0���8	�O��z� ���#�� ��=��9���辎ɾ��˓��pU�j���6��'Ҽ��/<�=Ĝ9=*�3=T=�<�q�;z�
������P���`�Am��#-ľ���j;	�$���� �ʪ#� ��@��<����6ξ��ϓ�(wU�����>���>Ҽx/<�=(�9=��3=�>�<P��;��
��   �   p*/���������`Q�@���鹧��Aþ@�ؾX�sx꾼��A�վְ����������B�v��������8<f�	=��D=̮O=��(=`ԙ<�����)�����X�Y��˜�4�ѾRT�����6��I���T�T�X�T��G���4�T���;���;� ��HS����͂�X9����<�a=:5=�`=�L�< ǩ��   �   �'	��,-���� ��/�F�[�������������E���ǘ�6x��>�x��GN�����ݽ�r��HS��X�1<,C=|X=��p=��[=��=pC�;�*��aֽ�_>��"��F�;����)�χJ�U�g��`~�~c��O������M2}��f�+�H�K(�,C��r˾毐��=���׽J,6��dO��<tQ,=�^6="+=��<�   �   �< E������́��½�\ �#��)�0��B=�eH@��+9�$l(����p8���%-��}� �<��/=��s=��=j��=��^=���<��+�d҉�� ���v���������>'���O���v������;��<Ȣ�����?|��θ��q!���u���N���&�(l��︾?Ty����1�������R�<��=NB=��==�x=�   �   �� =�a�<�n�;�\��|o�L�k����r^��nŽ�tǽN׻��䢽�*}���#�聼8<�=D.V=�4�=���=Z��=Yp�=�[=�Ʊ<d�Լʹ��7�9������޾L�H�E�`t����l��볿�½��������􅳿� ���M���
t�دE�����߾�ę�F�A�Zkӽ��"��˒;�=�E=�xY=��J=�   �   �]=dR7=|=E�<`%�;��� �����T���Ll�����px���5<���<�$>=���=yu�=�|�=��=j�=�:�=��S=(\j<��$��P콀e\�x���.��Y�-��f`��4��O&��9(���oʿ!uտ�0ٿkLտ�3ʿ�������q\���a��.�*����HNg�*��0j��|л ��<�0C=@�j=dop=�   �   l{�=��p=�lQ=��,=�"=��<P�<@�K<�8)<(�:<�%�<�¾<F	=M;=�q=��=쓬=�0�=:��=�y�=��=��=&L=��<�5S�*��m�w� �¾���l�>��Vu���������Yɿ,ܿ���,�违ܿUiɿcֱ�,*���v�^i@�3��oȾ�{������y����x����<u>=�	t=�H�=�   �   �ҍ=)��=�}=^�c=T�I=<�1="F==N�=�2=�&=��@=�c=.��=Y؜=���=I	�=���=�G�=P?�=L��=W̟=�F=��;lq�������q0Ͼ� ��xI�
V�������ź���ӿV�s��o\��r���o翟�ӿ>���U��	6��}�K�����?վ� ��D]&��ƣ��ګ�D#�<.M:=*�x=��=�   �   �Pf=
�b=�[=��S=4�M=��J=��K=�Q=x�\= �m=h>�=j�=��=ܲ=�<�=ڮ�=l��=�]�=���=�	�=���=���=��=V0
=�i���O���1��.���rؾ����A��0p�yk���3��(ʱ��ǻ��:���ѻ��豿�s��֎�{gq�B�C��I�=�޾�M���qF��_㽰M���滼ɲ<ƪ#=��M=�Qa=�   �   �vb=�^\=@R=��G=�c>= T8=̓6=�(:=��C=^T=<�j=�	�=JF�=�C�=zػ=(��=���=v��=�s�=n�=$��=<�=�/�=@=�n�SP����,�����fԾ�2��S>�~�k���m��:Į�j���U���ќ��ٮ�����`N���m���?�fS�r�پ�і��OA���۽~MB��ɩ��$�<��&=f�N=��_=�   �   P8V=�H=�05=@*!=x�=���<<��<���<��<Q=�q=�U<=�c= ��=C�=��=�d�=�b�=��=���=Y�= ս=�ɐ=p�=h2�[�������Q�Ǿ��	��4���_������W��|����R������GJ���Qg����uJ`�D85�����̾����k2��Mƽ80#� tH9�<b�.=FP=��Z=�   �   ��?=��#=��=h߻<0�k<���; �v:��+�`,Z� [��-�;��d<��<�� =,p\=���=�g�=]9�=��=U�=��=���=��=b�*=@옺��s�Jo���n�"鳾~L����#�4L���r�󨊿�-���̠�3����������������r��aL���$�D�������|�y��-�f����a�؉
<|'=b
:=
Q=��P=�   �   Z�=���<@�R<�OպK��H��$%�"�D��TS�:dN�f5��s�ĸ�����$��<p�=N�i=��=��=���=���=~��=���=��>=�f<�0�M0作�J��)����پ�~�Ye3�&V�j�t������A��ؐ�c��NE��
Gt�$�U�3��y�׭ھ :���Q�:Y��27s� �U�,D�<H%=R�E=�N=�>=�   �   ܂�< ��;�L]��D��n�|A��dWǽ�⽗"��%���ȽDˠ���_�4L缀ڹ��	�<t�>=u؄=u؞=~8�=�է=递=X�Q=P��<`�̼�۫��?"��~��k�����nt�Sv5��P��	e�Xr��v���q��8d��O�f]4��m�P�lj���~���$�����NR���q;4��<\�7=F�M=�D=��=�   �   ��;�꙼��F��v����轋��|�0��+F�V�R���U�p�M��Z;�I� �,J��)N����W��9��huV<d�=~bo=p�=Vu�=H�=N�`=<a�<`8⻲3e����KF������z����� |���)��';�O:F��I�|�E�}:�:(���`V�佾g����?A��m�4�f�`�6��ת<��'=z�N=x$P=�0=�H�<�   �   �����~U����HU���<�j�Z��㶘��Q��椾X���P��4���$BY��|(��d��V��4�㼀��;�=h#^=��=��=�%i=��=�� <�>�Q~����+X��Ó�U���徵S��N�,#����8l���Z[��1�׃��덾wL��'������u��0%Q<�=��P=l8`=�I=��=8�U<�   �   �::�ao��H@�ĨT��%������Kľ��پ��j%��T��1־+-���o�����b�C����3���g��7�;�=��T=��r=.6i=D�8=���<P]ͻ�/:�Ch���;��T��"��񨾄GľA�پ�美 �KP徐-־F)��Tl��B~����C�I���.���W�Pe�;��=��T=L�r=�4i=J�8=\��<@�ͻ�   �   �����P0X�4Ǔ�<
��M�2V�)Q��%�_���n�����]�i5������퍾�zL��*�#�������Q<��=��P=9`=F�I=��=V<u���rU�o��P��<�tj����𲘾qM���᤾`��M��ޚ��W<Y��w(��\�P���q㼀��;��=�&^=Z�=��=�#i=��=�� <�P��   �   ��FPF�}���~��J��n~�f�)�^*;�4=F���I�:�E�:�F<(�	���Y�潾gÌ��BA��q�^�f���6� Ӫ<`�'=��N=�%P=�0=pR�<�;�;�י���F�;o��o��@����0�l%F���R��U��~M��T;�֙ ��@��F��p�W��$����V<Z�=�fo=Dq�=�u�=�G�=�`=TX�< p⻮=e��   �   qC"����n��5��v��x5�TP�ze��Zr���v�A�q�J;d��O�H_4�]o��R�Ql����~�� %�����V���q;���<B�7=8�M=�D=n�=���<�*�;8']�9��n�J9��CNǽ?��R�;�	�w�Ƚ� �Ԇ_��2�������<��>=�ڄ=ڞ=`9�=�է=Q��=��Q=t��<@ͼ�૽�   �   1�J��+����پS��qg3�!V���t�O����B��eِ����mF��It�ΔU�m3��z�u�ھQ;����Q��[��<:s���U�0B�<"%=�E=�N=d>=P�=x��<��R<�6Ժ�5�����t%�t�D�XES��TN�h5��e���������<�=ȱi=���=ϰ�=銽=���=`��==��>=�R<f�0��5��   �   �n�J볾.O��;�#�!L���r�����.���͠�I�������v��d�����r��bL���$�o���������y�c.�J���d�Ї
<�'=�
:=BQ=��P=��?=��#=��=��<l<�8�; By:@X+��Y���X�P��;xe<��<�� =
w\=���=,j�=;�=	�=�U�=,��=l��=���=0�*=�����t��q��   �   Å�%�Ǿ�	��4�-�_������X��X���`S��k����J������g��'�K`��85�@��u�̾����Ik2��Mƽ0#� �H9��<�.=&GP=��Z=B:V=RH=�35=d.!=j�=̾�<���<԰�<���<�W=�x=,\<=ޗc=���=3E�=m�=�e�=�c�=���=D��=�X�=�Խ=�Ȑ=d�=hD���՚��   �   �����Ծ�3��T>���k�Y󋿚m���Į�㗸�����&���Fٮ�͟��xN���m��?�RS�9�پ�і�JOA���۽LB� ����&�<��&=l�N=��_=�wb=�`\=BR=\�G=Vf>=W8=�6=.,:=<�C=�T=��j=Q�=�G�= E�=kٻ=��=\��=���=�s�=X�=���=��=/�=d== �n��R��C�,��   �   l/��qsؾ<��A�y1p��k��4��Lʱ��ǻ��:���ѻ�f豿_s���Վ��fq�ƈC�:I�i�޾M���pF��]��M����Ͳ<�#=��M=�Ra=NQf=��b=ȧ[=��S=��M=^�J=H�K=F�Q=��\=B�m=b>�=	j�=��=�۲=�<�=���= ��=*]�=���=�	�=��=��=1��=$.
=@o���Q���1��   �   �����Ծ�2��S>�n�k����l���î��������V���خ�����M���m���?��R��پ�Ж��MA���۽(IB�`����*�<&�&=�N=�_=yb=�a\=CR=N�G=6g>=�W8=��6=�,:=��C=0T=��j=t�=�G�=E�=�ٻ=��=v��=���= t�=��=$��=�=�/�=2?=��n�Q���,��   �   `�����Ǿ��	�64��_�d���8W�������Q��؅��oI����uf�����H`��65�й�6�̾�����h2�Jƽd*#� (M9,��<$�.=�IP=t�Z=�<V=�H=�55=D0!= �=���<D��<��<���<�X=@y=�\<=J�c=���=eE�=��=,f�=2d�=��=���=�Y�=yս=�ɐ=��=01�s���   �   ��n�H賾NK����#�,L�i�r�,����,���ˠ��������h��~�����r��_L��$�z���y�����y��*�����S� �
<�,=N:=Q=(�P=��?=��#=��=4�<�l<�I�; �y:�?+�@kY���X�@��;�e<$�<H� =�w\=���=vj�=l;�=�	�=XV�=��=���==��=��*= ���T�s�vn��   �   ̗J�e(��'�پq}��c3�zV�q�t�܌��a@���֐�	���C��wDt���U��3��w���ھ�7���Q�S���-s��U�PQ�<H+=*�E=&N=�>=6�=���<��R< �Ӻ@0�����X%���D��CS��SN�Z5��d����� �����<<=��i=��=X��=���=���=Ȧ�=풓=��>=s<�0��-��   �   �="��~��i������r�lt5�kP�$e�TUr�?�v���q��5d��O��Z4��k�;L�<g����~���$�M���6H��3r;���<�7=�M=�D=
�=$��<`J�;p]��5�jn��7��MǽB��z��z���ȽP ��_�1� n��t�<��>=pۄ=�ڞ=:�=Jק=���=�Q=X��<(�̼Wث��   �   �~HF�z����w������z�n�)��$;��7F�+�I���E��:�K7(�����Q�DཾK����:A��e콦�f�؏6���<�'=�O=�+P=
 0=�[�<�^�;�ϙ���F�ym����轏����0��$F�G�R���U��~M�tT;��� �D@���E����W��"��ЙV<��=@ho=er�=iw�=�I�=l�`=�j�<�	�0,e��   �   :y�����&X�F�������}Q�
L�� ����mi�`���X�-�����獾JqL�#�]����]��xLQ<8�=@�P=�?`="�I=�=X$V<�l���nU��뾽�O�)�<��j�d������?M���᤾<���L��Ú��(<Y��w(��\�>P��p� ��;z�=�(^=��=�=*i=��=б <$/��   �   &:��a���7�!�T������zCľǫپ羔�NK徺(־�$��3h���z����C�$��"&���<𼰽�;ж=��T=��r=�<i=��8=��<�;ͻ,:��f���:�P�T�9"����FGľ�پ��i �/P�y-־.)��Al��.~����C���.���U� q�;��=v�T=d�r=�:i=~�8= ��<�ͻ�   �   �b��LgU�E澽&L���<�Pj�,�����RI���ݤ����H�����Y5Y��q(�LR��G���T��S�;��=�.^=	�=o�=R+i=V�=Щ <�7�|���V*X��Ó����徚S�lN�#����+l���P[��1�ȃ���ꍾ�vL��'�X��� s��X,Q<n�=@�P=�=`=j�I= �=�/V<�   �   @}�;�Ù�@�F��g�������ʝ0�F���R�%�U�
xM��M;��� �65���;����W����V<��=2oo=�t�=<y�=K�=F�`=xi�<@⻞0e���KF�N���Iz�������{���)�x';�B:F��I�r�E�u:��9(���PV��㽾V����?A�m�*�f�`�6�Dܪ<��'=��N=�*P=L 0=�_�<�   �   ���<�n�;@�\��,�(�m�1��Eǽ*�⽨�H�"���Ƚָ���t_�`� ȶ��2�<�>=߄=�ݞ=�<�=�ا=l��=x�Q=��<��̼lګ�H?"���~��k��O��Vt�@v5��P��	e�Xr��v���q��8d��O�`]4��m�P�_j����~���$�<���Q���q;,��<��7=X�M=�D=&�=�   �   �=��<��R<�Ӻ������h%�2�D�J5S�TDN���4��U���� q�@�<X=�i=���=4��=���=7��= ��=���=�>=�q<��0�W/�.�J�s)����پu~�He3�V�_�t������A��ؐ�a��ME��Gt� �U�3��y�ͭھ:����Q��X��H6s�ؽU��G�<(=2�E=LN=�>=�   �   ��?=��#=��=���<@1l<���; �{: �*� �X���U��ߣ; 0e<T)�<�� =�\=x�=�m�=>�=��=X�=\��=���=���=��*=@����s��n�v�n� 鳾`L����#�*L���r�見�}-���̠�0����������������r��aL���$�>�������g�y��-����`�(�
<x)=2:=Q=��P=�   �   �<V=tH=�75=�2!=|�=H��<p��<���<0��<x_=�=�c<=Ξc=���=!H�=	�=Kh�=f�=l��=���=�Z�=Rֽ={ʐ=��=h-��s��~���<�Ǿ��	��4���_������W��{����R������EJ��~�Qg����uJ`�@85�����̾{���k2��Mƽ�/#� DI9���<.�.=�HP=��Z=�   �   �xb=�a\=�CR=,�G=�h>=�Y8=��6=b/:=��C=dT=*�j=$�=dI�=�F�= ۻ=U��=���=���=u�=p�=���=��=d0�=�@=��n�P��v�,�����\Ծ�2��S>�{�k���m��9Į�j���W���М��ٮ�����_N���m���?�dS�o�پ�і��OA�r�۽.MB��ũ�$&�<z�&=��N=D�_=�   �   p��<lY�<���<h��<�>
=�(=T4=�.N=k=��=[��=Q0�=fB�=tS�=$��=0?�=�+�=^>b�>1� >���=r��=�n�=B�v=�d�<����Ľ̉7��k���l˾��8P)�]�J���h����N���U;������w)����h��~K��}*�°��Ѿ����>O�����Y���U ������QF<�ح<���<���<�   �   �S�<Н�</�<�\�<h� =<=��%=��==F-Y=vrw=s6�=(�=�u�=�6�=�\�=���=���=l��=t >dY�=�=N�=#��=��x=\�<��⼋a��`
3��P���QǾ�<��%&��G��fd�(�{��5���Ň�f:���{�Z�d���G�f6'����ש̾|K����I��y��$���I���(�}_<�̷<�'�<T��<�   �   ��<l��<��<�ſ<0��<<��<th�<�V=jO"=f
>=Zv^=n��=ՠ�=Z��=M�=4��=2��=0��=:��=���=���= o�=͡�=f=Td�<P���u���&�}Y��5r��Lg��\��\M<�g9X�uFn�tf|�4����Z|��?n�|QX�/�<�ڲ�n���忾xH���:����6*t�dߴ�@�>;�Փ<��<��<�X�<�   �   �R�<hϱ<� �<�e<��<<��(<H7-<�L<��<��<�"�<Xa!=��N=�2�==��=�=��=��=`
�=pK�=L��=��=W	�=�΃=�B�<�MZ�����Z���j���������~+�2E��|Y��wf���j�aNf�9;Y���D�e+�����e�� �� Yu�N|"�)��"�;�9�0d;<p��<���<�}=���<�   �   |�<�z�<���;��8�P����c��뒼�U���P���e�0�л�S�;�P�<f
=��E=�=(�=��=q�=���=�<�=���=�߱=��=�=`4�"�]��H��IH�F���B�ľ�0���5�i-��?���J�8nN��DJ���>�>\,������- ľ�͒���M���3C���� d;�f�<� =v(=�,=HQ�<�   �   ��< ��;�T������:��x�C�0�k����3p���
����d��s2�i߼�K��L<�=��W=���=�j�=��=��=�ֿ=�3�=��=X�/=k<��������!���p�Ҧ����оמ������E!�{+��J.�1�*��] �`������y�;R렾7�l��!��½n:�H�����<�S=7+=b/=`�=`��<�   �   2<0�ĔQ��#������n�ὦ.��b ����
���i�ؽ�����kw��c��뾻t��<~n1="=���=�t�=�ׯ=�.�=���=��C=0K�<V������Xv��|�<����!P���n˾;���p��n
����ú	�V����P�ƾ�١���x�E�1�h��pt�(�����R<�
= �<=�M=��C=n�"=@c�<�   �    ֺ�����k�-F��vy��n����5���I���U��tW���N�',<�85!�42 ������n[�t���@9;<��=f'h=YĎ=�D�=#=�=rw�=�~Q=0_�<@���#�g׭��S��qD��u�FE�������eɾJ�վ5`پ%�Ӿ��žt�k����n�L�1��������4�˼��<�	=�J=vyj=��k=(~Q=�s=�<�   �   �ט�p.\�\<���m�1U8�ptc�<���*i���\�����h���:)����y��iO��b �`�)���~Ҽd�;a=v�W=96�=�+�=JF�=�HV=��=s5<ʘ� %\�6���i�hP8��nc�����e��5Y����������&����y��dO�t^ �� ό����mҼ���;�e=ްW=U7�=:,�=GF�=�GV=��=�`5<�   �   ��#��ܭ��W�2vD�z{�}H�������iɾF�վ1dپ��Ӿ)�ž����)��1�n��1�q��|���غ˼�<�	=x}J=�wj=(�k=�~Q=�u=��<�aպh�弮�k��?���q��̥�p�5�(�I���U��nW��N��&<�U0!��- ������b[�@{��8W;<L�=�+h=�Ŏ=vE�=w=�=*w�=�|Q=�W�<�g��   �   3����|����<�%��,S��{r˾���r��p
���ʼ	�5�U��1�ƾ�ۡ���x�D�1��彤wt�\�����R<X�
=0�<=�M=��C=��"=h�<�!2<H����^Q�^��(����Ὅ%������������ؽ�y���]w��W�@������<�t1=�&=���=v�=�د=�.�=��=��C=XB�<\c���   �   �����!��p�x�����оp�������G!��+��L.�6�*��_ �������ž;&��l��!�.�½":� ����<�Q=�5+=�a/=��=\��<�<���;�%��0������"�C�R�k�� ���h��0����d��e2��O߼����L<�=f�W=V=�l�=P�=��=�ֿ=b3�=��=<�/=HW<����   �   �M�QMH�b���مľ�3��>7�M-��?���J�/pN�FJ�^�>��],�H������!ľ�Β�V�M�f��#E����� B;�c�<�=�'=�,=S�<�<Ā�<��; `7�0e��ic�tؒ��@��h:����d���л���;�c�<�=^�E=!�=���=t��=�r�=���==�=Ԉ�=*߱=��=~�= b4�~�]��   �   ���j��� �j��a�+��3E��~Y�Lyf���j��Of��<Y���D�f+�����f㾸��BZu�0}"�a*����;�x9��_;<���<���<v}=���<@U�<Tӱ<�&�<�)e<��<<)<(R-<�M<���<�ȴ<�2�<�h!=h�N=�5�=☙=Z�=��=��=`�=L�=���=��=��=�̓=�;�<�aZ�-����   �   �&��Z���s��=i��w���N<��:X��Gn��g|�͟���[|�r@n�@RX�Ȥ<�N�����忾�H��C�:���彶*t�$഼��>;pՓ<���<�<�Y�<D�<��<��<�ʿ<���<���<q�<�[=rT"=�>=\{^=ʛ�=���=E��=�N�=���=L��= ��=���=��=���=�n�='��=@=�]�<X%���x���   �   �3��Q��SǾ�=�G&&��G��gd���{�G6���Ň��:��d�{���d���G�u6'������̾VK��`�I�]y��#���G��(��~_<�ͷ<�(�<\��<XU�<���<�1�<�_�<>� =T!=֟%=(�==�/Y= uw=�7�=F�=�v�=�7�=�]�=j��=d��=���=� >XY�=��=��=p��=��x=���<��d���   �   ֊7�l���m˾e���P)���J��h����\���V;������^)����h�4~K�1}*�f��6Ѿ{����=O�"��aX���S ��s�� WF<�ڭ<H�<���<���<�Z�<��<���<~?
=)=�4=N/N=Pk=��=a��=<0�=JB�=LS�=���=�>�=B+�=9>7�>� >N��=���=6n�=�v=4`�<󼦝Ľ�   �   �
3�Q���QǾ�<�v%&��G��fd�ʐ{��5��:Ň�	:��7�{���d���G��5'�?����̾tJ���I�Aw���!���B��(�(�_<|ѷ<d,�<���<�X�<��<�4�<�b�<�� =t"=ؠ%=��==�0Y=�uw=�7�=w�=�v�=�7�=�]�=���=���=���=� >�Y�= �=8�==�x=��<���#b���   �   �&�4Y���q���f������L<��8X��En�de|������Y|�4>n�-PX��<����k���㿾G����:����\$t��մ��?;Lݓ<$��<�<T`�<�
�<d��<��<Tп<���<P��<�t�<2]=�U"=�>=8|^=*��=L��=���=�N�=���=���=@��=��=B��=>��=�o�=��=�=de�<���2u���   �   [���j�3�����B���}+��0E�t{Y�vf�M�j��Lf�}9Y���D��c+����3c������Uu��y"��$���;���8��x;<���<���<Z�=`��<H^�<ܱ<�.�<�8e<0�<<@)<�\-<`M<\��<�˴<5�<�i!=:�N=26�=0��=��=�=F�=��=�L�=<��=���=
�=�σ=(F�<�DZ�2����   �   �E�HH��󑾘�ľ�.��>4��	-��?�ܐJ�>lN��BJ���>�OZ,�?��{��mľA˒�ȾM���_>����@�;�r�<R&=.=�2=d^�<$�<D��< >�; @6��T��[c�DҒ��;�� 6����d�p�л ��;�e�<�="�E=z�=��=㩹=s�=���=�=�=���=��=:�=έ= �3���]��   �   Z|��0�!���p�ण�,�о��������C!�o+�]H.��*��[ �V������#�;u蠾q�l��!���½N�9����䦒<Z=J=+=vh/=P�=� �<��<p�;����P���.��8�C���k�+����g��;��H�d��d2��M߼���L<�=<�W=�=bm�=��=ܖ�=*ؿ=/5�=j�=2�/=�}<ڳ��   �   ]���q��*�<�����M���k˾ɒ��n��l
������	�2���羡�ƾH֡�&�x���1����^dt��y����R<h=<=��M=��C=4�"=�t�<@:2<���z�NQ���,���^��%$���n�������ؽy���\w��V�P���d��<�u1=�'=U��=w�=�ٯ=h0�=���=�C= V�<�H���   �   �#��ѭ��P�|mD��p�[B������&bɾR�վ\پ�Ӿ��ž�ﯾ�����n��1�Ֆ�ò����˼�<�	=V�J=Z�j=��k=��Q=&|=h�<@�Ժ@��p�k�H=��bo��ڤ���5�|�I�2�U�|nW���N�s&<�0!��- �����a[��y���Z;<^�= -h=�Ǝ=�F�=;?�=�y�=��Q=�j�< ���   �   ����h\��/���e��K8�xic����mb���U��ً��I���s"��	�y��^O�
Y �2���􅽰SҼ���;�n=��W=�:�=�/�=�I�=2OV=��=Љ5<4����\��3���h�nO8�nc�����}e���X��[���ײ���%����y�tdO�F^ �* �V���4lҼП�;g=��W=�8�=�-�=�H�=�MV=��=��5<�   �   �XԺ���¬k��8��Fi����|5�T�I���U��hW���N�� <��*!��( �*����R[��_��8�;<��=�3h=gɎ=�H�=�@�=�z�=L�Q=�i�< ��ܵ#�)խ��R��pD�u��D�������eɾ�վ`پ�Ӿ��ž\�V��o�n� �1�:�𽔹��X�˼ �<(	= �J=\|j=��k=ڃQ=�{=��<�   �   @2<H���o��P�>����������~��|�+���r�ؽp��6Lw�H�p/��࿥<�~1=6/=6�=Ny�=�ۯ=�1�=T��=��C=TT�<�M������zt����<�:���O���n˾����p��n
������	�K���@�ƾy١���x��1�� pt�@�����R<��
=p�<=��M=��C=�"=�t�<�   �   T��<�,�;���x�������C���k������`������<�d��U2�`1߼���M<�=��W=eƎ=Tp�=Z�=���=�ٿ=(6�=��=b�/=�y<6��w~����!��p�����P�о��������E!�l+�yJ.�(�*��] �Y������k�;B렾�l��!���½� :���d��<�U=�9+=f/=��=���<�   �   $�<l��<pP�;�P5��?��@c������(��P!����d�P;л
�;{�<�=�E=c�=q��=���=Zu�=p��=h?�="��=��=��=�=��3�x�]��G�pIH�����ľn0��o5�Z-��?���J�0nN��DJ���>�:\,������" ľ�͒�n�M�����B��H���t;�i�<�"=t+=1=t\�<�   �   l]�<�ܱ<@1�<Be<��<<00)<�r-<P6M<̴�<T۴<�D�<�q!=��N=�9�=p��=�=��=d�=��=N�=j��=v��=�
�=-Ѓ=4G�<PEZ���������j�����������~+�2E��|Y��wf���j�\Nf�6;Y���D�e+�����e�� ���Xu�7|"��(����;��9��h;<���< ��<��=���<�   �   t	�< ��<��<�ҿ<p�<���<�{�<6a=>Z"=r>=D�^=���=���=܌�=Q�=���=4��=���=H��=T��=$��=Dp�=¢�==\g�<���u���&�^Y��r��4g��R��RM<�a9X�pFn�pf|�2����Z|��?n�{QX�,�<�ٲ�i��~忾qH����:�p���)t�\޴���>;�ד<���<�	�<�]�<�   �   `W�<��<\4�<$c�<"� =x#=:�%=��==�2Y=�ww=9�=��=x�=9�=�^�=���=n��=���=� >>Z�=��=��=���=x�x=��<@��?a��>
3��P���QǾ�<�~%&��G��fd�%�{��5���Ň�f:����{�Z�d���G�e6'����ԩ̾yK����I��y���#��I� �(��~_<4η<�)�<���<�   �   `���P���0���@i� ��98�C<HC�<��=DOP=���=H��=��=ֻ�=^��=\�=,T�=�>:�>�Z	>��>�p>d"�=(f�= u�=*{U=��c<�(�m)½<�*�����𮾬�߾���FC��9.�"9���<�{.9��`.����ۨ����6���=��| D�Z���Ϋ�PtQ��.���;�� ��D����蜼hȳ��   �    ��܂���\���� � ����-<h��<`=�D=@sw=,�=�d�=b_�=���=p��=���=��> $>^�>�>�>�=^��=¥�="�W= �u<����s����&��tz��^����۾�?�RD�A�*�J�5��X9���5��+������Z4޾� ���	����>��l�!���BF�8�弈r��H{^� l�P!���ͦ��   �   4̕�����ǁ�p -� wE����;�G�<X��<V�!=P�P=7�=�V�=���=7��=Fl�=|��=�B�=�� >��>8>��=���=P,�=p�=g]=��<H�����2�m�j�0���ξR��"���e!�^�+�B/��|+�JU!�������о�����w��/�_��v����%�����`_3��������8%H�t���   �   @X�@�z� @x��YO��l� q�.�;p<��<�=��:=|^i=n��=Fv�=E�=��=
��=<��=�m�=8��=<
�=85�=���=7��=��d=<�<8����E���'	�h'R��7�������� �-��w���������6�R��'E�zL��W���N�Z�����Ž�Wf�L��8�&�@���@��: ƣ��`������   �   p6��PGO�4��8j��\���Tq���3� ����:�Q&<�3�<�y= �7=��n=P��=�]�=�F�=���=�*�=du�=��=|[�=���=��="�k=���<�.��^j��]���3�I�z��`��xJƾ�\�p���J��t�
�
���(��BG�ľ�e����x���5�i��^���8D��C�@;v;��;<��T<�N&<��;��Ժ�   �   @S�pTA��$����Ӽ����K��S�L���<��$���hf��\��@P<�o�<�s8=��y=\��=��=@��=�w�=�K�={�=�(�=��=�6o=�=�f�� �*�y��8�&�O�T ��0���������վ�W�
�羽�� 0ӾT¼��ߠ�$��NF��C�qҲ�p�>�x�|�`^�;��<�\�<�!�<�}�< 0k<0D�;�   �   �Np��Mf� Z޼ �"�<�Q��<z��-��Z{��1�������r��H;�ا������8<F�=\�O=�=�=���=L��=��=R+�=�ԯ=��=r4l=�=���;�߼OA����-$�*@W�PC�����-����������~��8ᦾ����Cy�j�E����n�����X�TE�� 
�;P�<T6=�"$=6O=~�=�h�<�@<�   �    ��x���$�j�u�������ƽ���	���M~��������#ν�>���we��-�� �x��4�<B,=��r==Nz�=�L�=X4�=�p�=P�`=b0=�,Q<Hfx� �A��⩽�����#�
�I�1�j��G��8쉾䈋�Ԇ�8Yx�tY��2�o��EV��:KY����Pg<�A�<�J7=̯V=�,]=��M=,=TW�<0sy<�   �   0[ֻ�d�p�����%���)��F;�� E� �E���<�^�*�'��(�v�����9��=h��6W<Z!=81U=Bm�=� �=GL�=F�w=�8K=�e=�!�<Bֻ��{p�Ч�����	��)�dB;���D�;�E���<��*����!�c�����9��h�@QW<�&=�5U= o�=["�=^M�=Ɯw=�9K=�e=��<�   �   �wx�~�A�<穽� ����#�T�I�k��J��������ֆ�8^x��Y��2�����[���SY�(����P<�8�<�F7=��V=`*]=��M=�,=<V�<Xuy<����q��X$���u�������ƽ���f���Bz�������콄ν�7��nke�����9x�0C�<8,=P�r=ڲ�=�{�=�M�=%5�=.q�=L�`=D/=�"Q<�   �   �#߼*E����X0$�:DW��E��y�����������l����㦾A���Vy�ԘE��������̥X��P��`��;��<3=
 $=�L=��=@f�<0@<�p�(Ef��R޼j�"���Q��3z� (��Ju������j�����q�<;��뼰��P"9<��=��O=G@�=���=恵=��=8,�=bկ=4��=�3l= = l�;�   �   H +�������O�t"������\�����վ�Z��羚�ᾥ2Ӿ�ļ��ᠾ�%���PF��E��ղ���>�h�|�0B�;���<�V�<��<4y�<H)k<0<�;�S�pPA�  ���~Ӽ<����D�tK����(��tv��@�e� "�XeP<P��<�z8=��y=軚=��=���=&y�=�L�=�{�=")�=��=�5o=�= 짺�   �   ej�&b潼�3���z�c���Lƾ�_�@������ړ
�]��4+��]I��ľ5g��O�x���5�-�������G���C�`v;��;<(�T<F&<0֛;��Ժp;��8FO����<e����� Aq��q3��յ����:�p&< C�<�=�7=�n=��=�_�=�H�=\��=�+�=Zv�=���=�[�=���=(�=h�k=��<�.��   �   �H���)	�*R��9������!"�f�����������7�*���F㾘M��5�����Z������ŽZf������&� ��� ��: ���@m��X��@X���z��=x�hSO� c�@��N�;0+p<���<��=&�:=�ci=馌=�x�=G�=��=p��=X��=�n�=ئ�=�
�=X5�=t��=���=��d=�5�<@����   �   ��� ���j������ξ�S�����f!�G�+�/�H}+��U!�(������i�о����2�w���/��� ��� �%�l����c3�P ��H��h)H���T͕�,��<ǁ��-��]E� ��;�L�<���<��!=��P=��=�X�=p��=���=�m�=���=tC�=/� >�>A8>��=t��=�+�=��=�d]=��<����   �   .v���&�Bvz��_����۾[@��D���*�Ѧ5�PY9�]�5��+�9�����r4޾� ���	����>�vl�� ��nBF���弈r���{^�0l��!��Φ�(�������[���� � �����-<`��<=��D=uw=�=�e�="`�=J��= ��=��=��>$>j�>�>؜>��=���=��=4�W=Щu<���   �   �*½�*�����4�߾���{C��9.�""9���<�j.9�x`.�a�����3�⾰��=����C�����ͫ�xrQ��+��X9��@���p眼@ǳ�T���0�������f� G�9X�C<4D�<��=�OP=���=S��=
��=û�=8��=�[�=�S�=�>�>rZ	>��>�p>�!�=�e�=vt�=|yU=x�c<+��   �   [t����&��tz��^���۾�?�#D���*��5�gX9�w�5�+�p��5��?3޾������v�>�ck����z?F�t��xm���q^�H�k�����Ȧ�H���}��HW��@� � �����-<@��<:=��D=�uw=b�=�e�=U`�=p��=$��=@��=��>*$>{�>0�>��>�=J��=���=��W= �u<F���   �   ������j����p�ξ%Q�����e!���+�c/��{+�UT!����N��� �о����w���/���꽢���D�%�0��� P3��������(H�����Õ�����h���H-��"E����;XR�<��<��!=Z�P=��="Y�=���=���=�m�=���=�C�=M� >�>g8>�=��=�,�=��=�g]=h�<���   �   D���&	��%R��6���	��r�� �-��X�����e���5����B�pJ������E�Z�.���|Ž�Pf�h���&��"�� ��: ^���7�������W��z�%x��<O��N��x躠m�;�7p<���<��=֖:=*ei=u��=�x�=nG�=��=���=���=,o�=F��=*�=6�=|��=��=��d=�@�<�����   �   XYj��Z���3���z�[_���Hƾ�Z���������
�����%��yD侊�þuc���x���5��������f<��dC� �v;��;<�T<�e&<��;��Ӻ����8'O������W�������+q��_3�@���@^�:�z&< G�<��=Z�7=�n=���=^`�=FI�=���=R,�=�v�=B��=�\�=ۍ�=��=0�k=��<��-��   �   ��*�w����"�O�������&�����վ�T��~羔���,Ӿb��� ݠ��!���IF�@��̲���>�8e|�p��;��<(i�<�.�<Ȋ�<�Lk<Ђ�;��R��.A�(�� pӼ�����>��F����!�� q��h�e�@���jP<���<�{8=��y=W��=�=c��=�y�=`M�=�|�=�*�=���=�:o="= ����   �   �	߼�<��b��)$�M<W�A��D��\�����֏��d{��ަ����y���E�ۜ�y����X��1���L�;$#�< ==v)$=�U=��=lx�<06@<��m��"f�tB޼�"�
�Q��-z��%��:s������
����q�P:;��� ��x&9<��=~�O=�@�=��=���=��=J-�=�֯=2��=$9l=b=���;�   �   �Ex�x�A�ݩ�<���,�#���I�<�j�8E��R鉾酋�ц�gSx��Y��2�����N��>Y��}��(�<@R�<�Q7=��V=�3]=��M=z,=�g�<H�y< ��Ta���
$���u������ƽh��r���ty�]�����콯ν 7��Zje����`+x��D�<,=Z�r=t��=�|�=�N�=�6�=s�=��`=Z6=�HQ<�   �   ��ջ^�pp�a�������H�)�h=;���D�χE�V�<���*�-����j����t9���g�XzW<|/=4=U=wr�=�%�=�P�=��w= AK= n=�1�< ֻp�tp�����
��Ԧ)��A;�A�D���E�I�<���*����!�������9��h��TW<�'=�6U=�o�=M#�=�N�=\�w=~>K=&l=D0�<�   �   @��@_���$���u�����g�ƽ��佚����u�>���r��u�ͽ)/���[e����� vw�pX�<P,=6�r=T��=�~�=�P�=C8�=}t�=��`=�7=�IQ<�Jx�f�A��ߩ����ƺ#���I�L�j��G���뉾�����ӆ��Xx�2Y��2�;���U��xJY�d����j<�C�<�K7=��V=:/]=��M=^,=�b�<�y<�   �    /n��"f�D?޼��"���Q��&z�!���m��쉔�~x���q��,;�dt�h\�hQ9<,�=��O=8D�=��=���=��=/�=:د=H��=�:l=$=0��; ߼�>��<��+$� ?W��B��q�����ܦ��˒��i~��ᦾ����y�>�E�Ƞ�����X��C����;��<�7=�$$=�Q=�=|r�<�-@<�   �   ��R��1A�,��lӼ�����9��?��d���\����e� ��X�P<|��<��8=L�y=���=��=���=�{�=O�=!~�=�+�=���=<o=�=�ɦ�j�*�E��3�:�O����ن��S���Y�վ�W��羢���/Ӿ?¼��ߠ��#���MF�C�"Ҳ�δ>���|��e�;<��<�_�<8&�<l��<�?k<�n�;�   �    ��H,O�h��� V������q��L3� ���@7�:��&<�V�<��=�7=.�n=ٛ�=Qc�=�K�= �=@.�=�x�=���=�]�=Ԏ�=��=6�k=���<x�-� [j�!\�&�3���z��`��9Jƾ�\�I���:��h�
� ���(��4G�ľ�e����x���5�-������C� }C� Iv;x�;<�T<�W&< ��;�
Ժ�   �   ��W���z��'x�(<O�pJ��6����;pGp<���<��=R�:=�ji=-��=�{�=�I�=�=���=\��=�p�=���=B�=7�=L��=®�=��d=�A�<ĝ���D��&'	��&R��7���
������ ���l���������6�M��!E�qL��O���<�Z����׀Ž6Wf�H�优�&�@���@�: ��� O������   �   dǕ����� ���p-��E����;�U�<���<d�!=� Q=K�=�Z�=���=���=do�=>��=�D�=�� >��>�8>��=���=b-�=p��=�h]=H�<Ȇ������j�
����ξ�Q�����e!�X�+�>/�|+�GU!���������о�����w���/�?��R�����%����� ]3���������H�����   �   �������X��0� � ���H�-<`��<$=��D=Hww=.�=�f�=6a�=V��= ��=��=[�>�$>��>z�>:�>��=���=>��=�W=��u<£��s��t�&�ntz��^����۾�?�ND�@�*�I�5��X9���5��+������Y4޾� ���	����>��l�� ���BF�Ф� r���y^�@l�����˦��   �   4�н�Sʽf��Tq��@f��g���G���(<R�=n�R=n�=L�=:t�=�s�=�P�=�>ɿ>JN>��>.1>��>���=L��=��=�A�=De?=�$?<`:��x,��Ҿ��M�W_����ƾfHݾ5쾨^�6G���ݾ�Ǿ���k����u]��'����V��a����X���Q��Ai���q��
M���ʽ�   �   E�ʽŽ��8���&b���x�L��l<4��<��K=��=��=�0�=6N�= i�=^8>�$>��
>mS>�">L�>:�=�w�=*0�=��=�<@=H�J<�򼗱��A~
���I�ю������¾_�ؾ$v�h�pv�j�ؾY�¾�W���u����W�ve"��뽙���j�x�h�L��F���]�j���lڜ�	�jĽ�   �   ;ҹ�Q�����fA��r�W�܄
��a`� ��;�y�<�6=��{=.�=�'�=f��=���=��=�J>O�>H�>��>�>�U�=�r�= O�=&��=NB=�j<p�Ҽ�򔽷/���<�H�z�2���Ɲ��̾�پ�e޾��پ��˾r���{d�������G����M�Խ_ܔ��U��+�l&��<�rde��ފ�򙡽]`���   �   z'���~������.���зJ��"
�4����:|�<|=��P=Ҳ�=6��=���=�I�=�)�=6!�=���=g3>
>> ,�=��=L6�=�ܼ=!��=�C=L��<������sQ�ΰ)��b��r���䤾�6���ľ=�Ⱦ�þ����pq��AX��<Mb���.��D��"����k��Y�tb����`}��n/��^�"u���ߖ��   �   �)��턽����g���@�j������� ��;0�<$^=��J=C��=d\�=f��=<��=�v�=~��=���=��=��=8��=��=)�=m�=�7@=���<�i�RX�U�Ľ�O���C��Ms��Ԏ��v���穾{��񌨾�᜾�T����k��<�0���Eɽ�D�����������S�X�E�P@���kּM��E��Oj��   �   �TA��UT�TZ��<S�ޘA�� '��"�D���x�A� r980Y<���<0)=�c=�Í=gK�=^�=�=2e�=z.�=`��=-�=�w�=��=�6�=PW6=l�< ����-��\������"�EVJ��2m�� ���d��l|��L���a���`��;�6�r�Խ���!���A��� �;���;@��:����������!��   �   z�� �%���=�VM�nnS��_Q��F�Z�3��������������,S<@��<d	8=z�u=�ѕ=���=]Ǻ=d��=a��=CL�=oͫ=b��=N�l=t^"=�ϔ<�Ի����[��AĽ��� �!��<�WQ���\�|�^��U��mC�K�(�
��,ͽ�5����y?����;���<8f�<ą�<ԗ�<�?< �V:<3�x���   �   4G������2��2Z���{��Ί�\���2q�����Mρ��5Y��> ��&����v���{<�.
=XcM=�A�=MM�=(��=� �=�y�=��=D"z=��C=F�=ؼZ< -滰a�x�V�������̽w���^��<P�5$�dO#��U�X�	��D�󉰽�Zn� r�������~w<d��<��&=$�8=�P5=*�=P��<?�<���;���   �   pT=��":��~�g���8��΅ѽ�߽���;Lܽ�ɽv쪽�׃�ܜ-�觝� W;d��<��%=6HY=�y=�x�=��}=��e=��?==$է<<�;8W=��鼼:�~~�:����4��ɀѽI�߽Z���Eܽ�ɽl檽D҃��-����� ~W;��<�%=�LY=y=�z�=��}=8�e=��?=$=Dڧ<�J�;�   �   p1��e�h�V�������̽����_���S��8$�S#�Y���	�K�e���^dn����0滻�gw<`��<N�&=�8=dL5=�=P��<h7�< ��;0���J��V��2�0Z�z�{��ˊ�m����l���	���Ɂ��*Y�Z4 �����Dv�X�{<x5
=iM=fD�=sO�=��=��=H{�=Z�=�$z=�C=��=��Z<�   �   �,Ի��r^���DĽ^����!�w�<�
Q���\�r�^���U�bqC���(�����ͽ�9��b��?� ��;��<�]�<8}�< ��<��?< �U:pL3����T����%���=�6M��kS�~[Q�>�F�P{3�(����ἴ����X��LS<�	�<�8=�u=.ԕ=���=0ɺ=��=���=�M�=�Ϋ=Z��=��l=_"=�Δ<�   �   �����-��_��"�n�"�bYJ�D6m��"���f��p~��<��me�)�`�{;����M�Խ>�$��*���̼��ߺ;���;@m�:� ���������!�XA�XT��Z�=S���A���&��������A� �x9KY<���<F6)=֐c=:ƍ=�M�=W�=� �=�f�=�/�=���=&�=fx�=l�=�6�=W6=��<�   �    �i��VX���Ľ�Q�d�C��Ps�k֎��x���驾a������N㜾qV���k�)�<�ޖ�gHɽ�F����������S�8�E�$H���sּFQ� E��Sj��+��x���fg���@�lh�P���Ș���;�'�<&c=��J=���=�^�=d��=��=0x�=���=���=��=��=���=�=o�=d�=�6@=Љ�<�   �   ����p���T�ز)�d b�t��V椾�8����ľڈȾ��þ�����r��9Y���Nb�D�.��F�������k��\��gＤ�弈��0r/�t^��v���ᖽ)��B�������������J��!
����� ��:d$�<�=6�P=���=ꦢ=���=�J�=�*�=L"�=��=�3>\>>�,�=F��=�6�=�ܼ=Ԩ�=VC=���<�   �   �Ҽ����&1���<�S�z�U�������E̾)�پ�f޾ʃپ��˾6���e�������G�*��)�Խݔ���U���+�(&�0�<��fe��ߊ�<����a��`ӹ�A��Ƹ���A����W�t�
��]`� ��;�}�<(�6=�{=9/�=�(�=h��=���=Ƙ�=K>��>��>��>>�U�=�r�=�N�=���=�B=�j<�   �   <�`���X
��I�����ȁ���¾#�ؾ�v����v���ؾ��¾�W���u����W�ne"��뽃���t�x���L���F���]������ڜ���kĽ��ʽzŽ[��18���&b�n�пL�p<\��<� L=<�=R�={1�=�N�=`i�=�8>�$>��
>zS>�">G�>�9�=�w�=�/�=��=B;@=��J<�   �   �>���-�������M��_��慨Hƾ�Hݾ$5쾬^�G�̖ݾ�Ǿ[�����Lu]�1'�y��U�������X���Q��@i�W�9���L��޵ʽ��н�Sʽ�e��q���f�g���G�@�(<��=��R=��=L�=3t�=�s�=�P�=�>��>3N>��>1>l�>���=��=J�=FA�=�c?=h?<�   �   �򼭱��D~
���I�����ր���¾��ؾ�u��~쾵u羟�ؾ��¾�V��u��J�W�7d"���뽾���V�x���L���F���]�D���Dٜ��쳽�iĽ��ʽ�Ž�	���6���#b���x�L�w<(��<�L=��=��=�1�=�N�=�i�=�8>�$>��
>�S>�">^�>,:�=�w�=00�=��=�<@=��J<�   �   �Ҽ��/��<�>�z���������
̾нپd޾m�پb�˾$���?c�������G����=�Խ�ٔ�p�U��+�x&�H�<�t`e�y܊�����^���Ϲ�� ��s����>���W��
��M`����;��<N�6=��{=�/�=H)�=ʪ�=��=��=1K>��>��>��>4>\V�=*s�=�O�=���=�B=�j<�   �   �������N�N�)� b��q���㤾�5���ľ��ȾM�þ�����o���V��bJb�x�.�v@��]��<�k�(T��WＨ��<x�ti/�>^�r���ܖ�$��d{�����u���V�J�N
����� ��:�+�<�=��P=���=���=��=nK�=X+�=�"�=8��=�3>�>>-�=��=N7�= ޼=I��=HC=@��<�   �   ��i�&LX���Ľ�M�V�C��Js�ӎ�u���婾t�������ߜ�S����k���<�V���@ɽV@��~��8���x�S�`�E�4���^ּ6F��E��Gj��%���脽��:�f�|�@��`��񶼨��p3�;�.�<�e=ЯJ=���=G_�=���=��=�x�=6��=`��=�=x��=���=��=��=%�=�;@=���<�   �   k�T�-��X������"�SJ�/m�����b��6z�����]�ؘ`��;��{�g�Խ�鋽����� ]���6�;���;�̡:@�����lz��!�.KA�|KT���Y�2S���A�F�&���������A� v|9hWY<���<,8)=V�c=�ƍ=9N�=��=,!�=&g�=L0�=*��=��=vy�=��=�8�=Z\6=��<�   �   ��ӻ��V���;Ľ�����!�J�<�4Q�W�\���^���U�liC�-�(�B��Yͽ�/����hT?��"�;|�<8t�<���<襦<��?<��X:�3�X�*�� �%���=�M��aS��RQ���F�8u3�0�����`z��`1�`TS<��<8=,�u=�ԕ=��=�ɺ=���=|��=hN�=�ϫ=�=��l=|d"=,ݔ<�   �    �� O�(�V�󂜽��̽}������.L��0$�K#�6Q�*�	�"=�ł��Nn�4[���_��8�w<,��<�&=�8=VW5=@�=t��<xO�<�<�; L뻬1����|2�f%Z���{��Ǌ�禒��i��-��ȁ��'Y�2 ��� .v��{<�6
=�iM=�D�=�O�=���=M�=|�=k�=�'z=�C=�=(�Z<�   �   �3=�d��&�9���}������-���yѽ��߽z���=ܽ�ɽ�ު�˃�΅-��~���&X;���<R�%=fTY=�y=~�=�}=f=P�?=,=$�<`��;�(=�X��.�9���}������0���}ѽ��߽9��"DܽPɽ_媽rу���-�`��� �W;Й�<��%=�MY=y=Q{�=�}=* f=��?=�=��<�|�;�   �   �8������2��$Z���{�tŊ�ȣ���e������Y��& �������u�8|<�>
=VqM=H�=�R�=2�=��=T~�=��=�+z=��C=|�=��Z<��� N�B�V�u����̽4������O�$4$��N#��T���	�>D�d���Zn�Tp��Щ�� �w<��<��&=F�8=�Q5=�=���<XE�<0�;�n��   �   z��~�%��=��M��`S�PQ�x�F�6o3����Pu��h��@��hwS<d�<�8=�u=�ו=Վ�=*̺=���=���=QP�=�ѫ=�Ĕ=��l=g"= �<��ӻZ��W���=Ľd����!���<�kQ���\��^���U�omC��(�����ͽu5��� �(v?� ��;X��<h�<��<���<��?< �W:�-3� ����   �   �OA�rOT���Y��3S��A���&����}���vA� N�98rY<|��<?)=��c=�ɍ=Q�=^"�=r#�=2i�="2�=���=��=�z�=<�=:�=f^6=��<Xi�"�-��Y����"�4UJ��1m�X ���d��3|�� ���a�Ĝ`��;�
�"�Խ�
�D �� -����; ��;��:��������X����!��   �   (���ꄽ���p�f���@�T`��x�0P�;�7�<�j=��J=��=�a�=T��=���=�z�=��=��=��=ڍ�=���=.�=��=,�=L=@=���<��i�MX���Ľ�N�РC��Ls�[Ԏ��v���穾S��ь���᜾�T��q�k���<���kEɽcD����������S���E��>�� iּvK��E��Lj��   �   0&��=}����������ʱJ��
�����@��:h0�<�=��P=P��=y��=���=2M�=�,�=$$�=���=�4>?>(.�=��=H8�=�޼=��=�C= ��<`���2	���O��)�Ib�Tr���䤾�6���ľ"�Ⱦ��þw���bq��5X��'Mb��.��D�����v�k��Y��a���弾|��m/��^�bt���ޖ��   �   jѹ�<�������?����W�`�
��M`����;`��<�6=��{=1�=t*�=���=��=(��=�K>+�>�>P�>�>W�=�s�=HP�=u��=�B= j<��Ҽ~�4/�p�<���z���������̾վپ�e޾��پ��˾j���td�������G����0�Խ@ܔ�̿U�±+�&���<��ce�*ފ�|����_���   �   ��ʽ�Žk
��D7���$b�����L�8w<���<�L=�=4�=Q2�=|O�=.j�=�8>%> �
>�S>#>��>�:�=vx�=�0�='�= >@=H�J<,����~
�n�I�����퀥��¾S�ؾv�^�jv�f�ؾU�¾�W���u����W�oe"��뽅���P�x�P�L��F���]�M���Eڜ����jĽ�   �   ��a��>\��L���2������ݽ���L:�`GB��z�<�Y=��=��=d��=|��=�\>_�
>�,>=U>�>FI
> �>��=z��=�&�=s�="�5=0�p<������m��̽����L<��-b����*���l��b͉����b�d���B�h��*��R�ý� ���G������;���Q�ɽ���c��b6��M� ]\��   �   ڎ\��IW���G�/�����Gٽ�*���C���:�(M�<J�U=-�=2o�=��=��=_>V	>� >4>��>(	>D�>d��=���=E�=)��=p4=Ѐq<P���p}h��ǽ���Y8�>c]��z�ۼ���𪆾)�z��G_�D�=�;��d0�֖��������~N��8��F�½[���=)�61� �G�W��   �   ހM�	I�A�:��$�<�V�̽���J�	� F5�4�<��K=�C�=5ڵ=���=� �=�K�=��>�j	>�
>ƈ	>�>�)�=\��=�4�=�i�=1��=�.=��p<�L��x�Y�݁����(	-�(�O�R�j��,|��䀾:{��i��O��
/�$r� ܽ@�۞��vd��bh��
������p�ݽ�g	�*L#�N9�T�G��   �   �^6��53�e+'��{�I��+ƥy�� ���_�,�<b�8=BO�=���=P�=�(�=���=S�=�?> �>D�>V��=�2�=��=���=R�=l�~=jO#=PDd<H~~�DE�f���SD�����:���R�T�a�2�e��<_�oN��5��
����괷�,���l�K�lq+��w/��)V�9��B���뽶���+"��c0��   �   ����S�J�F"���pսJ��x-c�<w��P����Z�<v|=\�e=�g�=R~�=V��=a�=���=.��=��=��=$<�=(��=$k�=u�=�ו=�c=T�=��;<�`p��0�ڕ���ӽ6d��!���4�l�@�v>C��7<�0k,�|��B���bǽ��p��FI<������~ż�̼�q	��F�4��������佮j����   �   �|��,x��H��j�ս����E���&T�8]�h�=�`��;x��<~k0=��p=�\�=���=dE�=��=���=�=&/�=|*�=�-�=���=r��=� ~=t�9=�<���;�����#�t��ȵ��7�,��m��?�����p������kD���ւ�4�)�d���HW#�@Mu� ���F��Iм�v/�L��'�����ʽτ��   �   �ѵ�Yj��5��P诽�p��������S�v���ӱ��_ŻD <L��<p�&=$�a=͡�=IF�=�γ=�a�=nk�=���=/�=a�=��=h1{=��@=�� =`�n<� L�D����<$� Ep�􈜽U��Q#ؽ*n꽲��S��0ܽ���������`�N�
�0m�@k�:h'N<���<6�<�$,<�V���߅���	���Q�2Љ��<���   �   �x�����*�������X���,��8�g��C���$�μ�A���6;�q�<�=B�A=��t=4��=(�=P�=�=�w�=MX�=��b=��-=0��<�3T<�>�,����� ���7�d�j��ߋ��h��ꢫ���� Y������=̑�$�k��'���� `����G<(��<��=�+"=\=B�=Б�<8�<P7�����������M��   �   �����?���a��t{�6���M��u����ꃽ��p���M�>^�(ͼ���; $�<r�=�G=��g=f�v=��s=r=_=~#;="�
=��<`�;0�#��uļ��n�?��a��u{��5��EL��@����烽��p�J�M�xV��ͼ���`A�;x0�< �=2�G=��g=�v=P�s=fB_=�(;=ę
=��<0�;@�#�Hjļ�   �   D���.� ���7�8�j�����k��ᥫ����C]������Б�ֵk���'�ذ�������iG<P��<��='"=R	=�}=P��<P�<�l�����������M�x�t"���,��뢑�$Y��H,��z�g�ړC���� �μH�@� B7;`~�<��=�B=��t=|��=�*�=R�=��=�y�=�Z�=|�b=��-=4��<�FT<����   �     L�����d=$�fGp������W���&ؽir�]���W��5ܽ6���叚���`�*�
�XHm� ��:N<���<�+�<�,< ���셼��	���Q�ԉ�{@��lյ��m�����"꯽�q��ㆅ�L�S�ج�\̱��;ŻX <���<��&= �a=��=kH�=�г=�c�=>m�=V��=�0�=�b�=w�=X5{=��@=�� =дn<�   �   `��;������#�,���ʵ��:�1��������0�s����/H��ڂ���)�����xj#���u�@<��G��Uмd}/�n��������ʽʈ�u����{��+�뽣�ս���F��v&T��[���=�0��;���<~o0=��p=�^�=���=G�=���=��=t�=�0�=�+�=T/�=��=穜=�~=��9=d�<�   �   ��;<`fp���0�ܕ���ӽ�e�� !���4�̰@��@C�:<�Xm,�j������Mʽ�'s���M<�����Ȇż��̼dv	�j�F�4���W���E�佑l�{����:U��K��$��4rս@��$.c�Dv�� ���0_�<=P�e=+i�=��=���=Tb�=6��=R��=��=�=<=�=<��=2l�=
v�=�ؕ=�c=��=�   �   H@d<�~�VE�����G�X��֫:���R�l�a�@�e��>_��pN�s�5�<����ض��܎����K��t+�0{/��-V�`������>��*-"�(e0�`6��63��,'��|����%ﹽ��y��� ���_���<,�8=FP�=���=T�=�)�=���=�S�=J@>��>��>��=P3�=>�=���=��=��~=6O#=�   �   h�p<Q��~�Y�у�����
-���O���j�{.|�z倾�;{�$�i��O�f/��r�4ܽ:�˟��^d��dh�������2�ݽ�h	�FM#�v9��G��M�	I�-�:��$����̽��V�	��>5���<��K=�D�=�ڵ=J��=X�=$L�=Ǖ>�j	>=�
>��	>�><*�=���=�4�=
j�=��=2�.=�   �   �zq<d���
�h���ǽ����Z8�Ad]��z�R����E�����z��G_���=�^���0�򖼽$���I���N������½.����)��61���G��W�n�\�(JW���G�b/����(Hٽ�*���C� �:�TN�<��U=��=�o�=P��=��=|>$V	>� >)4>��>(	>H�>b��=n��=�D�=̔�=`4=�   �   �p<�����m��̽��pM<�.b���>���o��T͉�����d�d�B����)��}�ý����'G��@���諢��ɽ���T��Z6��M��\\���a��>\��L���2����d�ݽ����9�@@B��{�<�Y=��=��=`��=n��=�\>R�
>�,>'U>�>+I
>ݳ>8�= ��=*&�=��=Ȩ5=�   �   �q<����}h�ͷǽ����Y8��b]�Z�z�~���&p����z�rF_�,�=�.��r.����m������;M�����½����(�^51�8�G�?W���\��HW���G�*/����GFٽ')��DA���:��Q�<4�U=��=�o�=���=�=�>5V	>� >84>��> (	>]�>���=���=8E�=U��=�4=�   �   `�p<H����Y�[�����-��O���j�X+|��〾T8{��i���N��/��p�.�۽������$d��^h��������;�ݽSf	��J#��9���G�FM�jI���:�D$���z�̽��z�	�  5��<�K=�E�=�۵=���=��=xL�=�>�j	>\�
>�	>;�>�*�=��=�5�=�j�=��=ܤ.=�   �   �Sd<Hm~��E�����SA����:�{�R��a���e�Z:_��lN���5������G���≇�~�K��k+�rr/�Z$V�d��7���������)"�ma0��\6�D33�()'�\y���3깽b�y�<� �`�_����<|�8=�Q�=���=�=*�=��=XT�=v@>��>̛>v��=�3�=��=b��=��=��~=�R#=�   �    <<�Hp�P�0�\֕���ӽ�a��!���4���@��;C��4<�^h,����?����½�sl���A<������qż��̼Lk	�d�F��������K��Lh�	����P�ZG����^kս\��8$c�f���o���i�<�=`�e=Uj�=���=f��=�b�=���=���=�=l�=�=�=ʳ�=�l�=w�=�ٕ=hc=p�=�   �   ���;����d�#�� ��@õ�d2�^��v��"����pm����	�
?���т�N�)�@w���9#���t�pޕ��F�;м�n/�v��V���|�ʽ,��v��"r��+��]�ս���N@���T�S�0�=� ��;��<�r0=V�p=�_�=>��=�G�=%��=���=��=1�=z,�=�/�=䋵=���=j~=|�9=,�<�   �   ��K�4���$3$��:p�}���AO��<ؽ�g�1��zL�*ܽ\�������@�`�`�
�m��q�:�EN<��<D�<�A,<�`���΅���	���Q��ʉ��6���˵��c������᯽j��o���f�S���ཱ�pŻ j <���<:�&=�a=ޤ�=I�=`ѳ=!d�=�m�=Ӫ�=n1�=�c�=H�=�7{=x�@=Ԏ =��n<�   �   �~��R� ��7�2�j��ً��b����������R��'����ő�
�k�|t'���������G<��<�=
3"=N=p�=���<8<�����ƽ�0�M�X�w�^��9$������R��%&���g�J�C����$�μ��@�@w7;|��<��=8B=��t= ��=+�=�R�=���=�z�=;[�=�b=��-=���<pUT<@���   �   H��l�?���a�j{��/��2F�����pჽ��p��M��J�0�̼Pl�p��;PB�<.�=��G=��g=�w=��s=2I_=�/;=��
=8�<@a�;hk#��Sļ����?�\�a�Xg{�/���F�������ヽ��p�H�M��R���̼���`O�;L3�<*�=(�G=��g=��v=6�s=`C_=�);=4�
=�
�<�)�;��#��aļ�   �   �x�����&�����9S��\&����g�4�C�4��إμ8�@�@�7;`��<��=�B=��t=���=�-�=.U�=��=}�=�]�=��b=��-=���<�mT<�Q��t��$� ��7�ڴj��ً�d��О�����cV��n����ʑ���k��}'�𞹼PV��ЅG<���<~�=�,"=*=*�=ܓ�<P�<�)��@�������M��   �   �ϵ��g�����]䯽�k��V���t�S�J��������Ļ�} <x��<��&=��a=���=�K�=�ӳ=rf�=�o�=��=�3�=�e�=��=r<{=r�@=ȓ =0�n<�YK�$��d1$��:p�C����P���ؽ]k�n��9Q�/ܽ����ʊ��ֻ`�B�
��,m� ��:P*N<��<l7�<�',< :���݅�B�	� �Q��Ή�;���   �   {��$v�����D�ս�	���A���T��R�x�=� �;�
�<�v0=��p=�a�=j��=�I�=&��=x��=��=�2�=V.�=�1�=ڍ�=���=x
~=j�9=P �< ��;������#�D��]ĵ�k4����R��Z����p�D��8��C��\ւ�z�)�����T#��Cu�P��h�F�`Hмv/�:��s�����ʽ����   �    ���R�I�����mս���&c�g���j���l�<p�=>�e=�k�=]��=��=�d�=4��=D��=~�=��=6?�=X��=n�=�x�=eە=vc=&�=�<< Cp���0��֕� �ӽ�b��!���4���@��=C�X7<��j,�@������ǽ�Wp���H<������}ż0�̼,q	���F�豋�����%��Xj���   �   �^6��43��*'��z�C
���빽z�y�2� � �_���<�8=�R�=���=B�=B+�=@��=�U�=A>8�>]�>���=�4�=�=���=�=�~=U#=�Zd<�h~�<E����HB����>�:���R��a���e�~<_��nN���5��
�f�񽹴�������K�q+�jw/�\)V�������뽊��T+"�8c0��   �   ��M��I�Կ:�T$���ه̽�����	��5���<��K=F�=Aܵ=���=��=<M�=K�>Gk	>��
>�	>��>p+�=���=m6�=�k�=��=��.=P�p<�E��D�Y�h���
��-���O���j��,|��䀾�9{�ςi��O�|
/�r���۽ �����6d��bh��
��|���I�ݽng	�L#�*9�"�G��   �   ��\��IW�V�G��/�E��*Gٽ�)��B�`�:�PQ�<b�U=:�=4p�=���=l�=�>lV	>� >s4>��>c(	>��>4��=Z��=�E�=��=:4=��q<􊛼�{h�X�ǽ����Y8�
c]�±z�ʼ���媆��z��G_�;�=�0��R0�Ŗ��� ��oN��.��0�½C���0)�61���G��W��   �   ��Ⱦ�ľ����$죾�늾��]��c$��ٽ�Xg���L�pa�<Jmf=>֦=Qb�=H�=?> f	>ft>X�>#e>B�	>��>�W�=n1�=:)�=��=���=
 6=H�< `c��	��\Ki�OV����׽\���	����	�������߽�꼽�꛽�����o��~�Q-��K]ͽ�5
��T6���g��]��e㤾����ľ�   �   b�ľu���������`��MY��� �ܤԽ�`��2>����<.�e=!��=��=�|�=H1>�l>4e>̀>�>�R>iH>���=��=���=���=��= 1=p'�<@x���ge�H���l(ӽ�}���e��
������ؽy��4����z��/d�Pr������ƽ��$m1�6b�����=�����d���   �   ����Fʴ��$���閾j��)L���(;ƽ1N��B�\�<�d=''�=~��=��=���=�j>� 	>l�	>�>��>���=�y�=��=*��=s��=�p=�F!=,�<0ǣ�$６[�ְ����Žf��3T��W�������ὅ�ý::����Z�V���A�~O�A災�����r-#���Q���������Ƞ��Dp���   �   �	���Ţ�@n�������f�
�7�yn�f˰��b3�`)��h��<2�^=6��=��=D��=�/�=�- >�u>��>VL>D��=t]�=d��=���=fi�=�[�= �M=|A=8.R< � ��;�=N�����&s����̽��۽�i޽NIԽ J��}Ǣ��C����K�������x��z�H��菽�xͽ*����7�>�c�I8��Wۖ�4塾�   �   W����@��c����ak�o�G��8�B꽈嗽z�@�=�Դ�<�S=L�=K��=��=���=���=�k�=���=���=��=���=�Ž=v�=�1�=��X=v�=t�< ��;p]������D�w��[p��r2��Ad��:Ѷ������%���Vs�&8���Ph��d���<��� ��$)K��ǜ�/�,��R>���b�xw��0����   �   yi��f�!�Y��KC��Q&��&�$�Ľ`3�(����|���F�<�E?=�w�="e�=�c�=�e�=Dg�=^z�=���=P��=e�=�ϲ=@ �=�_�=<G=N�=Tʞ<@ٜ;���T��h(��F�`�o����ᓑ��O��o��84z��|M����H>����7��r��>; �� ���Լ��J�d�����㽜E��N4�	�N��Fa��   �   (�4��p4�R�+�Ð������ؽ܅���W�\Eܼ�E8���<d�=be=��=ڙ�=K��=k�=� �=�F�=�=�e�=׊=fH^=ԥ!=�%�<؞<�|�������6����l?���X��-j�er��p���a��G�~c ��=༐Uj�@���hJ&<ȳ�<0�<�6�<�QW<���4�>�;��Ɩ��nѽzM�����:,��   �   ����+�t�p��ѽ(ޮ������?���ݼ����)<`��<��/=tHg=��=(C�=\2�=*9�=��=)ڍ=��n=<?5=̃�<�83< K˻H���v����A�4�c��y�*���eA��P�x��Zf���K���)�
���[���BȻ�h�;���<T�<2�=�y/=2�+=��=�T�<�
�;8�[��}��yy��ޫ�M�Խ3��   �   [C��v���X���;����������o�<;����F��@�"���J<�k�<�%"=z;N=�n=@�~=:�}=F�i=@C=�a=��<����P����-���u�����QH�����\��?���������o�;;�L��h?�� �"� K<�t�<�)"=�?N=@n=��~=�}=X�i=�EC=h=���< I��>����-���u�k����   �   ��A��c��y���@����x��[f��K�8�)�����e���kȻ0@�;���<��<v�=4u/=:�+=Z�=tH�<p��;��[�ֆ��y�'䫽1�Խ�8󽓿�w.���\��ѽ$஽���ڔ?�X�ݼ���ȋ)<X��<��/=DLg=��=E�=\4�=@;�=:�=�܍=Z�n=�E5=��< X3<�˻������   �   ԁ���,�ִ��i?��X�<.j�:gr�p�$�a�� G��h ��H�Xkj��>��x6&<��<|��<�,�<�;W<����������;�r˖�tѽ|P���*>,�X�4��s4��+���r��W�ؽ{�����W�dEܼ`38���<��=He=6�=s��==�l�=^�=�H�=��=Dh�=�ي=XN^=@�!=$3�<�<�G���   �    ��;�����~'�rF�Np����	���CR���q���9z�:�M�*���H����7������; �ĸh%��Լ��J����]��ZH��Q4�D�N��Ia�X|i�2�f��Y�<NC��S&�b(�'�Ľ�5����� s��I�<�G?=y�=Vf�=2e�=�f�=�h�=�{�=f��=��=g�=�Ѳ=�"�=5b�=<AG=h�=�Ӟ<�   �   �
�<�̄;� ]����� �D����8r���4���f���Ӷ�Y����(���[s��*8�<���p������ȹ������.K��ʜ��2�n���T>���b��x����嬎�VB������dk�T�G�n:�,D��旽�� �=����<:�S=��=*��=֢�=���=� �=�l�=*��=X��=!�=9��=fǽ=�w�=�3�=L Y=��=�   �   �B=�0R<�� ��=�"?N�m���u��ȶ̽Z�۽2l޽�KԽ]L���ɢ��E���K�������� �H�H�%돽�{ͽ���t�7�l�c�~9���ܖ��桾�
��Ǣ�co�����H�f�M�7�eo��̰��c3��,�����<��^=���=���=���=�0�=\. >v>�>�L>H��=�^�=���=��=�j�=�\�=��M=�   �   <G!=��<Pͣ��&Ｒ[�/���U�Ž*��V��*���w��]��ýk;������N�V���A��O��聽� ����.#��Q�i���{�������<q������-˴��%��\ꖾ���	L���� <ƽ2N�(D�L\�<�d=u'�=���=R��=��=k>� 	>��	><>��>n��=^z�=Ʊ�=̇�=��=`p=�   �   �1=�%�<@$x���Xie�O����)ӽ�~��rf�Y
�H����c�ؽ���z���2z�j0d�r�����ƽS��m1��6b����g>��Z���d��ݸľ�u������V������fMY�!� �+�ԽD�`�p2>���<|�e=L��=��=�|�=_1>�l>Je>�>�>	S>�H>���= ��=܏�=���=���=�   �   �6=��<@uc�t���Li��V��\�׽�\��*�	�����	�������߽i꼽Y꛽	����o��~�	-��#]ͽ�5
��T6���g��]��i㤾����ľ��Ⱦ�ľ����죾o늾��]��c$�ĳٽ�Wg���L�4b�<�mf=L֦=Vb�=F�==>�e	>[t>H�>e>/�	>r�>�W�=*1�=�(�="�=?��=�   �   � 1=)�<�x���|fe������'ӽ�|��^e�>
�.��
��b�ؽ ��Å���z�L-d��r�Z����ƽ>��l1�P5b���x=��W���c��ɷľ{t������k������LY��� �O�ԽR�`�P)>���<��e=���=�=D}�=z1>�l>\e>�>�>S>�H>��=Z��=,��=���=x��=�   �   �I!= �<P�����2[������ŽE���Q������G��R�ý�7�����V���A��	O�Q偽�����4,#��Q�М������ʟ��7o��w���(ɴ��#���薾{��fL�u��r8ƽ`,N��2�c�<td=e(�=���=ڊ�=v��=4k>� 	>��	>W>��>���=�z�=0��=V��=���=Dp=�   �   :F=�AR<�� �1（7N����p��a�̽��۽bf޽�EԽ�F��?Ģ��@����K������h��F�H� 揽�uͽn����7� �c�
7���ٖ��㡾��<Ģ��l��&���f���7�Xl��ǰ�"\3�����<�<l�^=	��=���=���=01�=�. >Cv>�>�L>���=�^�=��=���=Wk�=�]�=v�M=�   �   ��< ��;��\�H����D����Ol��N.��	`��Ͷ�h����!��DOs��8�*���[��4���8�������"K��Ü��*����^O>���b��u��r�������?������H^k�B�G�6��<�����`��U=�4��<x�S=���=[��=���=:��= �=$m�=���=���=~!�=���=�ǽ=�x�=�4�=�Y=ʈ=�   �   ��;8��@��$��F���o�+������J��Lj���*z��sM�P���.��Xg7��� �; �����X�Լ��J�����Q�㽪B��K4�t�N��Ba�ui��f�6�Y�HC�eN&��#�G�Ľ�(�t����r��hU�<ZL?=�z�=�g�=.f�=�g�=8i�=J|�=���=v��=rg�=pҲ=7#�=�b�=2CG=�=�ڞ<�   �   y��t!����0a?���X��"j�\Zr��p�D�a�hG��Y � +��2j������h&<���<��<8D�< nW< �}��߫��~;�<����hѽ!J���7,��4��l4�K�+�،������ؽ�����W��0ܼ@�7���<��=�e=��=w��=���=hm�=��=YI�=���=�h�=6ڊ=�O^=ʭ!=7�<��<�,���   �   ��A�Аc�B
y��z��V;����x�@Of���K��)�����hH����ǻp��;x��<$*�<.�=��/=ި+=�=�c�<@L�;x�[�.s��my�
ث�,�Խh+󽸸��'�x����@�ѽ$׮�!��z�?�p�ݼ���(�)<���<��/=�Ng=��=�E�=�4�=�;�=��=ݍ=<�n=�F5=p��<�]3<p�ʻ�������   �   xA������U��Q8��6��������o��/;��~�H+�� "� /K<��<�1"=�FN=�n= �~=>�}=��i=�LC=�o=�	�<����(����-�N�u�Y��;������-Q��z4��B�������o��/;�0��1�� A"��K<{�<b,"=�AN=�n=Н~=֜}=2�i=�FC=�h=@��<�8��;���-�X�u������   �   ޻��*�*�M����ѽ�ٮ����ډ?���ݼа�0�)<���<0=.Sg=�=H�=J7�=)>�==�=�ߍ=f�n=�M5=ģ�<�3<`�ʻ}��(����A�F�c��y�x��49���x��Nf���K�ȅ)�����<R�� %ȻP�;ȟ�<��<l�=�z/=�+=��=8V�<��;�[��|�rxy��ݫ�W�Խ�1��   �   ��4�
p4�J�+�v����/�ؽ΁��.�W�T2ܼ �7�	�<H�=� e=H�=J��=���=fo�=��=�K�==[k�=*݊=V^=޴!=0F�<��<P0j�� �<���\?�6�X��!j�[r�Tp���a�DG�j_ ��7�@Lj� `���O&<쵗<��<48�<�TW<�X����;�5Ɩ�nѽ0M�^��h:,��   �   �xi�w�f�R�Y��JC��P&�~%��Ľ8,������~���V�< N?=�{�=�h�=�g�=.i�=�j�= ~�=���=r��=�i�=�Բ=�%�=�e�=FIG=@�= �< L�;Ȟ����0�
F���o��������M���l���0z�zM�����;��x�7��d��I; ܹ�����Լ�J����5��mE��N4���N�0Fa��   �   ,����@������`k���G��7��?��◽���e=�`��<Z�S=^��=J��=ͤ�=j��=h�=zn�=��=P��=@#�=���=ʽ=�z�=�6�=�Y=��=��<��;��\�P���:�D����Jm���/��5b���϶�Y���%���Us�%8���g��`���D���`���(K�Zǜ��.����Q>���b�`w������   �   u	���Ţ�n��O���f�J�7��m�tɰ��^3������<��^=u��=T��=h��=2�=
/ >�v>��>�M>���=b`�=���=N��=#m�=�_�=��M=~I=(MR<؄ �X.�7N�[����p��ײ̽��۽�h޽rHԽ{I��Ǣ�OC��
�K���V��"��(�H��菽�xͽ��x�7�(�c�<8��Fۖ�塾�   �   ~���/ʴ��$���閾���L�x���9ƽf.N�P7��a�<�d=�(�=���=R��=��=�k><!	>(�	>�>p�>���=�{�=`��=���=��=�p= L!=0�<����pＰ[�)���O�Ž@��QS������;��n�=�ý�9������V���A�LO�'災��� ��f-#�s�Q�������������8p���   �   Y�ľu�������H���LY��� �F�ԽĿ`��,>�� �<��e=���=G�=~}�=�1>�l>�e>*�>3>[S>�H>���=��=��=ǟ�=R��=�"1=\,�<��w����ee�r����'ӽ9}���e��
��������ؽ]������z��/d�.r�v����ƽ��m1�6b�����=�����d���   �   �n!�++�!��g��?��:߼�b'��-QR����G���8�����<<�|=�u�=�m�=���=KM>20
>�>�%
>+V>J� >���=܋�=Xl�=N²=��=.y=�<=���<(am<�7������8f�p���~5��a=�
�5��X#��2����p�\4�2�D�ō��XF�D�$�GLe�b엾����,0�����)��   �   �S�Q!����UM�8��-������M�^���`�m�
�<z~=-J�=t��=~F�=v>�	>�A
>�>\p>���=F�=�C�=S��=J�=�+�=��n=,P3=TW�<�W< �������~�$�/��6���-��C� ���༰�׼���9��3��߯ڽVB �1�_��v��;��F���0�����   �   Q��S�/�	�ʕ���Ծv*���a���R@��]��z�w�0�+���<i��=���=7�=Xd�=`�>��>�.>�>�g�=P��=�D�=�/�=JԳ=쨛=>�=�QN=dy=~�<��<0��pʊ��߼tY�:=�`!!�0z�&N �`�ϼ�n��0���(vǼ�z�dy��Ľ1���O��l�������fվ�g��{X	�|4��   �   �K����S���R�ƶ��<T��k�q���+���׽\P�����q=���=ڊ�=j�=�Z�=�x�=h >@z�=(��=���= +�=x!�=�=Ԑ�=�{=n_H=��=���<��H<�s=:��"��[��܃ټ�z �*��zb�(���ֱ�@�z�()�P�PoV���ͼ&B?�������	S5���u�sX���˿�� ߾GN���[��   �   6뾮�澧�ؾ�#þGq���\���P�����=��r� ���;p�=kT�=�l�=���=$��=��=ph�=�j�=,��=�=� �=�Р=���=��W=��"=X��<�d�<� �;����p�G�xv����ż������;޼�Y���1�� �#���7�`�1;Pi�;@��:��d���k���Ž�����M�7��x��dn����־���   �   ˤþvO���񴾄���������b�jw,�L��V�����0#<@�=Z2�=5�={�=���=bH�=��=x��=�t�=�+�=�I�=\�`=��!=L��<��&<`���U�T���t��x� �jl��_�H� ��O㼰/���7v���ջ !!;�R1<Ť<x�<�-�<�h<pq�����$툽�߽�!��nV�iƅ�q���>���v����   �   ��J똾93���ہ��^���4�\��GQ���KV�X�����Y<y=0�t=��=��=7�=���=,��=@��=T�=&�u=��0=�R�<��;�mD�.�j\)��WQ���i�Is���n�8�^�,E���#����l~��8A�`�G;��j<�?�<Z�=��=�=��<x�i<P��<���s����s]�xL��t�O���J���   �   *^h�$�f�<�Z�?�E���)���	�bн�����(��a~<^v=n_=+8�=�Ý=~ަ=��=nS�=ô�=��Q=�G=X:<`�@����T�i��`������q�˽��ҽ��νh������V���Tf^�<��̢�� o���{)<p��<��=2f;=�dQ=:T=΢@=�-=�K�<�Ŕ��

�!����iӽ v��10���K��=_��   �   �&"��#�l/�d|����� ʽ�\����O��+��갻Uo<��=d�?=�Qm=3.�=MM�=��=Ri=�2=l��< �:��Ҽ�6`�������qe�=��*"��#��2�u����cʽX_��N�O�(/༐찻�Xo<��=��?=�Tm=�/�=*O�=��=.Wi=&2=��<@/�:�Ҽ�*`�,������ra�"��   �   ��˽��ҽ��ν|������l���pb^�*��ġ��@u���t)<���<�=�b;=aQ=�5T= �@=(=�>�<P��
�ؿ��2pӽ�y��50�R�K�KB_��bh���f�P�Z�әE���)���	��н��������a~<dw=�o_=Q9�=0ŝ=$�=��=�U�=t��=2�Q=^O=(C:<�@�*����i�>Z�����   �   �LQ���i�>@s�l�n�|�^�.�D�n�#���p���G�`[G;�j<(9�<ޡ=��=r=T��< ~i<0��z���x�����`��L���t����0M������혾r5���݁�9�^�J�4�`��"T��~OV�<��� �Y<ty=V�t=��=��=��=���=�=���=�=��u=�0=�c�<���;0DD�P�\Q)��   �   ��T�x箼���D� ��h��]�b� ��P�p2��x@v��	ֻ � ;�E1<@Ō<��<@%�<V<`���n��8񈽂߽�"!�WrV�tȅ������������V�þ�Q���������K�����b��y,�d��j�������<�=�2�=�5�=�{�=��=�I�=L�=V��=�v�=).�=�L�=0�`=:"=���<�'<�
��   �   Hp�<�J�; ���0�G�(r����ż���<���?޼�^��87��X�#�@8��i1; N�;@H�:��T���k���Ž�����M��Å��z���p����־s�徂8������ؾ�%þ�r��@^��"�P����?���� ���;�=�T�=Lm�=<��=��=��=�i�=Hl�=���=�=��=UӠ=���=��W=�"=���<�   �   ~�=,��<�H< �=: �"��[��\�ټ"| ����d�8�� ܱ�ȶz��)�`�X{V�l�ͼFF?�z
������T5�
�u��Y��lͿ�]"߾8P���\��L�����T��eT�"���WU��$�q�0�+�w�׽�P����\q=���=��=��=v[�=�y�=� >@{�=d��=
��=�,�=L#�=﫮=蒖=�{=�cH=�   �   �SN={=l��<�<���`ˊ��߼�Z��>�B#!�|�P ���ϼr������zǼ8}�gy�ҟĽY��DO��m������	hվi��1Y	�85��Q�XT�ӆ	�����Ծ<+��xb���S@�6_����w�x�+�L��<j��=ƈ�=N7�=�d�=��>��>"/>F�>dh�=T��=�E�=�0�=�ճ=*��=j	�=�   �   ��n=�P3=�W�<�W< �4���漒�@�/��6�x�-��D����,��׼����9�C4��ΰڽ�B ���_�w���򻾑G�"�����W��S��!�L���M���ᾆ��%��F�M�M^�X��@�m�
�<�~=BJ�=���=�F�=+v>�	>�A
>@�>�p>d��=��=D�=���=��=V,�=�   �   ny=8�<=���<�]m< V�������g� ���~5��a=���5��X#�J2�|��d��3���D�����VF�P�$�^Le�n엾*����30����)��n!�"+���X����߼�B'���PR����򤍽4���ؤ�<l�|=�u�=�m�=���=HM>+0
>�>�%
>V>6� >f��=���=l�=²=���=�   �   p�n=�Q3=Z�<( W<@���������h�/�� 6���-��A�����༰�׼ ���9��2��Ӯڽ�A ���_�!v����[F�s������)S�� �����L�x�ᾂ��N���M�B]������m���<�~=�J�=��=�F�=@v>		>�A
>J�>�p>���=��=@D�=���=�=�,�=�   �   HUN="}=h��<�<����Ê�\	߼�U��9��!��v��J �p�ϼ�g�������oǼ�w��`y��Ľ��~O��k�������eվ}f���W	��3�YP��R�m�	�\�����ԾK)���`��,Q@�0[��֥w� �+���<���=���=�7�=,e�=��>%�>@/>^�>�h�=���=F�=;1�=�ճ=���=

�=�   �   ¤=ػ�<�H<��>: x"�8P��lxټu ����(]�����̱�0�z���(�����]V���ͼZ=?�:�����&Q5�d�u�W��>ʿ��߾VL���Z��J����Q���P�����R����q���+���׽�O��╻"v=� �=d��=���=$\�=z�=
 >�{�=���=R��=
-�=�#�=R��=m��=!{=@eH=�   �   �u�<�d�;�|���G�0f��,�ż\��d���-޼�L���$����#� �7���1;Г�;�f�:`|����p�k�!�Žf��.�M�����w��Hl��/�־��徔3�&��3�ؾT!þ+o��[���P�����8���� ��/;��=�V�=�n�=Z��=̜�=���=j�=�l�=8��=_�=:�=�Ӡ=���=�W=~�"=���<�   �   �T�D஼��� �,b�V��� �H>���Xv���ջ@�!;�l1<x،<0��<89�<Ѐ<�=������舽߽�!�BkV�_ą�(�������ˌ���þ�L��1﴾���M�����b��s,�8��,�������@<|�=5�=h7�=2}�=���=^J�=��=���=w�=�.�=M�=�`=B"=8��<X'< ���   �   JQ�N�i��;s���n��^���D���#������k������G;��j<`M�<��=��=�=���<P�i<�z⻀���n�����Y�T	L�j�t�����G��>
���蘾�0��2ف�>�^�p�4�����J���@V��⌼ЩY<�=&�t=|�=&�=��=L��=��=���=p�=d�u=��0=�e�<P�; ?D���(O)��   �   S�˽��ҽظνު������ж��ZZ^�@��؎���&��؜)<���<��=�l;=�jQ=,@T=�@=@4=�Z�< ���x 
�7����bӽ,r�,-0���K�x8_��Xh�դf��Z�T�E�m�)�f�	�н<������ ����~<�}=pt_=
;�=rƝ=�=� �=3V�=᷆=��Q=P=F:<��@�4��P�i�pY�����   �   U&"�#�|.�9{���B�ɽ�X����O�t�ࢰ��yo<
�=��?=�Zm=�2�=R�=�
�=�]i="-2=D��<@\�: �Ҽ`�퐫�o��]�l�""��#��*��w�U�����ɽ�U��:�O��ༀ���xwo<`�= �?=�Wm=�0�=P�=H�= Xi=�&2=p��<�D�:��Ҽ�)`����� ��a����   �   �]h���f�p�Z�@�E���)��	�3н%��r����� �~<�~=(v_=A<�=�ǝ=��=�"�=�X�=���=��Q=�W=`j:<�@�d��Rxi�vR��w鸽#�˽��ҽ~�νG���V���3���@U^�6��P����(��Ȗ)<���<��=�h;=�fQ=�;T=��@=v.=M�<�����	
�ӹ��5iӽ�u�`10���K�>=_��   �   ���똾�2��Vہ��^�|�4�
��XN���EV�茼0�Y<�=.�t=^�=V�=��=��=��=d��=C�=��u=��0=8w�< R�;�D����TC)�L>Q�"�i��1s��n���^�D�D�r�#�,���tk���#�@�G;��j<F�<��=|�=�=��<��i<�⻮��ns����R]�QL���t�3���J���   �   ��þLO����4���6���کb�_v,����ϐ��h�Ἐ9<��=<5�=�7�=~�=��=�K�=~�=���=fy�=C1�=>P�=2�`=:"=���<='<`Q�@�T��ή���� � ��\�fR�ʸ ��<�p ���v���ջ�X!;0]1< Ќ<,�<�/�<�k<�l��R���숽P߽�!��nV�Zƅ�b���+���\����   �   	6뾑��}�ؾk#þ q���\��V�P�����;��Z� � ;��=�V�=2o�=��=���=���=dk�=<n�=��=��=��=�֠=��=��W=��"=���<���<p��;�M��p�G��^��H�ż�༌��00޼�P���*����#�@�7��1;pq�;�֬:���h�鼞�k���Ž�����M�,��x��Zn��t�־ ���   �   �K�����R���R྘���T����q�P�+�]�׽l P���u=� �=���= ��=�\�=�z�=� >�|�=��=���=�.�=�%�=���=ꕖ=:&{=|jH=ک=P��< �H< �?:�m"��L��4wټ~u ����<_� ��ӱ���z�)�X�8mV���ͼ�A?���������R5���u�lX���˿�� ߾@N���[��   �   Q��S�(�	������ԾR*���a��|R@�$]����w�8�+���<z��=���=28�=�e�=�>v�>�/>֤>�i�=Ċ�=�G�=�2�=�׳=g��=��=�XN=h�=X��<�<�옻����|߼V��:�N!��x��L ���ϼ8m��(���TuǼ�z��cy��Ľ%���O��l�������fվ�g��yX	�{4��   �   �S�O!����PM�+���������M��]����h�m�$�<|~=�J�=��=G�=cv>5	>B
>��>�p>4��=��=E�=���=�=�-�=��n=�S3=�]�<�&W<����������ʟ/��6���-�@C���� ��׼����9��3��ϯڽRB �-�_��v��9��F���.�����   �   k{q�`�l��{_�I�J��0�$u�|��BQ��8|p��������B���=��=��=L�=n��=~>y1>"w>�  >"��=�X�=���=Xf�=nB�=��=F�=��h=��D=�-"=(p=Ln�< Ġ<�^�<�a<��X< �^<(�`<h%C< I�;	ƻ4���w�Egݽj@0�⸁�/���L��ϒ��0�4�J�:�_���l��   �   �m�\�h��j[���F�T�,�����T�z���.k���n�����'�x�=���=���=p0�=�B�=�G>��>br>H_�=n��=���={��=l��=��=���=��}=�]Y=ޝ6==�S�<��<�\�<(�y<��`<h-`<��l< �s<��Z<p( <���h�̼Nl��սhp+�dA}�,���^��g��:M-���F�f[�{�h��   �   |_`�J\�3�O��<��R#����V"־�e��$�[����H{����=��=s�=�Z�=X/�=�5�=Pq�=F��=���=n��=���=�}�=+��=ϋ=`p=�PK=��)="V=�m�<P��<(Q�< Or<��Z<�E\<ؼr<TE�<��<�ǎ<�PO<@Y�:�>����I�6'��0u��Lk� E����ؾ�6�I|#�M�;��nO��[��   �   "}L���H��*=�9+�#����ǰ��=l��Y�C�8�� �L����:$m+=���=��=��=r@�=��=��=���=0t�=��=�ӧ=�z�=0}n=T�@=�T=���<���<�~<�=;<��<p��;�� <H�<x(I<`$�<<�<0��<���<�[�<p�*<���������l��DKO�.����¾)���-�c�*�K�<�bH��   �   E?3�p�/���%�J������q־����v�
�%�$5�����X�&<�w==��=�{�=��=���=4�=��=&=�=Z_�=j=�=+m=�h0=��<x��<�g�;@ ^��ХG��RR���9�7���Z� -&;HJ<쀅<�C�<���<$��<�X�<Ȋ�<@��;�����e��׽=�+��3x�1����Ծ�� �����%�/��   �   &����ڃ���o�پ�0��؈����J��%�v	���N��p-�<WN=�n�=�U�=�K�=��=Ê�=s�=+۞=J	=N�6=���<�^�;pC5�<oټxt�0�?��P� bO�خ?���#��=��餼�U� �M;��n<8�<(0=�`=�R =�=p��< ����}�������E���B����վ����~Y
�#t��   �   ��򾶣�_����ʾ�Ȯ��2��R*]�� ���Ƚ��F��;޻XX�<��Z='�=z��=���=�
�=fX�=��=��Z=X`=��<��z��*#���������ý�ԽNxؽ��Ͻz���寠��}�Bs3��μ�h� !<���<r=�^9=�#H=��>=�=���<��ϻ��,��.������O��l��3Ȩ���ž�pݾ����   �   ���?���������k˅���Y��p&��轠������c�;��= `=�.�=��=�=�*�=���=�?=���<�<�D���b��Atǽ
l����-+�X�3��p3�_P*����!9�lҽQ���0E������5�:��<bI=�O=ܚk=\�o=DhX=t�"=�%�<��'��\A�Zݺ����yE��z�`Ӕ�����մ��   �   �x��m����:{��`b�y�A������,���@/��R<��|<��=(L\=V�=�Z�=T�=�n=�.=ҡ<�� J6�����' �S�)���O�V�n�ˁ��{��^ ���?{��eb���A�R��y��0��@F/��`<�h|<,�=�L\=&�=�[�=�U�=��n=�.=L�<���.>6�ꄫ��# �u�)�>�O���n��ǁ��   �   ?�3��k3��K*����5��ҽ�L��X*E�\��� ��:��<0I=�O=ʘk=n�o=^dX=^�"=��<((�gA��㺽���~E�(z�m֔���aٴ�v��$C���ì�۷���ͅ���Y�t&���������"輀O�;��=:`=n/�=��=q��=�,�=!��=��?=H��<�u;�����[���kǽpg����(+��   �   �Խtpؽz�Ͻ�������X�}��l3���μ�Q軈!<T��<�=X]9=!H=��>=��=H��<��ϻR�,�F4��T��-$O�\o��˨��ƾctݾ���z��I�����ʾwˮ��4���-]�*#�D�Ƚ��F�PT޻,U�<��Z=c'�=>��=2÷=@�=�Z�=ެ�=¾Z=�h=�<�Qz� #� ��� ��@�ý�   �   ��?���O� WO�4�?��#�81���ߤ��I�@�M;��n<L7�<�.=�^=P =�=,�< H���A���X�� �E������D����վ����B[
��u��������	���پ�2������<�J��'����U���)�<VVN=�n�=NV�=�L�=B��=���=^u�=�ݞ="=~�6=���<0��;p5�hVټ�g��   �   �k]�����G�07R�(�9��%� tZ�@K&;hM<���<,B�<���<X��<�S�<̄�<�y�;�ꝼ� e��׽��+�7x�3��Q�Ծ� ���8%�ŀ/��@3��/�z�%��������s־n	����v���%��7�������&<�v==��=H|�=���=���=x5�=h�=V?�=b�=�@�=H2m=�p0=���<�<���;�   �   P��<��<X,~<P;<H�<0��;�� <�<0)I<�#�<d�<���<���<�W�<@�*<�*�����I����wMO�������¾2���.���*���<��cH��~L�b�H�,=��:+�%��������Cm��حC�D�齶�L� {�:^l+=���=��="�=,A�=��=^��=r��=v�=��=b֧=j}�=^�n=ʫ@=t[=�   �   fTK=D�)=:Y=�r�<@��<�S�<XRr<��Z<HE\<Ⱥr<�C�<���<(Ŏ<�JO<��:$C����I�')��tv�yNk�F���ؾ�7�&}#�B�;��oO�!�[��``�I\��O��<�QS#�=��C#־�f��+�[�s��{�����n�=��=:s�=([�=�/�=6�=r�=L��=0��=֔�=<��=Y�=��=ы=Zp=�   �   V�}=f_Y= �6=�=�T�<|�<�\�<��y<��`<�+`<0�l< �s<`�Z<�% < ����̼�l�3�սq+�ZB}�Ƥ����թ��M-�[�F��f[�	�h�Tm�ݖh�,k[�Q�F���,�ͪ�U�Ƽ���k�+	����� �'�^�=���=���=�0�=C�=
H>�>�r>�_�=��=���=N��=H��=d�={��=�   �   �=��h=
�D=�,"=�o=m�<� <^�<�a<8�X<�^<��`<�%C<�J�; ƻ ���w�dgݽ�@0�����K���j�����"�0�A�J�B�_���l�g{q�V�l��{_�6�J��0�u�R��Q���{p�������h�B��=��=��=V�=l��=~>t1>w>�  >��=�X�=n��=0f�=AB�=��=�   �   �}=`Y=ڟ6=�=HW�<T�<$`�<��y<�`<�3`<0�l<0�s<��Z<P. <���`�̼�
l�9�ս�o+��@}�ǣ��������L-�e�F��e[��h�8m�ɕh�#j[�`�F���,����S�һ��k������x'��=B��=G��=�0�=DC�=!H>�>�r>�_�=&��=���=h��=k��=��=���=�   �   vUK=��)=�Z=�v�<���<LY�<h^r<�Z<PS\<��r<`K�<���<�̎<h[O<���:�8����I�i%��t�xKk�&D����ؾ46��{#�p�;��mO��[�j^`�8\�(�O��<��Q#�ޔ�� ־�d��Z�[�Q����z��г���=��=t�=�[�=80�=l6�=\r�=z��=^��= ��=h��=��=S��=Vы=.p=�   �   <��<0�<`5~< [;<h�<��;�<h�<�<I<�-�<�&�<\��<���<Xc�<p�*<����f����Ԙ�LIO�󋒾�¾R���,�)�*��<��`H��{L���H�I)=�(8+�����������j���C�^���L� I�:q+=Q��= �=��=�A�=\��=���=���=Xv�=0�=�֧=�}�=�n=��@=�\=�   �    Q]�X��P{G��)R���9����#Z� �&;�d<��<�N�<ġ�<���<�a�<��<��;֝�<e�%�׽ּ+��0x�F/����Ծq� ����
%�Y}/��=3���/�>�%������Eo־�����v�0�%��0��<����&<z|==��=�}�=ʎ�=X��=�5�=��=�?�=Jb�=�@�=�2m=~q0=��<��< ��;�   �   ��?�R�O�@TO���?���#�|'���Ԥ��1��dN;��n<0E�<6=f=�W =�=T�<  �����y����b�E��򇾛?��*�վy����W
�Hr�@������� ��]�پ�-������˶J��"�h���>���:�<�\N=;q�=�W�=�M�=
��=��=�u�=Xޞ=�=�6=0��<���;@5�@TټTf��   �   �ԽVoؽ�ϽN���a���p�}�"g3���μP�;!<��<�=�d9=)H=4�>=��=���<��ϻ��,�O)������O�ej��[Ũ�k�žYmݾ�������ྎ�ʾ�Ů��/���%]����Ƚ,�F�@�ݻ�f�<��Z=�)�=洬=`ķ=�=8[�=N��=��Z=�i=8<HOz�x#�8��7 ����ý�   �   ��3�.k3�*K*����4�~ҽ%J��z$E��w���U�:t!�<DP=#O=��k=��o=nX=��"=84�<�'��QA��ֺ��	�/uE�Kz�TД�w��hҴ�b��1<��X���б��wȅ���Y�dl&�I��8�����@��;�	=n`=�1�=i�=���=�-�=���=��?=���< l;�j��k[���kǽDg����~(+��   �   ox��5����9{�6`b���A�������q)��;/��:<��0|<,�=S\=��=�^�=�X�=��n=�.=��<��<26��}��j ���)���O�z�n��ā�Ru��,���64{�[b��A�������$���4/��)<�(:|<��=�R\=2�=o]�=�V�=�n=�.=��<����=6������# �W�)��O�P�n��ǁ��   �   ����?������ƴ��˅�	�Y��o&�������L����;p	=>`=%2�=i�=��=�/�=M��=(�?=���< �:�R��HT��zcǽ�b����K#+���3�f3�\F*�����0�?ҽ:E��.E��m��@��:$$�<DP=�!O=v�k=��o= jX=��"=�'�<�'��[A�ݺ����yE��z�RӔ�����մ��   �   ��򾖣�4����ʾ�Ȯ�S2��|)]���y�ȽH�F��޻Lb�<"�Z=�)�=���=�ŷ=��=j]�=��=l�Z=r=�?<�z��#�������ýv�ԽgؽH�ϽP���Y�����}�z_3���μp 軰B!<��<:=:c9=�&H=��>=��=��<@�ϻ�,�.������O��l��(Ȩ���ž�pݾ����   �    ����˃����9�پf0������ܹJ��$����8G���5�<V[N=7q�=`X�=�N�=d��=��=x�=-�=�=P�6=T��<0�;P�4��:ټ�X�^�?�Z�O�&HO�֖?�xy#����`ɤ��!���N;�o<�D�<�4=d=U =�=���< 0�.��}��{����E����A����վ����zY
�t��   �   B?3�m�/���%�<��s���q־�����v�n�%��3������&<{==��=�}�=j��=^��=b7�=��=�A�=�d�=D�=B:m=�y0=t��<��<@�;`�\�(���VG��	R��9����`�Y���&;�j<���<�M�<О�<\��<\\�<x��<���;�ߝ�e�ؕ׽(�+��3x�1����Ծ�� �����%�/��   �   !}L���H��*=�u9+����������l���C�;��ڜL� ��:�o+=��=@�=d�=|B�=Z��= ��=Z��=Sx�=���=T٧=���=��n=Ƴ@=�c=ܩ�<@�<�O~<Hr;<��<��;�<p�<@I<�-�<<%�<X��<���<�^�<0�*<`��\��}��Z��4KO�(��� �¾&���-�a�*�J�<�bH��   �   {_`�J\�2�O��<��R#����?"־�e���[�r���{�0᳻��=��=t�=\�=�0�=7�=8s�=���=���=���=6��=���=���=�Ӌ=!p=JZK=:�)=2_=�~�<���<�^�<�er<��Z<8U\<��r<�I�<X��<ʎ<@TO<@m�:�=��h�I�'��"u��Lk��D����ؾ�6�H|#�M�;��nO��[��   �   �m�\�h��j[���F�S�,�����T�m���k������ ~'�4�=	��=>��=�0�=xC�=JH>+�>�r>�`�=���=���=p��=���=��=���=x�}=�bY=B�6=$=[�<h�<db�<��y<`�`<83`<h�l<X�s<вZ< * <P���̼"l��ս`p+�_A}�+���\��h��:M-���F�f[�|�h��   �   >���'���(��-��v|��-T�{*��9��T��z�x�9[���}�� ���8=���=Ru�=^4�=R1�=tX�=f1�=���=���=���=�Ͻ=�۫=��=�ʋ=B�}=�h=�X=�L=.�D=��@=�@=h�C=,�G=�J=�F=�Z8=��=�,�<�P.��@#�ľ�n�)���������ǎ�,�R3U�}��7���-��$���   �   |M��&F��m��������w�[XP�9N'�<f���z��{-s�i�dNs���:�<=��=D��=t�=^`�=�r�=*�=��=�<�=�;�=s,�=�R�=9��=U@�=Ԩf=z=R=�0C=�X9=�P4=�3=&`6=��;=:�B=�{G=��F=p:=֌=��<�V�`�Yط�5%��f��!ͽ�D����(�1>Q�dwx������h���=���   �   �����䛿-y���G���k��3E�����P����b����~�T����;��E=��=��=��=���=d��=P��=*��=���=r-�=�ϖ=h+�=[=�9=�=�=z>=8r�<�j=�<
=P�=�$=V�2=�1?=��D=RO>=�q$=�"�<Ъ�;������������r�5���,Q��%+�^�E�n+k��8��i\��eϛ��   �   �`���Î�2����u�m�V���3�8����پ����.�I�����%���L<�S=��=>5�=���=+�=�}�=���=+ڵ=\`�=ŋ�=�H=�y=���<��}<�g< ��;0��;�"�;��,<4��< `�<hY�<G=�/=r�?=�=C=��2=��=�tP<P��H���O�.�U�*�d7ܾ�4���3�cV�(.u�Ć�����   �   Q���|�$6n�nwX�o�<��������%��>��`�)�B��2׼t�<2�c=��=��=�e�=L��=6n�=w��=x��=��I=,��<8U<@�s�Ғ�l�꼒H��r�&{�Џ��������*����:�c<���<�=��4=��E=��A=��!=d�<�E���8���νg�1�&��=���Ly��s���;���W�Jum�X�{��   �   ��Y��V�%J��g7������!Ҿ<�N{Y��U��0��@/� P�<Nr=Mɟ=���=�÷=��=���=��g=��=�HS<��=�J��l�����>����Ž�;ƽ�ں��r���n���]A� �伐��� <���<�v=d�B=�O=D�>=�=��=<�컼�X�����R�X�	X��˽Ͼ�R�h��6��I�^wU��   �   x�1�h.��$��	�\@�
�վG��6�w�б'�[�Ľ�8#��ț;�=�Y|=ce�=P��=l1�=Sj�=�}I=��<@`�@-	�Q����ʽ������p,�:p4�)3���(�TT��P���uĽu���`��%F�X':<���<��6=�V=�Y=��9=LM�< ��8�"�x׼�k	!�|yo�]u���RѾ�,���5�g?#�=�-��   �   f<
�j��j �x�a�Ǿ�e��	u�H�8�b��q���񌼄��<�P9=��=��=4j�=��|=N�7=���<��:�BH��p��_t	��M5���\���|�yK���鍾Z���LՃ���l�!�I��!�x�｝{���V&����@ח< �=��V=Non=D�c=� 4=P�<1�l S��tս<*���p����\���5��v���J���   �   l̾
$ɾ^���K���������n��6�ܼ���x��Ε��%;���<jM=�{=��=��n=x�1=���<��^��a��Խ"��V\����������;����ƾPp̾6(ɾG�������������n�2�6�8���[}��d����$;��<�M={=5��=`�n=̳1=@Ξ<��^�\{a��Խ6�!��P\�@�������~7��J�ƾ�   �   1捾����҃���l���I���!����Lv��O&����ݗ<��=��V=nn=��c=�4=h׸<pQ�(S��{սl@*��p�H���$���p��
�������>
����� �|���Ǿ�h���y���8�����t���������<LO9=��=��=�k�=\�|=��7=���<��:��H�ch��oo	�.H5�1�\���|��G���   �   fj4���2�V�(��O�hH���nĽ�o��TX�HF��7:<T��<��6=��V=B~Y=��9=XD�< ��8��"�#ݼ�!�/~o�Ex���UѾ�0���7��A#�Ƶ-��1��j.�j�$��4B�%�վ����w���'�{�Ľ>>#�p��;t�=LY|=�e�=���=V3�=�l�=��I=�+�<`���	�6퇽�
ʽ���|�k,��   �   ��Ľ>3ƽ�Һ�pk��Gh��*SA�ht�Pv�@� <���<Rx=��B=�O=N�>=�=��=<P���5]��b���X�fZ����Ͼ~T�l��6�f I��yU�G�Y�X
V�l'J��i7���4���#Ҿ2���;~Y��W�S3��p/�HL�<�
r=�ɟ=� �=jŷ=�=n��=��g=��=�sS<h�=��;�l�ڳ��F����   �   2;��e�2o�@z��8����*�@��: �c<��<�=v�4=��E=��A=��!=h�<h��8���ν�1��'��v���|�����;��W��wm���{�DR���
|�F8n�[yX� �<����>���'�����L�)��D���8׼���<��c=��=���=�f�=���=dp�=D��=���=ΤI=���<H7U<��r�,�������   �   ،<P�;P͟;�]�;(-<���<Dh�<T_�<I=� /=��?=J=C=��2=�=jP<�%��K��`Q�x�U���O9ܾ�5��3��dV��/u�qņ�y����a���Ď����u�бV���3�,��l�پ�����I�/�ླྀ�%�H�L<v�S=��=�5�=V��=8,�=D�=���=�ܵ=Vc�=<��=��H=H�=��<�#~<�   �   � =��=�C=8{�<ln=�?
=��=Z$=h�2=f2?=��D=�N>=�p$=$ �<`��;L���齣���^�r�[����R��,�h�E��,k�`9��]��Л���囿�y��9H���k��4E�6���xQ����b�r��J�T��{�;J�E=��=O��=p�=R��=^��=���=���=���=�/�=1Җ=.�=�[=��9=�   �   p�f=�?R= 3C=�Z9= R4=P�3=a6=|�;=��B=�{G=��F=,:=P�=L�< NV���pٷ��5%�g���ͽ����_�(��>Q�xx�񨍿/i���=���M��~F��im��ߕ��6 x��XP��N'��f��{���-s�_i��Ns��y:�<=&��=p��=Xt�=�`�=�r�=�*�=���=�=�=�<�=�-�=T�=���=�A�=�   �   �}=��h=X=hL=��D=��@=��@=�C=�G=bJ=��F=�Z8=��=�,�<�R.��@#�Kľ���)�э������ݎ�,�k3U�6}��7���-��$��>���'���(�� ���u|��-T��z*��9��T��'�x��Z�"�}� ���8=ӈ�=bu�=h4�=Z1�=vX�=^1�=���=���=���=�Ͻ=~۫=��=qʋ=�   �   ʫf=^@R=�3C=h[9=�R4=@�3=b6=��;=̋B=�|G=`�F=�:=�=�<��U�&��׷��4%�?f���̽�����(��=Q��vx�L���|h��5=��M���E���l��<����w��WP��M'�[e��z��a,s�Fh��Ks� �:r<=���=���=�t�=�`�=&s�=�*�=���=�=�==�=�-�=,T�=���=�A�=�   �   n =n�=�D=�}�<�o=tA
=��=�$=��2=�4?=��D=�Q>=�s$=p'�< ��;T���e������Jr�V���P��n*��E�h*k�%8���[���Λ�&���䛿|x��G���k��2E������O���b�T��6�T�@��;P�E=��=��=��=���=���=���=���=���=�/�=UҖ=9.�=[=b�9=�   �   ��<@��;�؟;�k�;�-<���<�m�<|e�<JL=*$/=��?=dAC=f�2=&�=��P<t��F��,N�4�U����5ܾ�3�_�3��aV��,u��Æ������_����?����u�ЮV�J�3�����پW�����I�O��.�%��M<��S=[�=�6�=��=�,�=��="��=�ܵ=�c�=h��=�H=��=��<�&~<�   �   @:�|d��m� v��@���H�*� ��:��c<���<�#=��4=��E=�A=�!=@�<`���8��ν�1��$��@����v������;���W�!sm��{��O��b|��3n�RuX���<�k��!���|#��j����)��=��d$׼H�<��c=��=��=�g�=���=�p�=���=.��=:�I=D��<�8U< �r����<���   �   b�Ľ�2ƽ�Ѻ�Qj���f��
PA�<m伈f�x� <���<L}=
�B=�O="�>=�=H�=<h߻��T������X��U���ϾQ�~��6��I��tU�-�Y�WV��"J�Ee7� ��޸�Ҿ�awY��R��+����.�T\�<|r=�˟=
�=[Ʒ=��=ⷕ=v�g=L�=�uS<ؕ=�;�R�l�����┶��   �   &j4�0�2��(�O�G��mĽ�m��`T���E�`J:<t��<�6=��V=N�Y=N�9=HY�< ��8h�"��Ѽ��!�uo��r��2OѾ�(��e3�=#���-��1�e.���$���K>�q�վ?��<�w�Э'��Ľ�.#���;��=&_|=�g�=�=H4�=�m�=��I=8-�< ��	�퇽t
ʽ����{��j,��   �   捾�����у�(�l�Z�I�ՠ!����bt���J&��s���<��=��V=�tn=��c=�&4=T�< ���R�nս�7*�k�p�哝���������������9
���� ��s�u�Ǿ�b��Do���8�����j���݌����<FW9=�	�=��=m�=<�|=��7=H��<��:�"H�/h��Zo	�H5��\���|��G���   �   �k̾�#ɾ8������\�����n�N�6�!����v������g%;|��<�M=p�{=���=R�n=��1=Dޞ<0�^��na�^�Խ}�!�2K\�����}��m3����ƾ�g̾�ɾ*~��_������V�n��~6����pq���� �%;<��<M=
�{=	��=��n=��1=�О<��^��za�޻Խ"�!��P\�:�������s7��<�ƾ�   �   `<
�`��\ ��w�*�Ǿ�e��gt���8����Ro���錼D��<|U9=�	�=K�=�n�=��|=�7=H��<�r:�H�.`���j	��B5���\���|�4D��j⍾���h΃��l�ފI�2�!�N�ｂn��"B&�h[���< �=�V=�sn=��c=�"4=\�<�,���R��tս�;*���p�����X���0��p���F���   �   v�1�	h.�
�$��	�G@���վ����w�$�'�פĽV5#���;\�=v^|=`h�=��=6�=.p�=N�I=�>�< �
��	� 函Qʽ���fv�e,�4d4�Z�2�e�(��I�3>���eĽ�g���J��E�p]:<<��<H�6=��V=؃Y=��9=Q�< ��80�"�+׼�P	!�dyo�Uu��zRѾ�,���5�f?#�<�-��   �   ��Y��V�%J��g7�������� Ҿ��zY�U�)/�� /�W�<`r=�˟=��=�Ƿ=�
�=���=��g=�=��S<�c=��,�*ql�֪������"�Ľ~)ƽ[ɺ��b��`��pDA��Z估I�8� <���<.=��B=O=j�>=
=Щ=<�껼�X��n��=�X��W��ŽϾ�R�f��6��I�_wU��   �   Q���|�$6n�iwX�f�<��������%�����)��@��p-׼��<`�c=��=���=�h�=��=�r�=Q��=���=n�I=���<�dU< r������f�L,��V��`��^���z���p*����:��c<|��<B&= �4=��E=:�A=J�!=��<=��$�8�h�νR�1�&��6���Jy��s���;���W�Mum�Z�{��   �   �`���Î�3����u�i�V���3�.����پ����ڇI�K��<�%�xM<l�S=?�=7�=ĝ�=�-�=(��=(��=Zߵ=�f�=䒀=
�H=t�=���<�M~<(�<�H�;�!�;@��;�3-<̲�<�w�<�l�<�N=�%/="�?=&AC=|�2=��=(yP<���@H���O��U�"�^7ܾ�4���3�cV�*.u��Ć������   �   �����䛿.y���G���k��3E�����P����b����Z�T���;2�E=��=.��=Z�=d��=���=��=���=���=2�=�Ԗ=1�=2 [=��9=� =��=�J=���<�t=zE
=��=�$=l�2=�5?=��D=�Q>=(s$=�$�<���;����ܻ�������r�2���*Q��#+�\�E�m+k��8��j\��fϛ��   �   }M��'F��m��������w�YXP�6N'�5f���z��d-s�i��Ms���:�<=���=���=�t�=<a�=�s�=x+�=���=�>�=.>�=�.�=�U�=2=kC�=�f=�CR=�6C=J^9=|U4=f�3=�c6=��;=��B=z}G=��F=�:=��=��<��U�&�Bط��4%��f��ͽ�D����(�1>Q�dwx������h���=���   �   �]�[�N�Կ�y¿�\��Q:���l��7�����e���ri�5'���>/�0?�<��k=���= H�=ʹ�=,��=(��=x��=4��=��=x��=�ێ=��|=jnb=��O=�E=�yC=�sH=2fS=$�b=T#t=�ɂ=�҉=,��=j�=�=w=�P>=,=�<P�f������uyz�"A���Q	�[=9��m��ܑ��ë���¿^�ԿfV��   �   3��G�ܿ&ѿ�;���y��c�����g���3��������2d������%�h��<�m=(�=�U�=i�=�=r��=���=���=���=sd�=@I�=��_=*7D=�1=�'=:P'=��.=B�<=O=<d=H�x=�/�=4߉=���=��v=PM@=���< �F�n���^��wt�� ��y��K�5��hi�
I���˨� Y��`!ѿb�ܿ�   �   Bwտw�ѿ��ƿs˵����+v����[��)�����l���HT�њ޽���]�<��r=�"�=nU�=�L�=µ�=N��=:^�=,�=���=��_=��/=j�=l*�<�&�<�O�<D¡<���<���<8?=��2=�^R=��m=�A�=sm�=. t=ܘE=4��<�׻�g�n��c��)��_;����+���\��ʇ�r+�� ���'�ƿm�ѿ�   �   V&Ŀ ���(���S����ؒ�6x���H�Ք��G������;�脽��
ü���<��x=4C�=$��=���=0*�=��=��=�e=z.!=dV�< 4�;�����e���������D��8)� \� �,<d��<�	=>�;=*^^=�:q=F�m=�8L=�L=@��:\�2�Ktݽ*�G�����l�	��h!I�!x�P���秦�Lj��7����   �   �����!$��8����ꁿ
�Z�N0�� �jþ���<���⓽��7���=|Q~=5s�=r��=2v�=���=�|=~/=���< H���¼N�4�z�x�M��(=������ᒽtQw���8��޼�e�P�+<��<np*=d�Q=V%a=�FQ=�P= �K<X.߼$����%��򅾢ž_f��0�:?Z�,q���q�������Ϫ��   �   ���9j��֣���|��>]���9�����c�bۡ�X�T����?K�`/#;֑ =�=��=c|�=[�=�W=0�<�y�;�ϼ"h�������$��c��|�#�\�!�<�����Cٽ���R7P������%;@X�<&�#=�K=��Q=��0=���<����{k�����?�V�?����J����)b8�,�[�u3{�������   �   f(u�J�p�+�c��<O�v�4����a�,���~�x,"�����ڼ,܂<��7=h,{=���=�bz=��==�>�<������5�bͮ�,Y��b.��0U��wt�����#	��1膾%8}��b�z�>�z����ڽ�ۉ�ԛ�� �F� B�<��(=�J=�C=�= }<D��[��7��dLz�"��������2�nM�̀b�"-p��   �   oJA�X�=�Ql3��"�sb�~�������>��j�;����jR�� �����<�H=2�m=��e=��0=���<ȱV���a�3�ֽ��#�i�^�Mi���}���k��DAɾ��ξ67˾�D�����uj��.+o���5����S��:��`�};�%�<b`8=BN=0�6=��< �@��e>��ԽO3��c��Lس��v徿�
�o� �b�1�!=��   �   �K����U���j��PҾ�����{��~�B�f����Ŋ�`���Pb<�K=�CP=�6W=��/=D��<�7��=d����
�4���j���n̾����=���N�a������o�#UҾv���~���B�;����ʊ�����a<�I=�CP=9W=��/= ��<h�7�d1d������4�j�@f��yj̾������c���   �   �ξr2˾@��n���f��(%o�ً5�k���WM���)����};<,�<�a8=dAN=��6=|��<@VA��o>���Խ�S3��f���۳�{�C�
�>� �k�1�.$=��MA�y�=�Eo3���"��d�}�����A��>�;�t�!R��F�����<lH=��m=�e=<�0=<��<��V���a�M�ֽ�#���^�e��Iy��g��p<ɾ�   �   1��X䆾�0}���a���>����áڽsՉ�4��� *@��J�< �(=J=�C=�=Xh<����`�����GQz�5%��|��p�m�2�qM� �b�v0p��+u���p�C�c��?O���4���e�����~�j/"�& ����ڼpւ<�7=@-{=9�=bgz=x>=�P�<�����5�gĮ��S�`\.��)U�Jpt�ڮ���   �   f�#�j�!�������:ٽP��+P�������;@b�<P�#=lK=��Q=0�0=��<���k�$�����V�����N����zd8���[�h6{�*	����������k��[���ٱ|�$A]�ī9�V���f�gݡ�H�T����hDK���";�� =j�=��='~�=��=�W=��<�֖;P�μl�g�W�`��[��X���   �   %4��͌���ؒ�tBw�z�8�|�޼0A���+<���<t*=��Q="&a=FQ="O=8�K<p8߼ӥ����%�u��ž�g��0�bAZ�ir��#s��o���IѪ�{������%��|����끿��Z��O0�"��kþ�����哽X�7�\�=�Q~=�s�=�°=.x�=k��=� |=�/=T�< ����¼Xx4�N�x�D���   �   �휼����-��h)��5Z��,<���<�=��;=�`^=�;q=��m=�7L=
K= G�:ʛ2�~wݽf�G������n�P���"I��"x�[�������k��z����'ĿY���L���]����ْ��x�$�H�֕�'I����t�;�ㆽ��ü���<l�x=�C�=��=b��=&,�=���=#�=p'e=n7!=�j�<���;�D��Ppe��   �   \6�<_�<|С<��<���<D=��2=�aR=$�m=lB�=�m�=F t=:�E=t��<�$׻j�g���Xc��*���<����+���\��ˇ�7,�������ƿW�ѿ,xտV�ѿ��ƿ,̵�F���v��l�[���)����}m���IT��޽B��\�<��r=:#�=V�=�M�=��=���=?`�=�.�=���=�_=�/=��=:�<�   �   ��1=��'=|S'=��.=֐<=4O=�d=��x=o0�=~߉=��=r�v=�L@=���<��F�z��@_��xt��!����ݹ5�8ii�mI��K̨�wY���!ѿޒܿ��࿻�ܿo&ѿ�;���y������U�g���3����C����d�C��d�%� ��<��m=`�=2V�=�i�=��=B��=���=膿=[��= f�=�J�=�_=�:D=�   �   ��O=��E=LyC=rsH=�eS=Οb=�"t=rɂ=�҉=��=�i�=�=w=�P>=�<�<�f�h���>���yz�QA��R	�|=9�@�m��ܑ��ë���¿f�ԿkV࿠]�[�B�Կ�y¿n\��>:��tl��7�ݍ��e��Hri��&��*>/�T@�<4�k=���=H�=ֹ�=4��=*��=|��=2��=��=r��=�ێ=n�|=4nb=�   �   �1=��'=�S'=�.=\�<=�O=�d=T y=�0�=�߉=���=��v=ZN@=���< �F���� ^�Jwt�� ��=����5�hi��H���˨��X��� ѿ�ܿ���ɝܿ�%ѿ(;��y�� ���E�g�"�3�S��B���d�4���%���<b�m=��=�V�=�i�=��=X��=���=���=h��=f�=�J�=6�_=�:D=�   �   $7�<`�<�ѡ<�
�<���<*E=��2= cR=��m=RC�=�n�=�t=�E=���< �ֻ"�g�� �fc��(��B:��݃+���\�Fʇ��*��b���T�ƿ��ѿXvտ��ѿ��ƿ�ʵ����}u��d�[�)�)������k���FT�$�޽��4d�<4�r= $�=�V�=�M�=P��=#��=f`�=�.�=���=,�_=.�/=&�=�:�<�   �   �으ț��0,�� 
)� �Y�@�,<�ú<�=�;=&c^=�>q=�m=�;L=P=� ;�2��qݽT�G�ͅ��=k���� I�}x�_���ڦ��"i������%Ŀ����𾶿.����ג�cx�R�H�����E�S����;�b���( üx��<y=�D�=���=���=�,�=蜬=1#�=�'e=�7!=k�< ��;�B���ne��   �   �3��n���Iؒ�.Aw��8���޼�8��,<���<w*=�Q="*a=�JQ=&U=��K<p#߼����҄%�-񅾠že�90�E=Z�
p��~p������LΪ�u������"������L避��Z�<L0�U��gþ���|��hޓ�@�7���= V~=lu�=�ð=�x�=ߜ�=J!|=V�/=��<������¼.x4��x��C���   �   B�#�<�!�e������9ٽM���(P����� �;�h�<�#=�K=��Q=��0=d��<��.tk�������V����H���`8���[��0{���z��r����h��A��� �|�<]�\�9�����`��ء�r�T����6K�@�#;�� =H�=î�=C�=��=�W=��<@ږ;��μ$�g�<�G��N��C���   �   !��B䆾�0}���a�M�>�"����ڽԉ�D��� �<�XR�<��(=~J=vC=�=��<���JV������Gz�4������;�2�,kM��}b��)p�%u���p���c��9O���4����]����ك~��("����H�ڼ4�<Z�7=P2{=��=�iz=�>=�R�< �����5�BĮ��S�T\.��)U�Bpt�Ю���   �   �ξb2˾@��I���f���$o�L�5�&����K��#��@$~;�4�<�f8=
HN=:�6=`��< a@�z[>�_�Խ�J3��`���Գ��r�W�
��� �i�1��=�8GA�(�=�Ai3�0�"��_���!����;����;�[�⽚R�֧��
�<��H=�n=V�e=h�0=��<@�V��a��ֽ	�#���^�}e��Fy���f��i<ɾ�   �   �K����L���j��PҾ����s{����B�!����Ċ�����`b<nP=�IP=?W=D�/=���<n7�&%d������4�A	��b��'f̾А�,������H��������e�PLҾ����Sx����B���������@导�%b<�R=dJP=�=W=��/=��<@�7��0d���㽾�4�[�>f��yj̾������b���   �   oJA�V�=�Ml3���"�db�V�꾨����>����;����xR�P��t�<f�H=jn=2�e=V�0=���<h[V�
�a���ֽк#���^��a��u��nb���7ɾ�ξ�-˾a;�����b��Lo��5������E�������~;�<�<�h8=�GN=.�6=@��<`�@��d>���Խ O3��c��Gس��v徿�
�p� �c�1�!=��   �   i(u�K�p�(�c��<O�j�4���~a����{�~��+"������ڼ��<��7=�2{=��=�mz=�>=8c�<�>����5������N�QV.�'#U��ht�誄�&��U���0)}���a�?�>�����ڽ`͉��n�� T5�X\�<`�(=�J=�C=p�=��<h��[����NLz�"��������2�nM�πb�%-p��   �   ���;j��֣���|��>]���9�����c�4ۡ���T�����<K�@_#;�� =�=x��=΀�=�=��W=�1�<@3�;T�μ��g��粽��뽊��.���#�$�!����I��c0ٽH���rP�p����H;ht�<ڵ#=�K=X�Q=��0=��<����zk�Z���$�V�8����J����)b8�,�[�w3{�������   �   �����!$��9����ꁿ�Z�N0�� ��iþv��ۻ��ᓽ`�7���=zU~=�u�=�İ=�z�=q��=(|=�/=�)�<�!��<p¼Dh4�Оx��:���*��]����ϒ�V1w��~8���޼��(&,<���<V{*=��Q=h+a=�JQ=�S=H�K<�+߼������%��򅾝ž]f��0�9?Z�.q���q�������Ϫ��   �   Y&Ŀ#���)���T����ؒ�2x�ٝH�ϔ��G������;�:����ü@��<hy=&E�=���=<��=`.�=]��=B&�=4/e=�@!=\�<���;�����;e��Ҝ�P������H�(� cW�p�,<�Ѻ<t=Z�;=f^=�@q=��m=�;L=�N=@��:x�2�tݽ�G�����l���g!I�!x�P���駦�Lj��:����   �   Dwտy�ѿ��ƿs˵����*v����[��)�����l��tHT�Z�޽���`�<r�r=.$�=W�=�N�=~��=���=ib�=1�=t��=��_=x�/=��=�J�<�G�<Xp�<X�<��<��<�J=��2=�fR=��m=DD�=jo�=t=�E=��<P׻p�g�X��c��)��];����+���\��ʇ�q+��"���'�ƿo�ѿ�   �   5��I�ܿ	&ѿ�;���y��c�����g���3����󏵾d����d�%����<еm=��=�V�=&j�=l�=��=���=,��=ϸ�=�g�=�L�=�_=?D=�1= (=�W'=��.=��<=�!O=�d=Hy=�1�=x��=���=��v=NN@=���<h�F�L��u^��wt�� ��y��J�5��hi�	I���˨�Y��a!ѿc�ܿ�   �   NM�����.	�(��޿|B��� ��6ms�c�5�H �)槾�mE��ʺ�0/���R=W��=VA�=|��=l��=���=�b�=��=�B�=���=�W=��4=xC=�=8�	=>8=�=$=��==t\=ڑ|=:�=C��=�_�=��=D�=
O9=8
T<��'�ܽIkT�G����,�2�8�Tv�wF��U,��7�޿�w���8	�����   �   ���RJ�������fڿ$��N����(o�Jo2��=��yX��z�@�������( =�1�=��=���=�=bK�=j�=�)�=�Ӊ=(�b=J�5=�(=�Q�<@��<�8�<W�<��=�5 =�B=�g=`��=���=��=L�=�	�=nD:=`�f<'���ս�O��Ǫ�̈ �b5��q�����dﺿ��ڿjC�����JB��   �   
�	��S�c �Y.��Ͽ����ې�p�b���(����h��T�2�����(�.���=&��=>6�=J��=Lо=Oj�=A�=�s~=x�A=�=�
�<(g < 0�7Pu������ H"����;��<���<hF%=�JT=4l{=�0�=.�=�~=z<=���<���9����?�5���c��,�*���d�H�������Aп��F ��<��   �   �P�����(k쿺�ؿ�Y������ӄ�W3O����־Qꉾ"��������R�Z"=BЇ=��=?�=�4�=:3�=�NS=P=�5N<�~�μ�K#�fnL�T�_���[��CB�e�@��������L<�M�<Z&5=��a=��w=��n=$>=�l�<�M���h��d�'�7�����پ��[SP�='��SȢ�����"ؿV��)����   �   sy�y�ݿ�ҿ�����#���Y����j��;6��'�G[���k�0�<�H���;�.,=�=0��=Fό=�5l=�A"=X��<��)����Ie��Z��5z�j4������C�
��Ͻ�-���G`�@w�@Dj�x��<�=��F=��U=.�;=`��<���3s��	�6�q�鹻�e���6���j������������ѿXݿ�   �   (����Ҿ�0������Gّ���v��G���������.=���ĽD�����w<8�2=�k=Υo=^7G=�'�< y;i �L@���޽Ξ�t@:���V�e�i�ܳq��vm�H�]��LD�dm#��=���®�0�G��8���z><��=Ĳ/=�Y2=�V=@�;���Ͻ`�@��֙�؆�k��F��"u��ꐿY���GA��xU���   �   4栿�B���������kp��NJ��"�?����!��� o�����ۅ���C��%�<�"2=�H=��*=���<p7�4�<��C��i����L������k��?9���J���^����������!2��櫇��3Z��C#�l�ܽ<�y�p]��l<D(�<�=�=�5�<����oC���R��m�<����O���
!��HH�a)n�ᇿ�'�������   �   n-��Z|��n�<BY�3�=�����?��HE���/��e.������ ا;���<��'=p�=���<h����T��ؽ~�-��v�>���=ƾ�羫/���	��C���
�x��HL쾳�˾�0���d���:���d�Pl��0BF<p��<��=$��<���;���4��2�)��,������Y���,]��Y;�S�V�A�l�j{��   �   %8C�_�?��R5��|$�����?�� ��6����>����nc]�H#��{�<Ƈ=��=̊�<����ĩC�RX׽�5������������+P�N1"�y�3���>��;C���?�V5��$�u��;D����:���]>�}罘l]�`##��u�<x�=�=l��<@h��f�C�|P׽~5�d���ԡ�����HM�."���3�H�>��   �   |@���
�����F��˾�,��pa��d:�K��ļ���\���TF<���<N�=p��<pБ;v�j:����)��/��y�������_��\;���V��l�n {�v/��S|���n��EY�=�=�����C���H��\2���h.�� �����0��;���<2�'=R�=轧<���H�T�H�ؽЂ-��v����8ƾ��羯,���	��   �   fY������؊���-������-Z�r>#��ܽ��y�(K��Ȅ<p/�<<�=�=�.�<Ԝ��,H���U���m�`����S��Q!��KH��,n��⇿�)���Ý�Q蠿�D����o����np��QJ�S�"�ɳ��J$���o�v��5߅�(�C��"�<F#2=�H=�*=���< �滶�<�<:������L�����Wg��i4���E���   �   �q�2om���]��ED��g#��3������@�G�<%��(�><|�=J�/=Z2=:U=@յ;���Ͻֳ@�^ٙ���m���F��%u��쐿4���CC���W��;����Ծ���H����ڑ�Z�v���G����������p1=���Ľ����`�w<r�2=�k=�o=�=G=$9�< 1	;|Z �Z7��9޽����9:�2�V���i��   �   �� >�E���ϽH%��9`��^�`�i�,ǚ<X�=X�F=L�U=&�;=���<���D9s�e�	���q�,��������6��j�p���9������[�ѿ�Yݿ\{�S�ݿ��ҿ����$���Z����j�1=6��(�
]��.k��1�6�H� ߼;�.,=��=���=�ь=J<l=\J"=�օ<�x)���\���O��)o��(���   �   4�_��[��4B�lW��������(�L<\[�<�+5=��a=��w=��n=� >=i�<�T���k��h�'�������پ ��TP�9(��|ɢ����C$ؿ�������&R�����l��ؿ�Z��	����Ԅ��4O�߆��־N뉾p��H��� �R�"=�Ї=�=��=[7�=f6�=dVS=�"=�bN<��$�μ.<#�j^L��   �   �$��@[�� ����;��<���<�K%=�NT=fo{=�1�=��=J ~=�~<=�}�<@%��;����?�P������(�*��d��������9п�뿟F �b=���	��T��c �C/���Ͽc���ܐ�Q�b�R�(������.�2�̮��H�.���=���= 7�=h��=�Ѿ=Tl�=�!�=z~=��A=2�=��<�� < 0�7�   �   ě�<B�<�_�<� =9 ="�B=�g=T��=b��=���=��=�	�=�C:=(�f<�(���ս�O�VȪ�@� ��5�єq�����ﺿv�ڿD�����B�$���J�������zfڿl$������C)o��o2�9>���X��Ś@�k������H =�1�=
�=���=��=`L�=��=,+�=�Չ=�b=��5=>-=4[�<�   �   ��=�	=�7=6=$=X�==�s\=��|=�9�=��=�_�=�=�C�=�N9=8T<h���ܽ�kT�z����,�X�8�v��F��k,��K�޿�w���8	����LM�����.	�(��޿cB��z ��ms�9�5�& ��姾vmE�\ʺ��-��rS=���=pA�=���=z��=���=
c�="��=�B�=���=�W=��4=PC=�   �   ���<LB�< `�<� =d9 =~�B=ng=���=���=���=  �=L
�=vE:=(�f<�%���սO�]Ǫ��� �5���q�k���ﺿ��ڿ�B��t�� B���� J�V������eڿ�#��‘�,(o��n2��<���W��v�@����� ���!=U2�=j�=ĵ�=�=zL�=��=7+�=�Չ=$�b=��5=N-=D[�<�   �    #�� Y�� ��P
�;�<���<�L%=�OT=�p{=�2�=�	�=t"~=<=���<��28���?�t���W��x�*���d��������nп�뿇E �<<�t�	�ZS��b �K-�+�Ͽ���Cې�<�b���(�K��H����2�Q���X�.���=���=�7�=���=*Ҿ=�l�=�!�=Dz~=��A=L�=��<�� < 0�7�   �   �_���[�P4B��V�h��������L<<^�<&-5=��a=N�w=��n=�>=�s�<�E��Zf����'�����پ�
�RP�e&��QǢ�h��{!ؿ��뿚����N������i�L�ؿnX��뻢��҄��1O�����־�艾���r���`[R��"=B҇=��=��=�7�=�6�=�VS=#=�cN<`��μ<#�L^L��   �   ���
>���Z�Ͻ�$���7`��[뼠�i�˚<��=*�F=��U=��;=���<���,s��	�n}q�������k�6���j�����@���v����ѿ,Vݿ�w῔�ݿ!�ҿ7����!��pX����j��96�7&��X��Jk�~-���H���;<4,=��=병=qҌ=B=l=�J"=(ׅ< x)�ʰ�\���O��"o��(���   �   �q�om���]��ED�Dg#�;3��幮�p�G�� ����><��=H�/=P_2=@\=�"�;X	�p�ϽD�@��ԙ���Ai�ŖF�8 u�_鐿����]?��sS������о�5�������ב�Ùv��G�����ྨ���+=�w�Ľ`���P�w<`�2=� k=��o=Z?G=8;�<@;	;Z �<7��*޽����9:�0�V���i��   �   aY������ˊ���-������6-Z�>#�/�ܽr�y�F����<�7�<��=�	=�B�<8����>��^O���m�d����K���!�FH�/&n�E߇��%��ɿ��䠿@��
������8hp��KJ���"�,���e����n���օ��|C�P4�<b)2="�H=��*=��<����<�:�������L�����Yg��k4���E���   �   }@���
�����F���˾h,��Ca���:�G�𽊻���V���dF<ȴ�<P�=���<�:�;���-���)��)��7��������Z��V;���V�}�l�r{�f+��U|��n��>Y���=�#���:��qA���,��X`.��������;��< (=>�=�§<X��X�T���ؽ��-�xv����8ƾ��羲,���	��   �   (8C�`�?��R5��|$����q?�� �����Z>���潰`]� �"���<8�=��=p��<P��ؒC��H׽�5�A���靵�ո羅J��*"���3���>�r4C���?�O5�Py$����{:����±��T>�]��>V]���"�Č�<`�=J�=���< V�� �C�P׽^5�\���ѡ�����KM�."���3�K�>��   �   p-��\|��n�6BY�*�=�����?��E���/���d.�x�����P��;T��<�(=\�=xΧ<���|T���ؽh}-��v����84ƾB���)���	�P=���
����\A���˾4(���]��p:�ɳ�J���XE��{F<���<��=���< �;���q3���)��,������X���-]��Y;�X�V�E�l�n{��   �   8栿�B���������kp��NJ��"����r!��? o�>��Yڅ���C�P/�<P)2=\�H=X�*=h��<`��|�<�N1��2��J�L�̳���b���/���@��8T����������?)�����n&Z�u8#�8�ܽ��y��1��Э<H@�<��=�	=�=�<P����B��TR�Чm�4���{O���
!��HH�e)n�ᇿ�'�������   �   +����Ҿ�1������Fّ���v�w�G�	��ɇ�����Y.=���Ľt���x�w<¦2=f"k=�o= EG=�K�< �	;@L ��.���޽����2:���V���i��q�;gm�R�]��>D�a#��(�� ���n�G�T��`�><�=��/=�`2=�[=��;|�t�Ͻ2�@��֙�҆�k��F��"u��ꐿ\���IA��{U���   �   wy�{�ݿ��ҿ�����#���Y����j��;6��'�*[��jk��/�
�H���;L3,=��=4��=�Ԍ=tCl=<S"=H�< D)�F��S���E��&d�8����68�����Ͻ���*(`��A뼠�h��ۚ<��=2�F=0�U=��;=���<`�໎1s�ޙ	��q�๻�c���6���j������������ѿXݿ�   �   �P�����,k쿻�ؿ�Y������ӄ�Q3O�ۅ�z־4ꉾ־�������R�~"=g҇=��= !�=�9�=�9�=>^S=Z,=��N< ���μ�,#�NL�t�_�x�[��$B�hH��i���I��8�L<@m�<35=��a=(�w=*�n=>=�q�<\J��Gh��<�'�,�����پ��[SP�<'��TȢ�����"ؿZ��-����   �   
�	��S�c �[.��Ͽ����ې�n�b���(����U�� �2�@�����.���=���=(8�=�¿=�Ӿ=pn�=U$�=(�~=��A=V�=�.�<�� < '8�ρ���� ���S�;�(�<< �<�R%=�TT=dt{=4�=�
�=r#~=��<=p��<��z9���?�.���_��+�*���d�H�������Aп��F ��<��   �   ���RJ�������fڿ$��N����(o�Jo2��=��oX��b�@�ݘ��0�� !=62�=��=2��=��=fM�=��=�,�=u׉=�b=��5=2=Le�<0��<�L�<�i�<�=�= =�B=|g=ؘ�=���=���=� �=�
�=�E:=��f<|&�`�ս}O��Ǫ�ʈ �c5��q�����cﺿ��ڿjC�����LB��   �   8�8��5��+�.��\_
��k���¿�I���2i�'�U��?�����"�Z��0<��R=ԍ�= �=�f�=�t�=Q��=͊�=�Rm=|p9=^1
=H`�<�2�<�q<��y<l%�<d��<��=�4<=�h=6È=��='.�=><�=0�{=D= �~�<�����N?��\h澍,*��|l����wĿ�����
����<�+�Z�5��   �   ³5��X2�B�(���#�J�迉���[���_e���#��۾r1�����ڃQ���-<&
R=2�=d��=3��=���=�J�=Ĵ=��L=RX=���<��\<Pg�;�*S;@E;��<��<��<�A=��M=8�{=^r�=K�=9�=P�w=Bc=�#0����č�j����ᾞ�&��*h��8��!�����P��lE��(��N2��   �   LQ,��?)� O �P�����ݿ�q��>���Y�q��9�ξ��|�D��7���V<2�N=�;�=ꖥ=tS�=P�=��s=��1= 6�<0�	<�@b�����bm�4���,�̼(q�@��`�h<�D�<�8=dk=��=�ن=��k=t�= B0:�xf��&�|����Ӿ�g��[��G���o��TB޿��&���& �D)��   �   ���h�Jn����￵3̿�է��)���PF��������a�Xo�,l�|�<G=�V�=a�=u8�=��J=Xf�<� <Ņ�L$��u{��㠽�h���;½y����)��̺��h|J�H� ����݊<P�=ҫH=�Pb=j�T=�= R�;J�9����T�i�՚��Z���H�kڄ�E���G̿��������(-��   �   r���H
��Y����Aտ�ᵿ�����i��F.�q��㠾�=>�a���T¼�,�<@9=�<`=XUS=<�=t��<PH�r�6�Y|����j��V�*��;�ҢA�F�=��/�.i����z���Eg��]ʼ �X;���<�`!=W1==Я0<����_Ƚr�D��������/� 
j��ꔿ�c���eԿ���V��l�	��   �   GH�Ov�⿗�ϿP���WC���~���F�h����̾d��� Z�~f��P2=�@s�<4$ =�$=d_�<P�;<E�����)�־Y��ł�xR��/㟾Z��3M�����@����:c���3���_h��$�&�P��\��<�(�<���<��{<����͓��n��u��T�;i��"F��}�vV��_����}ο�rΏ���   �   ��ɿ+�ƿ�ռ��򬿙|���!��LgQ���!�d�>���SL��߽��1� �|��<DO�<LǦ< 3U��O#��]��<k���W�G��������2Ͼ�羪�������NG����꾯UӾ�����蓾^�b�X �Y�Ƚv�H��0>��T<�@�<( �< I��~�=�Kw⽂�L����H��r� �'�O���P��E���5���Fƿ�   �   #+������c���M��p�r�φL���$�����ɬ����s���������r��(<�@�<���< Y��D�+�o_��)%�\v�mh��;׾ ��\��U-(��2���6��3���)�'�����ݾ7���$���-�MнFfE�p�#�:J<@�<@7�;�봼˯������=p�R:��l���`"���I��p��ꈿ�H�������   �   h�y��wu�kh�\�S���8�U}�����N�.�(�l3��M� %0�оz<B�< �o�~N��Դ���#�#�
{��L�J��?6�KQ�jyf��kt��y�6|u�>oh�<�S��8�B���#������3���f�(�B9��hT��b0��z<�F�<�-n�(E��ʹ��#����v���F�1���6�P
Q�uf�gt��   �   ��6�/�3�@�)�������ݾ������-�-��Eнd\E��#�XEJ<�?�<`�;0���������Cp��=���p���c"�(�I��
p�툿�J�������-������-f���O��1�r�	�L�<�$�������\�s�������|��X<�C�<��<0����+�>W���#%�Uv�d����׾������)(�9�2��   �   ����A����@PӾ�����䓾�{b���T�Ƚ��H��>��,T<�D�<,��<`h��ا=�}⽸�L��"��2��� �7�O����a�����������ƿg�ɿ��ƿ�׼�����~���#��jQ��!��
����xVL�O߽��1� ���̮�< V�< Ԧ< �T�jB#��T���e���W����ʙ���,Ͼ֡�V����   �   'U��VH��U
������3c�f�3�ؽ�+`����&��l㻠��<�/�<|��<��{<X����Г��q�x��L�;b�Q%F�$�}�AX��i����ο'u�@���J��x��⿸�Ͽ3����D����~��F���m�̾���`\�.i�� <=�ts�<�& =�$=ln�<9�;8)������h)�*�Y�@����M��Hޟ��   �   ��A� �=�V�/� c�5����p���6g��Dʼ�,Y;\��<e!=pY1=R=8�0<@��FcȽI�D�$�������/�Vj��딿9e���gԿ���v����	�����I
��Z����4Cտ�⵿�����i�1H.�Vs���䠾@>�䥹�4¼D,�<�9=~@`=[S=D�=���<��G���6��r��*���x�*��;��   �   �1½����@ ��;���FmJ�0ἐ>���<��=��H=�Sb=� U=ڡ=B�;X�9����ѡi��������1H�kۄ�JF��[I̿+�����,.����i�2o�j���4̿�֧��*��RF���������a�`q�@n���<<�G=X�=!c�=Y;�=~�J=�y�<02 <����|�#�Pd{�`ڠ��^���   �   �`�Ę���̼��p� ��h<<R�<p9=� k=��=�چ=h�k=��= �/:�{f��'�r�����Ӿ�h�E�[��H���p��cC޿���Ҕ�L' �)�R,��@)��O �������ݿTr������Y�
���ξ��|��D�>�7���V<��N=�<�=D��=OU�=}R�=Чs=�1=�G�<�
<����J��ܡ��   �    �S;��;8�<���<��<�E=��M=��{=Is�=��=y9�=r�w=�b=�70����������˭�1�&��+h�,9���!��?�鿦���E���(�*O2�,�5�0Y2���(�b��#����ն�������e���#���۾�1����$�Q�`�-<�
R=��= ��=#��=ꈯ=bL�=΂=��L=(]=|��<h�\<���;�   �   `�q<��y<�$�<���<��=�4<=��h=È=��= .�=<�=ʳ{=�=��~�s<��@���?���h澷,*�,}l�9���wĿ�����
����D�+�\�5�6�8��5�
�+�"��N_
��k���¿�I��Z2i��'��Tྭ?��l��>�Z�3<Z�R=���=< �=�f�=u�=f��=֊�=�Rm=�p9=X1
= `�<`2�<�   �   ��S;@�;��<���< �<�E=�M= �{=�s�=<�=�9�=��w=8d=`0���m��,������\�&��*h�{8��� ��?���� E�¸(�\N2�X�5�dX2�ܵ(���4#�������믗��e���#���۾�0��Ρ�*�Q�H.<R=�=a��=R��=���=iL�="΂=��L=*]=p��<`�\<���;�   �   �`�������̼x�p�@➺��h<pS�<*9=p!k=��=�ۆ=��k=�= �0:�uf��%�ց����Ӿ�f�1�[�AG��3o��{A޿�������% ��)��P,�?)�FN ����~���ݿ�p������Y������ξ��|��B�~�7���V<~�N=^=�=�=�U�=�R�= �s=
�1=�G�<
<���J��ܡ��   �   �1½����% ������lJ�� �8���<F�=D�H=Vb=�U=�=pq�;�~9����Z�i�v���f��RH��ل�D���F̿ ������,,����g�Vm���"�S2̿[ԧ��(��POF�޸�떺�4a�k�Hf�h�<��G=(Y�=�c�=�;�=��J=z�<�2 <����~�#�hd{�gڠ��^���   �   ��A��=�I�/��b�����Gp���5g�hBʼ�DY;0��<�g!=�\1=B#=`�0<���[Ƚ��D�b�������)/��j�E锿b��#dԿ���B��F�	�B���G
��X����?տ�ߵ�R��?�i��D.�Ln���࠾�:>�Ԟ��¼�8�<49=.C`=�\S=V�=ૃ<x�G���6��r��9�����*��;��   �   )U��UH��O
������j3c�4�3����_����&� [�H��<�7�<\��<h|<z���ȓ��k��s����;� �� F�V�}��T��z���p{οgp�C���E��s�*��Y�ϿJ����A���~�8�F�n����̾&����V��a�� =�t��<Z+ =�$=8r�<�A�; (�s���ץ�i)�1�Y�E����M��Nޟ��   �   ����A����3PӾ�����䓾s{b�����Ƚ��H�@>��<T<�O�<��<����=��q⽞�L���Ƕ�.� �V�O����_�����آ���ƿF�ɿ��ƿӼ��𬿇z�� ��9dQ�Q�!�r�>����NL�߽D�1� ���0��<�_�<ڦ< |T�TA#��T��pe���W����ϙ���,Ͼޡ�^����   �   ��6�0�3�?�)������ݾ����X��ʣ-��Dн�YE� �#��ZJ<�N�<�t�; ڴ��������8p��6���g���]"�{�I��p��舿9F�� ����(�������a��RK��t�r�U�L���$���������s�d��A���^��p;<�Q�<,��< ��Ĵ+��V��m#%��Tv�d����׾�������)(�>�2��   �   p�y��wu�
kh�[�S���8�K}����͙��"󂾻�(�52���I� �/���z<8V�<�l�v:�Ǵ��|#����r���A�F��B6�zQ��pf��bt��y�Hsu��fh�W�S��8�1z����������(��+���@� �/���z<�S�<�#m��B�7ʹ��#����v���F�5���6�W
Q�%uf�%gt��   �   &+������c���M��k�r�ǆL���$���������J�s�'��C���(j���0<�R�< ��<�̜�N�+�AO��^%�\Nv��_����׾�����&(�f�2���6�K�3���)�[�����8ݾ����\��k�-��<н|NE��#�`jJ<�P�<�c�;�䴼����R���=p�H:��l���`"���I��p��ꈿ�H�������   �   ��ɿ-�ƿ�ռ��򬿗|���!��DgQ���!�F�����RL��
߽�1� W�����<�d�<��< �S��4#�SL��`�ңW�풎�����'Ͼ���������:���꾙JӾ�{������\tb����wȽ��H���=��ST<XU�<8�<�#����=�hv�@�L����C��r� �(�O���S��H���:���Jƿ�   �   LH�Sv�⿘�ϿP���UC���~���F�\����̾8����Y�e��X!=���<�, =� $=��<���;�� �J��
)���Y����4I��jٟ�*P��eC����������+c���3����V��2{&� 
�l��<X@�<(��<�|<,����˓�Fn��u��J�;g��"F��}�yV��b����}ο�r�����   �   t���H
��Y����Aտ�ᵿ�����i��F.�q���⠾�=>�D����¼d6�<�9=F`=�aS=��=ȿ�<H�G��6�i��)������*�x	;�.�A�ڱ=�Z�/��\�}���pf��*%g��'ʼ@�Y;���<�l!=`1=x$=8�0<���^Ƚ3�D��������/��	j��ꔿ�c���eԿ���X��n�	��   �   ���h�Ln����￴3̿�է��)���PF��������a��n��i�T�<��G=Z�=�e�=f>�=�J=0��<�_ <䎅��#�S{��Р��T���'½�������0����\J�T�� ۙ���<��=��H=�Yb=�U=��=�j�;P�9�
��*�i�ʚ��Y���H�kڄ�E���G̿������ �*-��   �   NQ,��?)� O �P�����ݿ�q��=���Y�k��*�ξh�|��C�j�7�x�V<b�N=�=�=ܙ�=HW�=�T�=̭s=,�1=�X�<�<
<`��$3��̈�T�L����̼жp� ����i<\b�<D	9=@&k=] �=�܆=��k=p�= �0:Xwf�x&�n���y�Ӿ�g��[��G���o��UB޿��&���& �F)��   �   ³5��X2�D�(���#�J�迊���Z���^e���#�x�۾f1�����*�Q�H�-<�R=H�=ّ�=��=��=�M�=�ς=��L=�a=�<h]<��;��S;`�;P	<�<�<`J=�N=2�{=�t�=*�=�:�=l�w=�d= 0�J�����d����ᾝ�&��*h��8��!�����P��lE��(��N2��   �   |.d��x_�
-R�t�>�.@'��}�!S뿀e���ꎿ�0O�}}�r]����K�!츽��}���	=Q́=P��=�#�=,�=�΍=B�f=0�+=���<�1l<�Q�; qM��Tɻ�i����:�V<�
�<�r=^�D=�w=�
�=c��=U5�=�@]=Ԫ�<@�ȼ��˽�`U������}���R�i֐�pw���d�li�t�'���>��OR��z_��   �   v�_��+[�pJN�~4;�py$��4�v�翢U���z���wK�:�
�x�����F�f���6k��	=��}=�u�=ak�=}ϖ=��=��F=i=\l�< ;%;��X��䍢��f��PJ� ���,<к�<P�$=��\=Gۃ=�#�=
@�=~8X=(��<�ོ��Ž�BP��´����,�N��E���;��l�D ��%��x;��SN� [��   �   &S��O��CC�2�1�*{�����ܿ�e��`��͡@�?��O٤�0�8�������7�L�=PIl=@j�=�ԉ=�Jn=�0=���<�7�;𶃼���T4G�ةn���~�v�2U��U ��C��`�Z�0�<�=�eI=�mn=� r=>cH=�y�<H���2T��ņA�0e���g��WC��ц��ְ���ݿ������1� C���N��   �   �`@���<�(�2��1#��'��r���c˿�L��9bt�;�/�mH���M�#�u���P߻`��<��L=��^=� B=�� =xl<_����;�iӖ���ɽF�����T�	�������Խ����@Z�<�Ѽ �:��<��=�<=ʭ+=�ʽ<�=h��9����*�yŗ��#�)�1�-Pv�#����˿������`�"��:2�P�<��   �   �*�P2'����M��� �zܿ�7���%��ҰW�����ξf�}�����]�����<�3=�A=�o�<X] �T)��B���n���#���H���e�J"y�PD��0X{�jj�>iN��+����볽��J�D��8'<,�<���<$�<�U
��u�ʝ�6���s�о{!��X�/b��%���fۿ@ �h��*����&��   �   �l��T������>޿�ƽ�����|�t�Z�6��`�e
��V�N�,(׽t
 � v�:�<@�< �;p(����{�����)��"e�������M⾾ԟ̾A�Ѿ
�;�V��yE��������m��2�Í�K������ h��0�x<8�s<@�k�V2��&߽��Q��m�����J7��!t����`�����ܿ������R��   �   h��[
�DD俣}ѿwS����������<�H����k�Ͼ^چ��/��O���μ W*;��<@i̺x��L����o���M�J����~���bᾮ�ީ��9���I�"'�V�1��%������U�
��t������ �ѻ ��; m��v弘̠�S��K��qTϾ��}G�t��O��;�����ϿZ��c)��   �   ?�Ŀ����#��@������/�{���K�-�*{�5/��6�G���mK�h�_� m :`���@"���Y����\`�a��|�׾�G�Y $���<�.mP��=]�� b��>^�ER��&?�՞&�!�
�A9ܾ����f�.)��C�����E� g���It�"hM�a^߽��F�>М�`;�=��H�I�7�x��I榿k���w����   �   �������b��� ���d�S�?������꾀���F�a�4���&��L<ڼ ��P���D�м����|�"�]�����.羍����<��a������B��C��������!��be����d���?�� �4�����d�a����=+���Eڼ����p���мR��xx�[�]�����)�q����<�Ia�\���L@���~���   �   ;�a��9^��@R��"?�I�&��
�E4ܾ� ���f��$��=������7� h��HXt��oM��d߽��F��Ӝ��?�����I�P�x�c��覿3���\���,�Ŀf����������F����{���K�����2��/�G��"��rK���_��� :�n������R��$���`�"��2�׾�D���#�p�<��hP�+9]��   �   :��}��#��e��4�������U�*��_�������ѻP��;�[m����Р�Ȯ��!���WϾi���G��w��Q��������Ͽ@��j,�u��W�G�9�ѿ�U�����������H�Ƕ�m�Ͼv܆��2�(S���μ b*;� <@|˺���V���Bj��M�����y���\�S�;���5��   �   <�Ѿ&�;Q��`@��&�����m�D2�̃򽭇��|�� |�8�x<0�s< l�f2� +߽bR�yp������	7��$t��������ܿ���J��\T�������������@@޿|Ƚ������t�[�6�hb�z���N�s+׽v ��t�:��<��<�G�;���"�{�)��p�)��e������詾�ܾ��̾�   �   �?���O{�=	j��aN�` +��Z⳽��J�d��`8'<��<���<�<0^
��u� ��ꣁ��о.#�H�X��c������hۿ` �������(�&�V*��3'�f���N��� �4ܿf9���&����W�!���ξ��}�Z���]� ����<8=�H=���<p+ �R	)�
9���b��B�#���H�9�e��y��   �   �N����y��Y�Խ����0Z�8�Ѽ�{:�%�<Z=��<=��+=\ʽ<�Fh�F<����*��Ɨ�&񾢞1�Rv�E$���˿�������~�"��;2���<�.b@��<�P�2��2#��(�5t���d˿�M���ct�O�/��I�����#����� ߻���<��L=h_=�'B=�� =��<pC��4�;��ɖ��ɽ������   �   ��~�v�u�>qU�I � -��@OZ�l��<P=�jI=�qn=�r="dH=y�<@���V��V�A�Zf��mh��XC�B҆��װ��ݿ��J����1�C���N�*S��O��DC��1��{�2����ܿFf���`����@�����٤���8�d���0�7�.�=NKl=�k�=׉=�Pn=J�0=<��<Њ�;T���|��(&G��n��   �   ����X��0�I��o�p�,<���<�$=��\=h܃=Z$�=@�=�8X= ��<�㽼ȋŽ�CP�Gô����ܳN�IF��k<���l鿢 ��%�
y;�lTN�� [��_�,[��JN��4;��y$��4�Α��U��{��xK�k�
�����6�F��f��h6k��	=��}=�v�={l�=�Ж=ޤ�=��F=n=�w�<��%;�d�(���   �   �Uɻ�j�� �:�U<T
�<�r=�D=�w=^
�=4��=$5�=&@]=���<�ȼ{�˽�`U�󯸾�}��R��֐��w���d�|i���'���>��OR�{_�|.d��x_��,R�d�>� @'��}��R�ae��bꎿ�0O�U}�3]����K��븽��}�Z�	=�́=r��=�#�=7,�=�΍=n�f=T�+=0��<�1l<�Q�;�rM��   �   ����X�� �I� n���,<P��<^�$=��\=�܃=�$�=�@�=�9X=`��<�޽��ŽvBP�D´�ǥ�߲N��E���;���k� �6%�,x;�nSN��[��_��*[��IN�4;�y$�V4�ڐ� U��bz��+wK���
�������F��d��-k�	=��}=�v�=�l�=і=褀=��F=n=�w�<��%;e�D���   �   �~�z�u�>qU��H ��,�� JZ�`��<�=VkI=�rn=�r=XfH=p�<�����R����A�md��g��VC�ц�Sְ��ݿ������1�@C���N� S��O��BC�\�1�rz���ݝܿ�d��a_����@�k��ؤ�w�8� ���H�7�=&Ml=dl�=u׉=�Pn=|�0=d��<���;`������J&G��n��   �   �N����y��G�ԽW��p0Z��Ѽ �:�'�<�=ָ<=��+=4ӽ<p,h�X7���*�Oė�J"��1��Nv�"��y�˿������Z�"�f92��<��_@�|�<��2��0#��&�+q��'b˿�K��[`t�Ƞ/�EF���
�#����0�޻���<�L=_=�(B=*� =��<,C��>�;�ʖ�*�ɽ������   �   �?���O{�@	j��aN�J +���⳽��J�� ��p?'<(��<���<�(�<�>
��u��������k�о �2�X��`�����&eۿ8 �:�����>�&�\*��0'����PL��� ��ܿR6��X$����W���#ξ��}�(���]�������<>;=pJ=܄�< ) �	)�9���b��N�#��H�L�e��y��   �   E�Ѿ+�;Q��Z@�����݆m�2�L��������� ��(�x<��s< �k��2��!߽��Q��k��F��=7�St�`��r���w�ܿ���r��XQ��������N����;޿xĽ�+�����t��6�!_����n�N�["׽@ ��y�:\�<l$�<�X�; ����{���n�)��e�����詾�ܾ��̾�   �   ?�����#��Z��$�����m�U�Ը�e��� �� sѻ�ڷ; )k��e�zǠ������KQϾ��
{G��p��M��𘷿q�Ͽ���l&�\��V�]A��zѿQ������'���>�H�`��ӮϾ�׆�,��I����ͼ@�*;@% <�˺�����j�
�M�����y���\�Z�B���5��   �   C�a��9^��@R��"?�E�&��
�04ܾ� ��οf�^$�g<������ ��X���&t��]M��W߽��F�<͜�a7侩���I�d�x��풿�㦿��������X�Ŀ����[ �����������{�=�K�W|��v��+��&�G��:aK� �_� �":�D��@	���Q��ީ��`���4�׾�D���#�w�<��hP�29]��   �   �������b��� ���d�N�?����~��]�����a�����$���1ڼ ж��*��L�м��dt��]�1��+%羋��y�<�<a�����=���{��c���G��S`��V����d���?����}�꾂�(�a��������%ڼྲྀ�`6����м���	x� �]�����)�t����<�Qa�a���Q@���~���   �   D�Ŀ����&��@���
���)�{���K�"�	{�	/����G�*ཎhK�0�_� �":�$��x���|K��m���`�(���:�׾�A�.�#�|�<�rdP��4]���a�J5^�F<R�y?���&���
��.ܾY���I�f����5�������@2���/t�dM�#]߽��F�(М�Y;�=��K�I�=�x��M榿q���}����   �   m��_
�GD俤}ѿwS����������1�H����H�Ͼ*چ�X/�N��μ��*;@0 <�Gʺ���{���*e���M������t��W������1�`����������S�����m����U�����������:ѻP��; k��k��ʠ�֪�)��cTϾ��}G�t��O��>����Ͽ`��i)��   �   �n��T������>޿�ƽ�󽛿v�t�Q�6��`�<
��ևN��&׽� � Q�:��<�-�< ��;X����{�����)�e������㩾#׾��̾?�Ѿ5�;fK��;��o����~m�m2��x�~��$�� �ٸ��x<x�s<��k�2�@%߽x�Q��m�����K7��!t���c�����ܿ������R��   �   �*�R2'����M��� �zܿ�7���%��˰W�����ξ�}�B��>]� ��(��<~>=<P=$��<p�����(��/���W����#��H��e��y��;���F{�� j��YN�h�*� �س���J�肼hd'< ��<���<�+�<�A
�^u�L�����d�оz!��X�/b��&���fۿB �j��,����&��   �   �`@���<�*�2��1#��'��r���c˿�L��5bt�4�/�XH�}���#�;���0�޻P��<L�L=

_=�.B=p� =P�<�(��r�;�������ɽ�����uH���Mn����Խ����Z�X}Ѽ��:�9�<x
=p�<=r�+=4ս<x/h��8��p�*�cŗ��#�(�1�.Pv�#����˿������b�"��:2�R�<��   �   (S��O��CC�4�1�*{�����ܿ�e��`��ȡ@�9��<٤���8�̓��8�7�� =@Nl=�m�=\ى="Vn=<�0=��<ڃ;\������4G�@�n�ؠ~�t�u��bU�|; ������Y��<=qI=�vn=�r=.hH=��<����zS����A�#e���g��WC��ц��ְ���ݿ������1� C���N��   �   t�_��+[�pJN��4;�ny$��4�v�翡U���z���wK�7�
�n�����F�f��x2k��	=��}=yw�=�m�=CҖ=���=��F=�r=���<`&;�I����q��HJ�� �I�`��-<���<��$=��\=ރ=�%�=�A�=�:X=���<x޽�(�Ž�BP��´����-�N��E���;��l�D ��%��x;��SN� [��   �   
������~N|���b���D���&�1	��ۿL����u�z�)�M^۾� ���� ���!��X�<�mO=�ʊ= c�=�o�=�Qk=��/=���<�Z,<`���O��8J��`jؼ�Nɼ�x���;�@��;<�<��= U=��='��=��}=�h7=�/<B<�����W@�p�,��{y��6���kݿp
�Ĺ'���E�)c�j�|�H����   �    ������/w��P^�}A���#�� �̈́׿fM���q���&�G�־�Z|��H���t�T�<)I=��=p��=d_=�XM=�"=c�<@�����H����A���,��c$����,���`�����8<���<7=�jh=��=(^r=0s1=��.<� 6���n'��g�۾��)���t��E��\�ٿR�.�$�`7B�h�^��Aw�����   �   P�}� $x�@�h�bR���7�r���� ��CͿ�$��.e�����Sʾll� ���*���<
�5=f�e=��a=�p7=���<�D�;�爼�!�4{u��/��L/��g������v������3�t`�����:��<�� =�K=r�N=B�=�'<%������?s��xξ�
 ���g�������ο|k�>����7�NR��h�~�w��   �   �e��`��pS�2�?�ܔ(�F��	e����WI���]Q��D������R�p̽��Жd<�0=ư&=6w=8Qk< s8���*�Oɗ�!ٽ��	��*!�Â0��Y6��2�*$�j��"��w����XA��/���i<�t�<x�=0��<2<���}�׽��X�����$�1hS�CU�����2��X(�La?�t�R�P`��   �   �oH�(�D�:9:�P�)����L ���ӿML�����-/8����h͝�Z�3��?���'��X�!<�b�<`ۑ<��E�P��������P转3$�hFS��}�ݮ��K����垾���L|���9��U�X��J*�~���=w��
�ĻX�R<��<���;����h��`X8��@��Ҝ���d9��B��<�����ӿ`���dk�z)�L\9��YD��   �   &�*��!(����J�ȗ�ݻݿ���d��ĴY���cѾy���;�PN�� $�� �#;`"Z;H\a���=������7Z�i���ܕ����Ͼ�D����k��]Y���꾕Ӿ"���=���a����1`Ƚ^bR����� 4H��s��`���)����=���2gҾh���Y�*��Y���qܿ�� � >������'��   �   ����"��l����ؿO�������P'n���1�ߜ�����ЕK��ݽbI�`]����0����Ab��ٽ�11�f��:~���9�za����.��9�x�=�wc:�
0���~
�Qg�U���]����6��⽪pr��FԼ�yH����f?R�{3���L�� ��-M��W1�o�l�⣖��f��{�ֿ7V��.��i��   �   Ԧ�4+�׿A_ſJ���fW��|�q��<��
�Ź��E�{�j��ޡ�����-����ؼoe�3eܽ<<9�N�����žҵ���#��C���`�(w��킿 ����u��[y���b���F�3Q&�2��Yɾ�t����=�G���o��Y��ة��������Xg���z�Q���N�	��g:�pXo��Œ�M���l�ÿ�տPJ��   �   	��+>��R^��e&���̆�/�c���7����Qξ������1�FPʽ��L��NԼ�3Ҽ�I�dTǽD</������˾E��i�5�B�`�9��3���##��Z�����/A��2a��)���Ά�B�c�D�7����oξ�Ì�˝1��Uʽ$�L�0QԼ�-Ҽ��I�Nǽz7/�������˾Y��Ζ5���`��6��{���7 ��Q����   �   N���'s��Uy�J�b�o�F��M&�J��wTɾ[q����=�G�J�o�\Q��ة��������j��z�%�����	��j:�p\o�Ȓ�����c�ÿK�տ�M�0�忀.�5׿bſك���Y��.�q��<�T�
������{�l��;������)����ؼ�de�4]ܽ�69�{�����ž���9�#���C��`��"w�낿�   �   ��=�_:��0�?���z
��a�RP��.Z��F�6�ˑ�Zer��8Լ�nH�(����DR�z8���L����IQ���Y1���l�����Ci��H�ֿSY�0�hk���������o��#�ؿ��������b*n��1�c�������
�K�ڌݽ"eI��[��P��X����4b���ؽ�+1�h���>y���3��]�2����.�|�9��   �   i���}R����꾠�Ҿ����9��}�`����MWȽlUR�8r����F�@A��<���,�����L���5jҾ|���Y����l���|sܿ�� ��?�|��n�'��*�t#(����dL����ݿ㷶��e���Y�����Ѿ���=�P��H$����#;��Z;�3a���=�j����z�Q/Z�ű��v�����ϾJ>�����   �   ��������w��65����X�%D*������n�����нû��R<��<���;x�强k���Z8��B�������f9�@D��Ւ����ӿ�����l�)�^9��[D��qH���D��::���)����M �-�ӿ�M��Ɔ��08�7���Ν�%�3�uA���(���"<pl�<��< %C�����K��eE��,$�v>S�%�}����8����   �   �R6��2��#$�j�����X����IA������<��<�=���<�1<��0�׽Y�����B%��iS�\V��*�����NY(��b?��R�`��e���`�rS�n�?���(���]f���,J��'_Q��E�L����R��q̽T��h�d<4=*�&=�~=�yk<H?8�*�ֿ��1�ؽ��	�8$!��{0��   �   �������m��|��Ȣ3��I�� ȓ:���<H� =�K=�N=\�=ع'<F%����QAs�zξ� �4�g�������οl� ����7�dR��h���w���}�d%x�\�h�NR�\�7���n� �yDͿM%��e�U��|Tʾ_l����R+����<B�5=��e=z�a=w7=��<`��;�ψ�X�!��ku��'���&���   �   ��,��[$���4����x��09<|��<�
7=hmh=��=:_r=ts1=��.<�6�ڠ�(��D�۾W�)���t�GF����ٿ����$��7B�
�^��Bw����| �����d0w�Q^�z}A���#�$��׿�M��T�q��&���־�Z|�I���t���<P*I=��=���=�b=�\M=�'=�n�<@�d搼�w��~9��   �   �jؼ�Nɼy���=����;��<��=�U=D�=�=>�}=h7=H�/<6	<�T�����@ྟ�,�*|y��6���kݿ(p
�ع'���E�,)c�x�|�K���
������nN|���b���D���&�1	��ۿ*����u�K�)�^۾T ���� ���!�Z�<JnO=�ʊ=%c�=p�=*Rk=�/=���<p[,<����O��0J���   �   ��,��[$���(����x���9<���<�
7=�mh=��=`r=�t1=P�.<��5�ʟ�8'���۾��)�z�t��E��	�ٿ���$��6B��^�HAw�9�����/��/w�P^��|A�B�#�� �7�׿�L��=�q�L�&�i�־QY|�G��r�8��<p+I=��=�=�b=]M=�'=�n�<�ẜ搼�w���9��   �   ʯ�����m��t����3�TI���ғ:���<� =K=��N=��=��'<�%����G>s��wξ�	 �
�g�%���	�ο k����7�ZR��~h�6�w���}��"x��h�TR���7����`� ��BͿ�#���e�ʜ�SRʾpl���<&�|��<d�5=2�e=B�a=tw7=p�<���;�ψ�t�!�"lu��'���&���   �   �R6��2��#$�g��m��3���IA�X����<���<�=���<E<�����׽��X�w���#��fS�gT��������W(�`?���R��`� e�>�`�oS���?���(�P��oc���EH��;\Q��C�J����R� l̽T��d<�6=��&=�= |k<X>8���*�࿗�G�ؽ��	�F$!��{0��   �   ��������w��65����X�D*�b���1n�������û �R<4��<�گ;Ԉ�e���U8�O?��y���^c9��A��Ꮸ�#�ӿY���.j�)��Z9��WD�
nH�R�D��7:���)�F�tK ���ӿ�J��/��:-8���L˝�N�3�;������"<\s�<��< �B�T���+��jE��,$��>S�:�}����D����   �   v����R����꾟�Ҿ����	9��Z�`�����VȽ�SR��l����E��u�� ��U%��D~�]����dҾ�
���Y����~����nܿL� ��<���ʍ'�H�*��(�4��TI�d��s�ݿ���Zb���Y�ݕ�LѾ9���8�I������-$;��Z;�*a�8�=�����z�R/Z�ʱ��������ϾY>�����   �   �=�_:��0�?���z
��a�AP��Z����6��⽌br�t0Լ�TH��梼6R��-��L�I����I���T1�V�l������d��ݦֿBS�H-��g�H���r��i����ؿ�򸿚����#n���1�����	���I�K�N�ݽ�VI�HI����̕���2b�1�ؽv+1�`���@y���3�^�9����.���9��   �   R���*s��Yy�L�b�l�F��M&�B��`Tɾ8q���=���:�o�E�(Ʃ�Έ�Ɓ���c���z�ׂ����	��d:��To��Ò�ũ����ÿ�տG�{���'��׿E\ſ�~��U��x�q��<�w�
�ֵ��n�{���*���L������ؼ�`e�\ܽG69�k�����ž²�>�#���C��`��"w�낿�   �   	��/>��V^��g&���̆�+�c���7���2ξ�����1�sNʽ��L��=ԼDҼX�I��Fǽ�2/�c�`˾���s�5���`�W4������c��S������";��f[���#��ʆ�ݮc�?�7�	���ξ\���[�1�<Hʽ��L�\8ԼHҼ<�I�hLǽ7/�l�����˾Y��і5� �`��6������= ��W����   �   צ�9+�׿@_ſH���dW��v�q��<���
�������{����o���4������ؼ�We�Uܽ"19�梌���žܯ���#���C�Z}`��w�p肿����}p��4y���b�"�F��I&�*��mOɾgm��v�=�
���o��9�é�f��L����f�D�z�<���J�	��g:�vXo��Œ�R���q�ÿ"�տWJ��   �   ����$��l����ؿM�������I'n���1�����췦�,�K��ݽ�[I��J���������2'b���ؽ�%1������t���-ᾨZ�n����.�!�9���=��Z:��0�O��(w
�t[�;K��V����6���⽰Ur��ԼDH��墼~9R��1�r�L�� �� M��W1�r�l�䣖��f����ֿ=V��.��i��   �   (�*��!(����J�ȗ�ܻݿ���	d����Y���<Ѿ8��2;��K����@J$;�[;Ha�,�=�(뼽�t��'Z�X���G�����Ͼ�7���p����K���|꾀�Ҿg���[4����`�N��MȽTER��X���TD����� ��C'��J�����gҾf���Y�+��\���qܿ�� �>�Ĥ���'��   �   �oH�,�D�<9:�R�)����L ���ӿLL�����%/8����8͝�ġ3��=�� ���"<�z�<���< c@��w��|v���:�Q&$��6S���}�N���7����۞������r���0����X�*=*�����d��H���ZûS<x �<@�;t���f���W8��@��Ü���d9��B��?�����ӿe���hk�|)�P\9��YD��   �   �e��`��pS�2�?�ڔ(�F��e����UI���]Q��D�����6�R��n̽����d<T9=t�&=Ć=��k<�8��w*�ö����ؽ��	��!��t0��K6��2��$�:��^�⽧���9A�p�����<$��<H
=t��< J<|��6�׽f�X������#�1hS�EU�����5�� X(�Na?�v�R�R`��   �   R�}� $x�@�h�dR���7�r���� ��CͿ�$��*e�����Sʾ*l�)��D(����<��5=�e=��a=f}7=��<���;���6�!�8]u����4�� ����䴽�e�����ʔ3�L1��@�:d�<�� =�K=�N=��=p�'<r%����F?s��xξ�
 ���g�������ο|k�>����7�PR��h���w��   �    ������/w��P^� }A���#�� �τ׿gM�� �q���&�>�־sZ|�kH���s�@��<�+I=}�=嬋=�e=�`M=n,=ty�<�N�dؐ�0h��\1�F�,�nS$�
��Ds��B���9<���<�7=&qh=?	�=�ar=�u1=8�.<��5���b'��b�۾��)���t��E��\�ٿR�0�$�`7B�h�^��Aw�����   �   �H���c��,e���Q����a�`$=����y#��Z������RC��.���R��8L!���x��;x"=L�o=Cr�=>q=:\A= =�Y[<P(���奼����(�V�5�X,�����{��` �8)<l1�<�l3=�c=$ev=��`=�m=�������&�~������
F��Ӎ�jq��ٓ��5��h>�(�b�ˢ��օ��Ui���   �   p����Ԛ�o/��R���X�]���9�<`�C0�;��������?�.:��������¬r���:n.=T�b=|�q=4EW=�) =,v�< ;�: M���l���J�>�o��~��s��Q�T� x���NѺH�<�=��H=�,c=R�S=L�=@������#�Fm���Y��[B��Q��e-���k��֍��:��i^��׀�@<��CϚ��   �   �&���Ɛ��!���r��Q���0�n� �翘!��谂��m5���뾓ތ���00a� ��:��=Z�:=��6=�=�i<����"��^v�+y��Yνrm��t�P��ODҽ�ծ�������@�R�H�.<�7�<�C(=:r,=��< k5��r�6�cۏ�ւ�e�7����Q����_�x��V.1�V�Q���q�l���m����   �   �ʄ����z�s�v�[�s?��M"����D�տ�ʣ�`Po�;A%�r�վ�=}���VIH� �k��
�<�<��< Y!��~�
퀽�˽8�	���*�>�D��U� �[���V�f�F���-�A����ҽMf��𫌻��<x��< �<࢑�j�W��a�� ���ؾ��&�r?q��Ѥ���ֿZ.��g"�84?�z [���r�g����   �   �f���a�̟T��A�ک)�Ԧ���>o��
Z��&S�b���u��T�Y�^@߽��-� \��ؑ< �^;����6�O�,��������H�v�}�sw���a�����HA�������㪾�x��
��$oM��k�ΏȽW_��	�� ,�8�q�;�	�j;��R潎�]����M���4T��ב�ɵ���J���(��@�r�S��a��   �   T3B���>���4� =%������:gο�Σ��qx�!�2�z�����2�r��V��8�X���K��f�̇������H�;�uς�Hũ���Ͼr����w������?��.�����ҾH���������@�[a���͒��,�(�y������?#�T����u5��l���F���\3�t�x�m���O�Ϳ%���*&��!$�̿3�XD>��   �   �r �j�����	�)��~�п�嫿H�����K��a��2þ t����9B���k�d\ּ4+(��>���	�-OW�;X��{�ξ�������^5�FH�'�T�tY�	JU�F�I��7�.i�Ģ���Ѿ5��r�[���r����1��.缨��ϥ���G�`Iu��zþDB�tXK�����۪�iOϿ�0�Σ�0�t_��   �   Bn�g����v�J�޿�0ſ���䇉��!W�� �5s�*��R7�bUϽva��3�:k8�RC������`�!>��ַ�.1�i<��\`� ������ڔ��֗��]��՟��F����b�G�>������b���Ozc�:�!����>��o��!d�c!нt7����Opྦ(�J�U��e�����9dÿ}�ܿC�����   �   Sʿ�-ǿ�F���q��4��Ϫ���oR�
�"��9�t����HV�Fj �&	����3�I3��珽���vT�w-��C�G!�MLP��U���������O����ƿ{Vʿ�0ǿ�I��|t���������sR��"�X>�٤���MV�@m �H����3��E3�|㏽ɣ���pT��)��) ��C!�AHP��S��X�������.}ƿ�   �   �ӗ��Z������C��7�b�R�>���¸�l����tc�F�;���=��o��&d�Z&н�7�����t྅+��U�3h������4gÿ��ܿ���l��&p����Nz�~�޿g3ſc��􉉿@%W�x ��v�����7�2YϽ"a��1��d8�l=��$��r`��9��C�澸-��d<�<X`�{��)���ؔ��   �   nY�EU���I�h7�ae����E�Ѿ����[�<����&�1�@(���������J��Mu�~þ�D��[K�v���iݪ�$RϿ�3򿐥�!�|a��t �l����ʷ	�,���п�竿������K��c��5þ�#t�����C��Dk��Rּ�!(�R7����	�9HW��S��ܼξ���Ą�QZ5��AH�2�T��   �   	��������x�����Ҿ<�������hz@�ZW��{ƒ��"���y�X����A#������x5��n��J��L_3���x�V�����Ϳ����'��#$���3��F>��5B��>���4��>%������Eiο/У�Dtx��2�:�����2�t�������X�({K�\[�������Q�;�˂����j�Ͼ��]��t��   �   x;��ہ��5ު��s������gM��e��Ƚ.H_�0��� p�80��;�	�;��U�p�]�Z�������6T�.ّ�����<���K�p�(�� @���S�a�2f���a�ȡT�2A�@�)����U￹p��3[���S����bw��Z�Y�`B߽��-��I����<� _;�㍼.vO��鿽>���H��z}�nr��K\��T����   �   �[��V��F���-�J����ҽ�戽����X����<8��<��<У��8�W�lc��!����ؾC�&�XAq��Ҥ��ֿJ/��h"��5?�,[���r�w���
̄�%���L�s���[�Nt?��N"�t��t�տ�ˣ��Qo�<B%�̑վ>?}���JH��=k��<�<��<����a�(䀽N˽�	��|*�ȁD�}U��   �   kｻz�6;ҽ_ͮ�1���P�0�R�Ф.<hD�<�H(=*u,=���<`s5���r�r�h܏�^��z�7����=����`�.��:/1�r�Q� r�3���C����'��^ǐ��"�� 	r�ЂQ�H�0���α�7"��_����n5�r��ߌ�b��0a�@Î:��=N;=,�6=X�=�;i<����\Ov��p���Oν�c��   �   �
~��s���Q���@j����к$"�<�=��H=�.c=��S=��=���󤂽�#��m��yZ���[B�DR���-��Ul��@����:�.j^�؀��<���Ϛ�旞�B՚��/������Ɩ]���9�v`��0��;��)�����?�}:���������r����:�/=p�b=D�q=�HW=X. =(��<�	�:<>���d��J��o��   �   f�5�*X,�̏�@|�� ��)<�0�<rl3=@c=�dv=&�`=2m= ������t�&�����F��
F��Ӎ��q�����65��h>�B�b�ע������Zi���H���c��"e���Q����a�H$=�~��O#��[Z������RC�1.��UR���K!���x� ";�"=��o=qr�=D>q=v\A=V =�Z[< '��l奼�����(��   �   �
~��s���Q���,j����кX"�<�=&�H=n/c=X�S=��=��j���`#�
m��(Y���ZB��Q��!-��Kk�������:�i^�g׀��;���Κ�����\Ԛ� /������]��9��_��/�;��������?�59���������r����:1=2�b=��q=IW=v. =,��<�	�:T>���d���J�*�o��   �   3k��z�O;ҽfͮ�%���2�(�R���.<�E�<�I(=�v,=���<`75���r�4��ڏ�݁ﾴ�7�Z�������^�����-1�h�Q���q����������%���Ő�!���r�؀Q�0����翲 ��4����l5���u݌�6�+a� 7�:8�=�;=
�6=̵=�<i<����xOv��p���Oν�c��   �    �[�/�V��F���-�F��t�ҽ�戽J���Q����<���<��<�y��(�W�T`����@~ؾ��&� >q��Ф�L�ֿ�-��f"��2?���Z���r�`����Ʉ������s�ʏ[��q?��L"����ɟտ�ɣ��No��?%�k�վ�:}���PBH���i�\�<��<��<�`�0a�䀽S˽ �	��|*�ځD�,}U��   �   �;��灶�=ު��s������gM�qe�ąȽ G_��� ��8���;���p;��N��]�@�������2T��֑�F���6��lI�z�(�@�v�S��a��f�B�a���T��A�R�)����c￁m���X���S�±�[s���Y�7;߽&�-����ص< E_;����zuO��鿽?����H��z}�{r��X\��c����   �   ��������|�����Ҿ5���w���;z@��V���Œ� ��y��ꁼR7#������r5�wj���C���Z3�Єx�����?�Ϳ�����$�( $�ؽ3�4B>�1B���>���4�.;%��������dο�̣��nx���2����6�2�Jl��d��`�X��jK��X�������@�;�˂����v�Ͼ��f��t��   �   yY�%EU���I�j7�_e����9�Ѿ�����[�Ȏ������1�p�4�������D�Eu��wþ9@��UK������ت��LϿ�-�$��X�x]��p �b����X�	��%����пy㫿]�����K��_�j/þt���!<���`�TEּ�(�6����	�HW��S���ξ���˄�ZZ5��AH�=�T��   �   �ӗ��Z��
����C��6�b�N�>������K���$tc����^�=��e�@d��нD�6�&���gl�&���U��c������iaÿV�ܿ���	���bl�����=s���޿�-ſL������CW� ��n��	��x7��MϽa��'�P^8�y;�����&`��9��A�澺-��d<�DX`����.���ؔ��   �   Sʿ�-ǿ�F���q��4��Ϊ���oR��"��9�G���@HV�Ti �/��l�3�;3�dݏ�����pkT�$&��w���@!��DP�LQ���~���﫿�
���yƿ�Oʿ<*ǿCC���n��u��f����kR���"��4ﾃ����BV��e � ��D�3��<3�����	���*pT��)�� ��C!�FHP��S��]�������5}ƿ�   �   Dn�l����v�K�޿�0ſ���⇉��!W�� �s�����7��RϽxa��'�bY8�{6�����]`��5����z*��`<��S`����d���Ք��З��W��-����@��l�b�%�>�6��������mc�$�Q룽�=��c�d��н�7�ϟ��8pྥ(�L�U��e�����?dÿ��ܿI�����   �   �r �l�����	�)��|�п�嫿E�����K��a��2þft�����>���a��>ּ�(��/����	��AW�}O����ξb����V5�%=H�R�T�s�X�+@U�ڗI��7�la�����Ѿ]	��Ŵ[����s��z�1�缨�������F��Hu��zþ>B�sXK�����۪�mOϿ�0�ң�4�x_��   �   V3B���>���4�=%������9gο�Σ��qx��2�U�����2�fo��D����X��SK�O��w��������;��Ƃ������Ͼ �񾿖�7p������ޖ�������Ҿ�}��8s@��K���������yy�,䁼�7#������t5�Vl���F���\3�u�x�p���Q�Ϳ*���,&��!$�п3�\D>��   �   �f���a�ΟT��A�ک)�Ԧ�~�=o��Z�� S�V���u����Y�`>߽��-�@����<��_;Hˍ��fO�࿽(����H��q}��m���V�������5��&|���ت��n��+���_M��^�`{Ƚ�6_��ت� l�8�ڱ;��V;��P���]�����F���4T��ב�̵���J���(��@�v�S��a��   �   �ʄ����z�s�v�[�s?��M"����C�տ�ʣ�]Po�3A%�U�վ(=}���DH� �i�p�<�&�<��<���HFۀ�)�ʽ.�	��u*�~zD�^uU�(�[�O�V���F��-�����ҽ�݈����������<���<��<`n���W�8a�� ���ؾ��&�s?q��Ѥ���ֿ\.��g"�:4?�~ [���r�i����   �   �&���Ɛ��!���r��Q���0�n��翘!��谂��m5�~��rތ�i�h-a��*�:��=�;=��6=R�=�^i<��� 	��@v�eh���FνFZ�Za�q��1ҽ�Į�g~�������R���.<\T�<,O(=�z,=X��< '5�<�r���Dۏ�Ȃ�d�7����R����_�z��X.1�X�Q���q�l���m����   �   p����Ԛ�p/��S���X�]���9�:`�D0�;��������?�&:�����ȝ�d�r� ��:Z1=j�b=�q=*LW=t2 =(��<@��:l0���\�R�J�
�o�^~���s��{Q�&��$[����Ϻ�-�<�=��H=N2c=p�S=J�=���P����#�9m��{Y��[B��Q��f-���k��֍��:��i^��׀�A<��EϚ��   �   �Ҷ�\i��p˥��
��&�z��3P��^)�v��I�Ͽ`���^~W�6��ɺ���;��垽X�����<��Q=t�h=�S=P| =��<`LA;�8��4��j>� @b��mo���d��B��;�`���@�:dn�<=X/K=�`=@�H=���<`�K������.?�ET���t�Y�p����ѿ���t�*�UQ�&�{��V��v���o���   �   ����/X�����ۏ�x�u��mL�,�&�~��z�̿����S�;)��7��"7��u�� !�80�<�D=�-T=Z�7=\y�<��9<�<!��$����J��ꃽ������󘽳>���2Q������A���<@+�<(/=�UK=Z�:=@y�<�UM�Z���u	;�����l��h�U�Ag���1ο��N�'��fM���v��������S���   �   ��������t��*߆�~�g���A�(m�������¿�x��YH�$O�g���|+��֑�X�,��Z�<N~=`�=�q�<`^n;����J�����jν������~����������ҽޠ�b,S�ܧļ@ϵ:lX�<��=�j=TC�< �V��闽p$/��Y����� J�쏐�c�ÿh���!�JDB���g�u܆��U������   �   ����d��jŇ�$Hs�ܥR�V�1�>����� (���}���6�7��y����1���]N��@[<�ם<(V<`*K��0�<m��ĭ�3!�zD�v�`�r�r�)uy���s��Ib�<�F��#����YŨ�$;�зq��u�;  �<�7< u�������*_��+��8�/G�����
��2:��1��pR�V�r�mw��	.���   �   ���kz�k�\iT��9�
���4���Ͽj.��Kh��K �>xϾ�x������j�XW���=������~9��<��$-+�T�e�����NP��\ν��˾��Ͼ��˾d�ʪ��:���i�$a.����x�����@�$���v���t�F3�5{�!Ѿ�5!�):i�r���lп�(��u��9�d�S��Dj�:�y��   �   ��U��Q�RFF���4��F���]�࿻����J��q[E����+���lM�2�ܽ�6S�X�Ѽ�d˼>;�IǮ�X��F�W���3���� ���WJ���:F"�0B���P���/�@�������[���4���pC���ڼ�/��{Z�7SཤoO�84��2��˸E��V���ʲ�[�\���y���3�HcE��cQ��   �   rf/��,���#�:������z㿢���Hx��I`��� �`�پ!��v�"�����`HH�Xo!�"�c�Ҷýb!�l�u�续���澈S��Y.�i/H�Ĝ\�T�i���n��ej�*�]���I�g�/����L�ں��J�x���#�~�ǽ�ij�*'�zuM�����#�L����ھj� �4�_�9���=Ǻ��6�������"�p,��   �   &��
����7c���ֿ�t������tNl�%�0�>���\��\�Q�K����ԏ��O��Nt��6Ľ��"�)�~�����v �|'���O���v�,���5���񢿥��9[���񚿶���]�x�>�Q��(�H���L��H���h�$���ƽ�x���R���5��x�Q����.����/�5k�����^;���Yտ��S�Zo
��   �   ��ܿ�ٿGWο'7���+������&!g�z�3����C��2?s����Ҋ����m��m�!ֱ��2�
�q��5��[���c2��te��댿�������ZͿčؿb�ܿ%ٿ�ZοT:��X.������@%g�Ğ3�(���F��NDs����@���,n���m��ѱ��.�5�q��1�����1`2�`pe�Y錿�󥿾���WͿ�ؿ�   �   h��X���돍�b�x���Q�~�(�r���H��$����$�D�ƽ�x���R�0�?;���Q��������, 0�)k�����3>��7]տ���U�dq
�8
��
�����f���ֿLw������Rl��0�^����_���Q�t����Տ��O��Gt�&0Ľ��"�5�~�b����s �Jx'�`�O���v�P����1��l�   �   �n�2`j��]�܆I�F�/�h���F�<���H�x���#���ǽ�aj��'��vM�3����#�����Wھ�� ���_�M ���ɺ��9⿔�����"��,��h/��,���#��F���}�꠻�#z���K`��� �m�پ#����"������GH�"j!��c���ýt\!�ۛu���������O��U.��*H���\���i��   �   �A"��=������o)�����k���[����X���teC�`�ڼ ,�~Z��V��rO��6��	��R�E�%X���̲��]�؋��{��3��eE�fQ�0�U���Q��HF���4�jH�(���࿅ ��KL���]E�<��-��oM�p�ܽ�6S��Ѽ�U˼&�:����������W�T��~���5��]��NF�����   �   ��Ͼj�˾�达CŪ��5��~i�|Z.�#��p��4��0�$� ͍�8u��tt�5�U{�m#Ѿj7!��<i�����Tп�)�Xw��9���S��Fj���y�̫��nz�Tk�PkT���9�L���5���Ͽ�/��Mh�UM �zϾ3x������j�|R�� ����������0����,&+���e������J��iȽ�c˾�   �   �ly�S�s��Ab��F���#��
��(����;��q�p��;�
�<87<`u�y���[��`��L��8�5H��8�����8;�V�1�DrR�P�r��x��H/��?���Pe��}Ƈ��Is�B�R�h�1������!)��h~���6��8��z�������PWN�HP[<\�<�z<��J�r�0��c��:���,!��wD�R�`���r��   �   ,�����إ���ҽ ֠��S��ļ��:lf�<��=n= F�<X�V�뗽�%/��Z�����I!J�����c�ÿ���X"�LEB���g�@݆�V��������������u���߆���g�b�A��m�����6�¿5y���YH��O����`}+�Bב���,�`�<|�=H�=|��< �n;�����J�8����`ν��������   �   �/:��L*Q� ����A��<�3�<B+/=XK=��:=�y�<�XM�^���Z
;�b������!�U��g��y2οP��ƒ'�>gM�J�v�S����~T��1����X������ۏ���u�nL�n�&������̿��S�S�e)��7��G7��u���!�83�<D=�0T=H�7=(��<��9<� !������J��僽�����   �   �mo���d�F�B�$<����� ؆:�m�<�=�.K=4`=ʽH=���<��K�;���/?��T������Y�����ѿ�����*�"UQ�D�{��V������o���Ҷ�Ui��e˥��
���z��3P��^)�^�� �Ͽ<���%~W�	������;�v垽H�����<`�Q=��h=d�S=�| =d��< PA;�8��4��j>�@b��   �   @:��V*Q�����A�P�<4�<�+/=�XK=|�:=�|�<`PM�����	;�k���=�� �U�g���1ο����'�BfM���v���� ��tS��#����W�����ۏ���u�mL���&�"���̿W��V�S��(��6��7�t��X!��5�<�D=n1T=��7=d��<��9<� !������J��僽�����   �   >���������ҽ ֠��S���ļ@��:�g�<��=�o=(K�<x�V��痽`#/�#Y��8��^J�h�����ÿ���� �|CB���g��ۆ��T�������������s��bކ�<�g���A�fl�l�����¿�w���WH�JN�1��{+�6ԑ�x�,��d�< �=2�=p��< o;�����J�K����`ν��������   �   �ly�h�s��Ab��F���#��
��
����;���q� ��;�<h7<�t�,����^����p8�gF��� �����Z9���1�:oR���r�Xv���,�������b��Fć�0Fs�F�R��1�@�����&���|��f�6��4�Vx�����p���AN��][<��<�<�J�,�0��c��F���,!�xD�h�`� �r��   �   ��Ͼx�˾�达JŪ��5��xi�lZ.�ܴ�o�������$�0����g��2t�1�T�z��Ѿ?4!�98i�*����п�'��t�`9�n�S�:Bj���y�`��Jiz��k�DgT�H�9����r3��Ͽ�,���Hh�5J ��uϾIx�Ġ���j��E��@��������o0�����.&+� �e������J��zȽ�u˾�   �   �A"�>������r)꾼���b���[�^��s����bC�$wڼ��sZ�&N�\lO��1������E�U��ɲ��X� ��<x��3�aE�aQ�
�U���Q��CF���4�E�V���࿳���BI���XE����(���hM�ܽ,S� �Ѽ�L˼|�:�߽��R����W�W������@��e��YF�����   �   *�n�<`j�!�]�߆I�H�/�i���F�+����x�(�#�%�ǽ�\j�v'�tkM����P�#������ ھ3� �G�_�]����ĺ��3�F���z�"�4,�$d/�|},�l�#�J������w����7v���E`�B� ���پH��d�"�����<H�
c!���c���ý\!���u���������O��U.��*H���\��i��   �   m��X����c�x��Q�{�(�j���H��𬀾n�$��ƽ��w���R��落/����Q�u�����=�/��k�X����8���Vտ���Q�Zm
���
�����_��ֿ�q��V��|Jl� �0�vz��sY��"�Q�P����͏�|�O��@t�.Ľ[�"���~�P����s �Mx'�f�O���v�U��� 2��r�   �   ��ܿ�ٿKWο*7���+������#!g�r�3�����B���>s����������m�2�m�˱��*���q��-�����\2�Ole��挿	񥿜����SͿ��ؿ��ܿ�ٿ�Sο�3���(�������g��3�Σ��>���8s����H�����m��m��α�.���q��1�����1`2�epe�]錿������WͿ!�ؿ�   �   *��
����:c���ֿ�t������oNl��0����\����Q�����TЏ�<�O��;t��(Ľ�"���~�����p ��t'�#�O���v������.��F뢿/���T���뚿���5�x�q�Q���(�`���C��|����{$�¥ƽ��w���R��ꐽ?3����Q�Y������/�7k�����c;��Zտ��S�^o
��   �   vf/��,���#�<������z㿠���Fx��I`��� �1�پ� ��_�"� ����=H�v_!�>�c�ɦýW!���u�`������\L�nQ.�&H���\���i���n��Zj���]��I���/�����@�=���p�x���#�R�ǽ�Rj�T'��jM������#������ھc� �4�_�;���?Ǻ��6�������"�t,��   �   ��U��Q�TFF���4��F���\�࿻����J��i[E���@+���kM�l�ܽ.S���Ѽ�@˼��:��������W���������Æ�_B�����="��9�����"����������Z�z��ƕ���VC��gڼx�ZsZ�yP��nO��3��&��ȸE��V���ʲ�[�^���y��3�NcE��cQ��   �   ���kz�k�^iT��9�
���4���Ͽi.��Kh��K �xϾWx����\�j��C��@_��������f(��_�罎+��e�􈏾�E���½�A˾7�Ͼ4�˾�⾾ǿ���0��i�jS.�����f�����p�$��~��Lc��t�=2��{�� Ѿ�5!�*:i�s���nп�(��u��9�h�S��Dj�<�y��   �   ����d��kŇ�$Hs�ܥR�T�1�>�����(���}���6��6y��[������AN��h[<8�<�<�J���0�kZ��8��&!��pD�b�`���r��cy�԰s�r9b�`�F�Ȼ#�����P���2;�XVq�`�;��<8-7<��t��������^����8�/G�������4:��1��pR�X�r�nw��	.���   �   ��������t��*߆�~�g���A�*m�������¿�x�� YH�O�G��R|+��Ց�@�,��g�<0�=4�=x��<@�o;�㱼��I�M����Wν��������z�E��қ��|�ѽ�͠�S�,xļ�>�:|w�<��=�s=PP�<��V� 藽�#/��Y����� J�폐�e�ÿj���!�JDB���g�u܆��U������   �   ����.X�����ۏ�x�u��mL�,�&�~��z�̿����S�5)��7���7��t��!�p6�<6D=�3T=��7= ��<�:<�!����Z�J�6ჽ�����鞽2阽C5��P!Q��{��A��<>�<�//=�[K=��:=��<�LM�����<	;�����j��g�U�Bg���1ο��L�'��fM���v��������S���   �   �B��q����0���֝����A]�3��4�Hwۿ펢�j�d��8��u��xL��y���ڍ��<t>=�`V=&{@=��
=���<�|��g��`)��Gb�����%��V2��F�d�p*,��ȼ`��"w<��=�<=��Q=��9=�<h����Z���mN�����8�f�e��b���ܿB����3���]��_��a��^E�������   �   �ܿ��N��k$���R��8J���Y��0����2�׿͟�Ӑ`�kZ�ｵ�K�G�rұ���(�<�0=��@=�K#= $�<��;�f���' ��p�����U��[�������阽�fs�4�#�쾕� �x;8J�<�=�5<=�+=�<����囵�J��<��XP�?�a�����0�ؿ�u���0�T�Y�ǅ��?t���-���L���   �   ����Ѯ�<���h`����v��FM��?'��1�AtͿ�ė�(�T�H�l��0};�И��dȔ��D�<�=@n�<j�<�kW��o����p��e��+h潗��l�=��Z��n��$S�e���::u��
��`ȑ�h	�<�
�<�n�<�<Գ��N ��z�=�H^�������U�_k��R9ο��Ȭ'��M�Xw��_����n����   �   ����?���J�� ���,�_�ȝ;�H��b������3%��RB�zI��}���(�O�������p��;��V<�:;p���|�V�%���6�Zj0��gU���r�*Ⴞ!>��f!���s�b�V���1���4̼�&�[��Ǯ��V�:`�C<���;���3��d�*����:�����B�񞋿�������Z��;��{_�����_���ś��   �   ���ӥ���Rz�_a�ND��J&��	���ڿo����u�:e*�N�ݾ녾KS�S����˼�(��&{�<s��r�����;���x�Y���t����˾(�ؾU�ݾ0Bپ¬˾�e���t����z��<�����5���i$��Ԇ�n+�@eռ6������N͆���޾P�*�U�v��O���ۿ^	��&�f�C��`���y��|���   �   j#c��^�&�Q���>���'��.����L���a����/Q�e��S�����^��6��0$y�v�	�(��\�`���Ž�8���i��j��q ̾����A]������(��?,��(��9��������|M;�{����k��� �XȽ��d��
����BT}��|��	�_�q*����`oQ�A��y���#f�R���R'�->��^Q��e^��   �   �K9��6��},�������8�U�ſ����g@m�#�*�B辬{��X�1��Ƚ��l�V�D��W��
m۽�0�n����j������!���N9�gT���i��xw��M|�I�w��[j�{*U�R:�ُ���� ��Ē��B�1��{ݽ���z�G���o��Hʽ`I2�;Δ�x�<�*��m��^��Pſn��lA��S��,�N�5��   �   L��F���
�,���t�ῇ�������y�+>;�<�����b�z��5䣽tQt�sq��Dt۽��1�"�����Ǿ�	�2���\�����|Ɣ��뢿@����.��e8���V���K��I����]���2�b�	���Ⱦ1)����2��ܽl��"�u�ϓ����V�b�����8��:�`y��'��b��>�����n
����   �   �H�}��ٿǿ���i��� !t��+>�P����ž�؂���#�Z�ǽ��� k��0�ǽ�J#�:���+5ž�y���=��4s�>���X���lƿ��ؿJ-�dL�π�aٿVǿ�	������L%t�%/>������žvۂ��#���ǽπ��Fi��w�ǽ�F#�*����0žw�<=�20s�����U��/iƿ�ؿs)��   �   +��5���S���H���F��5�]��2�i�	���Ⱦ�%��V�2�K�ܽLi����u�g������b�\�����F�:��y�*��e���������p
�:��~��j���
��������N������ݯy�A;�8>����ޑb�����壽fOt��m���m۽��1�z�����Ǿh 	�2��\�ܼ��zÔ�H袿�����   �   CH|���w��Vj��%U��:�"������)z�������1��tݽZ	��ГG�&�o��Kʽ�L2��Д��{�޺*�rm�$a���ſ���8C��U��,���5�PN9�6��,�������;￺�ſ~���sCm�k�*�OE��}��̑1�%�Ƚ(�l��D�QR���d۽4�0�t���Te��B���@��wJ9�bT�P�i�2sw��   �   R;,���(��5�%��+����G;�v��2�k��� ��OȽ��d���
�����V}�1���b�_�-���	�rQ���������h����nT'�X/>� aQ��h^�>&c�ֺ^���Q��>�T�'�(0���-���� ���1Q����p���z�^�H9��|$y���	�(����`�r�Ž�2���i��e��n̾����TY�����(��   �   ��ݾ�;پ��˾�_���o���z��<�.��O-��D]$�DĆ� \+��cռ��������Ά��޾%�*�ҏv�7Q���ۿ�	�!&�J�C�^�`���y�Q~������C���vUz�Daa��OD��K&��	�a�ڿ�����u��f*�=�ݾB셾uT��S�� �˼8�� {��e��i���� �n;�ʹx�4��������˾��ؾ�   �   �9�������s���V���1�H���¼���[�X����e�:h�C<�
�;4�������*�����v���5�B����������n�N�;�J}_��������1Ǜ�������L�������_��;�*�������� &��zB�K���}���(�����@���@��;h�V<`�:;ܜ���V���(�Oc0��_U� �r��܂��   �   ����|�>���I������+u� ���P|����<x�<4u�<�ń<����!���=�r_�������U�/l��]:ο�����'���M��w��`�����|�������Ү�#���)a���v��GM�*@'�"2��tͿŗ��T���
���};����Ɣ�(J�<J�=�z�<dz�<@�V�TV��rqp�]��j^�P�����   �   �U������嘽�]s�\�#�p�����x;�R�<b�=48<=�+=��<����
J��=���P��a� �����ؿv�*�0���Y�3����t��.��1M��ݿ�-O���$��#S���J���Y��0����{�׿@͟��`��Z�!���n�G�^ұ�L ��D�<00=��@=�O#=x.�<�5�;�W��� �pp�|������   �   %��^2��|�d��*,���ȼ���� w<�=d<=~�Q=x�9=��<,���][��YnN�G���8���e��b���ܿZ���3� �]��_��q��iE��Ť���B��k����0���֝����A]��3��4�wۿɎ��-�d�a8�du��L�y��ٍ�<�<zt>=\aV=�{@=$�
=���<�|�g��F)�zGb������   �   �U������嘽�]s�f�#�h���`�x;\S�<��=�8<=�+=`
�<ؓ��D����J��<��&P���a�l�����ؿlu�b�0��Y�|����s��	-��L���ۿ�N���#��AR���I���Y�,0�^����׿�̟��`��Y�"���"�G��б���� �< 0=(�@=�O#=�.�<�5�;�W��� ��p�����,���   �   ����|�L���I�����+u�����py�� �<t�<tx�<�ʄ<Ȭ��z��\�=��]��q����U��j���8ο���&�'�
�M�*w�_��.~��m�������Ю�@����_��|�v��EM��>'�1�;sͿ�×��T�b�&��T{;�镧����4O�<Ԙ=�|�<p{�< �V�0V���qp�#]���^�b�����   �   �9�������s���V���1�D��{¼�^�[����� ��:��C< (�;č��H����*�垛�����n�B� ����������t���;��y_�����.��ě�S�������I�����n�_�n�;�8���������$$���B�'G��^{����(�Z��� ������;8W<��:;|���̔V���*�\c0�`U�9�r��܂��   �   ��ݾ�;پ��˾�_���o���z�
�<����,���[$�����J+�Vռ`���`���ˆ�u�޾��*�O�v�JN��ۿL	�$&���C���`�F�y�l{������]���<Pz��\a�*LD�"I&��	���ڿ�����u�ac*���ݾ#酾aP�?N��|�˼` ���z�*d�Ti���� �m;�ҹx�>��������˾��ؾ�   �   \;,���(��5�+��2����G;�v���k��� ��NȽ��d��
�H��K}�Iw����_�(��T�mQ��	�������c�����P'�+>�&\Q�
c^�� c�\�^���Q�º>���'�*-����+��������,Q�h��s���Ŭ^�o0��
y�X�	�����~`���ŽL2���i��e��s̾����\Y�����(��   �   OH|���w��Vj��%U� :�#������z��������1�Hsݽ ��^�G���o��Bʽ�E2��˔��t��*��m�]���ſ�}?��Q�~,���5�RI9�>6��{,� ��*���5￵�ſc����<m�{�*�%>��x���1�A�Ƚ��l�~xD�P��pc۽֜0�Z���Ke��C���D��}J9�#bT�\�i�=sw��   �   %+��5���S���H���F��6�]��2�c�	���Ⱦ�%����2��ܽ�e����u�⍤�3���b��������:�� y�G%��U_���i����l
�������v�
�d����ῐ������y��:;��9����t�b�P��Lݣ�VDt�>j��hk۽��1�P�����Ǿd 	�!2���\�߼���Ô�O袿�����   �   �H�}��ٿǿ���j��� !t��+>�F����žz؂���#�)�ǽ�z��ec����ǽ&B#�1����,žSt��{=��+s�����R���eƿ_�ؿ�%俥D�-y�ٿ�ǿ�������gt��'>�[��>�žjՂ���#�{�ǽ&y��Cd��M�ǽ�E#�䇂��0ž�v�<=�60s�����U��5iƿ��ؿz)��   �   P��H���
�/���v�ῇ�������y�#>;��;�O���b����ߣ�Dt�}g���e۽b�1�����Ǿm��k2�{�\�F�������&墿�����'���1��qP���E���C��{�]��2�1�	���Ⱦ"����2�r�ܽb����u�{���i���b�����,���:�ay��'��b��D�����n
����   �   �K9��6��},�������8�T�ſ����a@m��*��A�W{��<�1�x�Ƚ��l��tD��K��3\۽��0�����s`��+������,F9�E]T��i��mw��B|��w�&Qj�� U��:�?��z����t��������1�kݽ�����G���o��DʽDH2��͔��w�5�*��m��^��Rſr��lA��S��,�T�5��   �   l#c� �^�&�Q���>���'��.����N���`����/Q�S������^�	4��Ly�H�	����s`�f�Ž�,��i�8a���̾����U�^����(��6,�F�(�o1�;��)����A;�q���k��� ��EȽ0�d�
�
����dK}��y��*�_�5*����\oQ�B��{���%f�R���R'�"->��^Q��e^��   �   ���ԥ���Rz�_a�ND��J&��	���ڿo����u�1e*�#�ݾ�ꅾ:R��O��Ȼ˼�����z��W��`�� � �v;�\�x�F������}˾�ؾ�ݾ!5پW�˾1Z��|j��<�z���<�$���#��"N$�����3+�Qռ��������̆�k�޾H�*�U�v��O���ۿ`	��&�h�C��`���y��|���   �   ����?���J�� ���,�_�ȝ;�H��b������1%��KB�_I���|��`�(����� ��� ��;XW<@I;;؃��x�V�Y鹽[��\0�YXU�ƶr�=؂�5��v���s�ĎV��1�,�L�����[����� ��:PD<�H�;���������*�ܟ�� �����B�𞋿�������Z��;��{_�����a���ś��   �   ����Ѯ�=���h`����v��FM��?'��1�@tͿ�ė�%�T�@�K���|;�G������ R�<(�=���<,��<@(V�D>��cp��T���T�,��u���^w��}��?�;����u�����%���)�<�#�<\��<pЄ<t������ �=�'^�������U�_k��S9ο��Ȭ'��M�Xw��_����n����   �   �ܿ��N��j$���R��7J���Y��0����2�׿͟�Ґ`�fZ�ཱུ��G��ѱ�|�����<X	0=��@=NS#=�7�<0c�;�J��� ��p��������P��k������NTs���#������Gy;�]�<��=�;<=0+=��<����$����J��<��VP�=�a�����1�ؿ�u���0�T�Y�ǅ��At��-���L���   �   	����0������[���!F��("b�\�6�V���߿ܥ���i�W��D��ztR�&2���n���f�<�6=��N=��8=*f=|a<��ӻL�ؼ��5�DMo����Z|��*��~�o���5��ټ��׻�M_< �=v�7=��M=�X5=�}�<`쩼�8��<S�"��������i������߿��X�6�h)b��H��+��������0���   �   Ek��̿�Oe������Z����]�^�3���0ܿ�	���ce����u���N��p���}����<��'=~�8=�=0��<��;�����-���}��ޞ�}P��]`��(^��5����5~��b-����� 6;�r�<.;=�
8=��&=�3�<骼or����N�DȺ�i���e�� ��R,ܿ ���3���]��]�����Nf��u̿��   �   �m��	���w�������G|��|Q��x*�ȳ��eѿ�њ�z8Y��K�0|����A�����`�w<(��<��<`�<��Ļn��#�*���6A��s�j��Xn�z��_���g�k���
������ɻ@�|< ��<ht�<er<8A���ఽ�B��ɯ��u��cY�3皿zѿ��f�*��Q�xL|�Ó��x��r	���   �   2v����I��������#d��-?�l��>�������Eꍿ11F�M�7����{.�e砽�ƽ��Β;�U/< �x9�P��D9e�,�½� �~6���[�WWy�8�������;���ey���[��.6��<���½��e����� 008�p+<O�;<���v����.�
ٞ��>�XF�|�������[�� ���2?�B'd�����ל��(����   �   =���x������4�e���G�v1)�&s���޿-*����z��.���⾩���Hf��Ȑ���㼘�E��ٔ��,�v���" �((A����S���Z����Ͼ`�ݾn��K�ݾH�Ͼ~��Y������DA�v��ۥ��-��r���zI��Q�������Vŉ��6��%.�B�z�J9���޿rx�R5)�J�G���e��������   �   �g�$!c��U�vB�z�*���-��b迿/���LU����#꽾h�d�5<��#���(�� �D�n�4vν��$�c�p�����q3Ѿ����Е��6"��9,�A�/�<,�r:"���/���q?Ѿ������p���$��ν�Go� ��j��#��/����Ke����)��
fU����m��𿨆��*��B� �U�
!c��   �   �<�xK9��d/��b �|������ȿ~Q��J�q��.��B�4����6�U�нPz��^Q�1|���4�N6��k��&��a���.R��[=�P�X�T{n�iG|������I|�1n�E�X� a=�"W����N-��r��x\6�YZ�)���p�Q�<{�7ѽ�7�T@��/j��*.�u�q�zX����ȿ_������b �Dd/�,K9��   �   0%���F��c��_�<Ŀ�C���~�ߵ>���� 	��	Zh�F0��ꪽ:����Y���㽒`7��4����̾�,�~6�Va��s���������R+���K��],����������u��hYa�U6� -�v�̾h2��*^7��㽇p��EȀ�+���Y���h��"��F����>��	~�HF��Ŀm_� c�������   �   WL�G��ܿm>ʿ�ϲ�+���>x��A����%�ɾ䅾�+(�BϽ5͏��؏��7Ͻ�E(��Q�ɾם�V�A��Dx�H��Ѳ��?ʿ�ܿ�I�KP��J迾�ܿ�Aʿ�Ҳ����WCx���A�>���ɾ�慾b/(��ϽΏ�׏�03Ͻ�A(�������ɾޚ���A�@x�����Ͳ�}<ʿY�ܿ�E��   �   �H���(�����쾗�s���Ta��
6��)���̾/���Y7�W���m��(Ȁ��-���\�r�h��&�����"�>�(~��H��""Ŀ�b��d���Ԍ�n'�:��R	�~e�,c�!ĿF��r~�ܸ>����7��^h��2�H쪽1���V��A��\[7��0����̾d)�u6�EQa��p����������'���   �   ����C|��yn�Q�X��\=�^S�����a(��_n��W6��R佹�����Q�v{�X:ѽ7��B��n�j-.���q��Z����ȿ������d ��f/��M9���<��M9��f/��d �8��u��W�ȿxS��e�q��.��E�]��Y�6�y�нdOz�jYQ��v���,�H6�wg��� ��˃��<N�DW=�8�X��un��A|��   �   ��/��7,�26"���N����9ѾĲ���p���$���νB<o�v��R��1$������*Oe�� �����hU�˰���������B��Ж*�FB���U��#c���g��#c���U��B�D�*�������L꿿����]NU�'��L콾��d��>��O���L���R�n��lνR�$�A�p�����O-Ѿw���ё�K2"�v5,��   �   ��⾨�ݾ �Ͼ���H���t���=A���ӥ��{-�b���hI��O�W�������Ɖ�a9��'.���z��:���޿�y��6)�<�G���e�ԏ����ʼ������(��n�e���G��2)�<t���޿�+����z�N.�{��܊��zg�ɐ�\���uE�`Ɣ�0�,�1��� ��� A�������z��~�Ͼ��ݾ�   �   ���D7���\y���[��'6��6���½�e����� �R8X�+<`e�;X���¡���.��ڞ�@��YF����������8��
4?�)d�����&��������w��P�����������P%d��.?�T����������덿`2F��0����|.��砽Lý���;�p/< -�9�6���(e�Ւ½��P6���[��Ny��3���   �   �h����|�^�䷺�t������Oɻ�}<���< {�<kr<`B��QⰽB��ʯ�fv�
eY�蚿&{ѿ���>�*�*�Q��M|��Ó��y���
���n�� 
���x��m�.I|��}Q�$y*�B��Kfѿ-Қ�C9Y�FL��|��%�A��X	����w<��<���<`�<VĻ~���A���G7�fn�����   �   �Z���X��B����,~��Z-�@��� �;�{�<�>=�8=�&=L4�<�ꪼ�s����N�ɺ����ʒe�w!���,ܿd����3�h�]��]��5���f��	Ϳ��k���̿��e��^��E[��,�]���3���|ܿ
�� de�1��v��N��p���{��0�<��'=�9=�=�ȸ<�A;���F�,���}��ٞ�$K���   �   a|��*����o���5���ټ`�׻HL_<��=�7=p�M=ZX5=�|�<�9���S�j������!�i�D�����߿��v�6��)b��H��;���Ï��1��	���|0������J���F��"b�@�6�<����߿Xܥ�y�i�&���C��tR��1��8m���g�<l�6=(�N=�8=~f=8}a< �ӻ��ؼd�5�Mo�����   �   [���X��O����,~��Z-�L�����;|�<�>=|8=��&=�6�<h檼�q��P�N�Ⱥ�7����e�� ��,ܿʢ�Ƙ3�R�]�?]��I���e���˿��j��o˿��d��s���Z���]�܏3�����ܿ]	��ce�p��u���N�o���w����<��'=B9=H=ɸ<�B;���R�,��}��ٞ�:K���   �   �h����(|�)^��x��x��`Mɻ}<���<X~�<`ur<(:��߰��B��ȯ��t�cY��暿ayѿ����*�,�Q�DK|�R��w��l���l�����v�������F|��{Q��w*� ���dѿ�К�;7Y��J��z����A��믽����w<d��<���<X	�<�SĻ\���P���]7�vn�����   �   ���P7���\y���[��'6��6���½��e�H��� �W8X�+<`��;ؘ������N�.��מ�>��VF����������	��6��n1?��%d���������ʒ���t����������e����!d�,?�T������:���1鍿�/F������zy.�`㠽Է����;�y/< ؁9 5��6(e���½��X6���[��Ny��3���   �   ��⾸�ݾ�Ͼ���Q���v���=A����ҥ�z-��\��xWI�4B��{��f���É��4�w$.�4�z��7��T�޿^w��3)���G�N�e�j������������������e���G��/)��q���޿�(��6�z��.���⾲���Pc��Ð���㼸dE� �����,�Ȋ����� A���� ��������Ͼ��ݾ�   �   ��/��7,�:6"���V����9Ѿ²����p��$���νp9o�������]������PHe�n��|���cU������𿿁��4���*��B���U�@c�&�g�Lc�|�U�0B���*�z�����7濿r���dIU����9罾"�d��5��y���������n�"lν�$�)�p�����R-Ѿ����ؑ�T2"��5,��   �   ����C|��yn�X�X��\=�aS�����V(��En���V6��Q�a���0�Q��{�J1ѽ@7��=���f�d(.�Y�q�V��p�ȿs��@���` � b/��H9�v�<��H9�Pb/��` ����a��?�ȿKO��ȕq��.��>�H����6�k�н�Cz��QQ�~t��;+佬G6�\g��� ��̃��>N�JW=�@�X��un��A|��   �   �H��)�����𾗿s���Ta��
6��)���̾�.���X7�&��6j����%��]V��h������ν>�~��C��PĿ,\�(a���r���"�؈�0��a�v\�:Ŀ-A��f�}���>�4��X��vTh�,��㪽����wR���㽵Z7��0����̾`)�v6�HQa��p����������'���   �   ^L�G��ܿq>ʿ�ϲ�-���>x��A������ɾ�ㅾ�*(�Ͻ)ȏ�я�K,Ͻ/=(��텾��ɾ$���A��;x�����ʲ�&9ʿ��ܿ'B�kH�C�\�ܿ�:ʿ_̲�j��Q:x�D�A������ɾ�����&(�LϽJƏ��я��/Ͻ�@(�������ɾך���A�@x�����Ͳ��<ʿ^�ܿF��   �   4%���H��c��_�>Ŀ�C���~�ڵ>�������6Yh��.�V檽y����O��R��V7�W-��,�̾Z&��6��La�"n������m���$��E���%��H
��仗�Mp��Pa��6��&���̾*+���S7�a��tf�������&���X���h��"��7����>��	~�IF��#Ŀr_�c�������   �   �<�zK9��d/��b �~������ȿ~Q��H�q��.�yB������6���н�Dz�0NQ�p���#�@B6��c������}��zJ��R=�N�X��pn�<|��|��+>|�[tn�@�X�,X=�nO����#��8j���P6�3I�	�����Q��{�p3ѽ�7�@��j�*.�s�q�zX����ȿ`������b �Hd/�.K9��   �   �g�&!c��U�xB�|�*���.��c迿/���LU�x���齾��d�T9��������d�@�n��cνR�$���p�����t'Ѿ������."�1,� �/�3,��1"���5���t3Ѿ������p�8�$�j�ν�,o���������K����Je������fU����n��𿪆��*� B�"�U�!c��   �   ?���y������6�e���G�x1)�&s���޿.*����z��.�W��X���2e�(Ő���㼠RE�����:�,�4���h���A��������	��F�Ͼ�ݾ���ݾ��Ͼ������r��/6A���Rɥ�Nl-��I���?I�=�p|�����ŉ��6��%.�@�z�L9���޿tx�T5)�L�G���e��������   �   1v����J��������#d��-?�l��@�������Fꍿ-1F�@�����:{.��䠽Է��`#�;p�/< *�9X���e���½��k6�ݍ[�Fy�/��d{���2��=Ty���[�� 6��0�U�½��e�r��  8��+<У�;�������P�.��؞��>�XF�}�������]�� ���2?�B'd�����؜��*����   �   �m��	���w�������G|��|Q��x*�ȳ��eѿ�њ�x8Y��K�|���A�$�0����w< ��<8��<,�<�Ļ<��p��~���-�+i�B���b�R���v�6T����x�vx�P�Ȼ�:}<0�<L��<��r<�7��M߰�-B��ɯ�~u��cY�4皿zѿ��f�*��Q�zL|�Ó��x��s	���   �   Fk��̿�Oe������Z����]�`�3���1ܿ�	���ce�����u���N�p��y����<�'=�9=�=Ҹ< �;H���P�,���}��Ԟ��E���U���S��*`#~�BR-�<�����;̆�<C=�8=\�&=L:�<p䪼�q��t�N�6Ⱥ�f���e�� ��T,ܿ����3���]��]�����Nf��t̿��   �   �?��B���A��0��vY����]���3�>��Y_ܿCC����e��r���~�M�eO���M�����<�:=:�R=�<=V"= �x<0u��&ȼ��+�ndd��$���#��`����~b�\e)�L¼�������<+
=�?=�=U=�==d�<(^���t����L�T����\���d�a����ۿ`9�T3��A]�%��B՝��.��ڝ���   �   �ٿ�$I��N)��(o�������Y���0��e���ؿ�u����a���1඾�yI�V����I�����<t,=��<=�e=H;�< �~;��� �#�v$s�:И�����W��8#��b̗�dqp�֖ �X~�����;X��<�Z"=��?=��.=��<\q��3Ȳ��BH����}���`�ܟ�j�׿���	0�|Y�.I���P��"��L���   �   �������{��
[���v�$�M�ڞ'�|���ο�N��$�U�Y������=�@(��l����6�<PU�<��<D3�<�򍻸5����t��p��f+�0x�6w����$!���*������ q�����@c�H��<4b�<_=�x�<p����~��M�;� F��K-���T�fҗ�OͿ\5�A'�4FM�V�v�e^�������ή��   �   ����u����,����q_���;�������D{������w�B�MQ���P���7*��=��|ǭ����;�KG<@F�:ȧ��ʀ[�$���o���1��V�0�s� ��H9��>�����r��uU�0�:8��?��EW�02�� �+; �R<���;8���ƙ��O)�����6���
*B�C1��E���������;��_�״��3H��G���   �   ����y���y���`���C��&��	��ۿ�8���`v���*��|޾�����c��9���Ҽ��'�dU����#���q�&�<��qz��c��FU���˾*6پ��ݾ��ؾ�˾Q���u���E�x�g7;�\"������  �`l~����μ�������X����ݾN|*��v����|�ڿ�	��H&�NJD�Za�Mz�Ƣ���   �   �c��_^��XQ��&>��K'����mU쿚{�������JQ�(���깾6~_�����!|�p���

�gd��ȽT� ��k�Pj��?:;^������ 0���(�h9,�N�(���� ]�N���:%̾hq���j�<M�A�Ža�Bb�
�F z�������^�ө��9��^>Q�X��)����� ,�n�'���>�H�Q��^��   �   zF9�R�5�� ,��N�><�uſ`Q����l�"�*��B辺����1�k�ɽ�o���F�hφ�-Jݽh�1�Z���p��������:��U�iOj�0�w��D|�rw�'�i�VdT�bM9�6�������i�����f�0��۽�~����D���m�-,ɽ��1������Z���*��Em�����V�ſ�2￦�����>x,�6��   �   �������j
�������Z�����G�x��:�s���Բ�\cb����?��vyu��D��)�ܽ|�2��#���Ⱦ�	���2���]�B��2D��1O��Y1��v(��Z����碿vÔ�򼂿��\��2����q�Ǿ<}��
�1�Jf۽Dv��Ƃt����_��t�b��"��A��?;�<�y����������Q���X�
�@��   �   �@��"�r�ؿPdƿQ�����O%s�vs=��j�ž�r��##�idǽ
L��Ix����ǽ��#��߂���ž~��I*>��t���������ǿ^ٿ@x俿D迻&��ؿ�gƿ�S�����)s��v=�xm��žQu���&#�hǽ�L��zv��5�ǽ��#��܂�3�ž����&>��t���������ǿ�ٿft��   �   %������䢿����[����\��2������Ǿ�y����1��`۽s����t�v��+���b�&��|C�C;�a�y�3�����W�����h�
�l������l
�������\��!���x��:�����ײ�Ngb�>��A��lwu�DA����ܽ^�2� ��&�Ⱦ��	���2���]�P?��/A���K���-���   �   ,?|�xlw�ܷi�z_T�I9����o���$e��_����0��|۽jz����D�ښm�`/ɽ �1�&����^��*�jIm�ʢ����ſ�5�v������z,��
6��H9���5�&,��P��=��w�ſSS����l�m�*��E�؟����1���ɽ�o��F�ʆ��Aݽ��1�^����j��8������:��U��Ij���w��   �   �4,��(����NY�����y̾�l��|�i��G� �Ž�
a��[���
��"z�E���� _�t���"���@Q���L���~�쿰-�R�'��>���Q��^�\ c��b^�8[Q�)>�~M'�*���W�~}��P���MQ�����칾_�S����!|�����
�RZd��Ƚ*� ��k�Le��64;X�������+�N�(��   �   N�ݾr�ؾ�˾����~�����x�s0;���?���| ��K~���μA���X�����*�ݾ~*�v�7��w�ڿ�	�(J&�0LD�d\a��Oz�=�������{����y���`���C�\&�		�cۿQ:���bv�N�*��~޾ډ���d�C:���Ҽ�'��B����#��蟽�k�ǭ<��hz��^��|O����˾�/پ�   �   �4���ۂ�q�r�nU�Jx0�l2�6���5W������,;H�R<���;H����Ǚ�?Q)����m����+B�Q2�����ˊ��&��ܝ;�ė_�쵁�vI����������Û����+���s_�Ҥ;����L���X|��υ����B��R���Q���8*�P>��(ĭ� ��;�fG<�y�: ���Tp[��i���1�'}V���s�����   �   ����������潺���v�p�̐�� �b����<�l�<Rb=`{�<x��������;�IG��'.���T�3ӗ�U�Ϳ 6��A'�HGM���v�B_�������Ϯ���������{���[��F�v��M�~�'�����οO���U�ܴ�B��T=��(��,���L<�<^�<|��<�C�<`�����\�t�h���!��r��q��   �   zR�����Ǘ�|hp��� ��p�� ߙ;$��<
^"=��?=�.=L�<�r��8ɲ��CH����D~�I�`��ܟ��׿d��D
0� Y��I��xQ���"���L��ڿ��I���)���o������Y���0�0f���ؿ0v��Ғa���c඾�yI�?����G��̡�<�,= �<=�i=�E�<�3;�����#�s�+˘�ϫ���   �   �#��g����~b��e)��L¼P���ؘ�<�*
=��?=r=U===�<�_��bu��^�L������\�+�d������ۿx9�p3�B]�6��R՝��.�������?��<���A�� ��dY����]�|�3�&��._ܿC��L�e���,����M��N��4L��Ժ�<��:=��R=j�<=�"=8�x< s���%ȼ��+�Ldd��$���   �   �R�����Ǘ��hp�� ��p���ߙ;l��<<^"=��?=��.= �<�n���ǲ��BH�����}�>�`��۟��׿���~	0�Y��H���P���!��|K���ؿ��H���(���n��T���Y�4�0��e��ؿ{u��Ƒa�2�`߶�jxI�����|C�����<�,=��<=�i=F�<@5;�����#�0s�9˘�߫���   �   �������Ƃ�ˏ��|�p����� �b�Ľ�<�n�<�c=���<p����|��2�;�bE���,���T��ї��~Ϳ�4�~@'�\EM�.�v��]��֍���ͮ����컮�z��+Z����v��M��'�֏��ο�M���U�q��X���=�U%�������A�<`a�<l��<�D�< ������X�t� h���!��r��q��   �   �4���ۂ���r�nU�Tx0�l2��5��x5W���� �,;��R<P	�; {��:Ù��M)�r��������(B�t0��5������2��V�;�z�_�ٳ��G�����2������W������o_�D�;����3����y���ۮB��N���N��E5*��9������@�;�oG<���:�����o[�݇���h���1�7}V���s�����   �   ^�ݾ��ؾ�˾����������x�p0;���ݱ�� ��A~�����μ ���@�������ݾ�z*��
v�O����ڿ�	�JG&��HD��Wa��Jz�X�������7x��b�y�B�`�
�C�x&��	��ۿd7��.^v���*�z޾�����`��4��h�Ҽ�z'�<=��j�#�o蟽�k���<��hz��^���O��ȗ˾�/پ�   �   �4,��(����UY�����}̾�l��k�i�[G�6�Ža�TW�v�
�$z�n����^�x������<Q����H�����쿲*���'���>���Q�j�^��c�<]^�<VQ��$>��I'�(���R�vy�����)HQ�*���繾z_�u���^|�B��4�	�lWd��Ƚ� ���k�Ge��54;`�������+�W�(��   �   6?|��lw��i��_T�I9����o���e��F�����0�g{۽'x����D�X�m�}&ɽ`�1�)���sW辎�*��Bm������ſ�/�������v,��6��C9��5���+��L�p:��q� ſ5O��J�l�z�*��>�ؚ��:�1���ɽLo���F��ǆ��@ݽ�1�B����j��4������:��U�Jj���w��   �   %������䢿����]����\��2������Ǿ�y����1�}^۽p���wt�	�������b�Q���>��<;�r�y�Y���O
����`���X�
� ��������h
����� �'W��E��#�x���:�����в��]b�����8��Nlu��=��G�ܽ��2�����Ⱦ��	���2���]�R?��2A���K��.���   �   �@��"�w�ؿTdƿQ�����Q%s�ws=��j��ž\r��("#�OaǽG���p��e�ǽL�#��ق�'�ž���#>��t�f��������ǿٿ�p��<���|ؿ�`ƿ�M������ s��o=��g��žHo��#��\ǽ8E��qq���ǽ��#�z܂��ž����&>��t���������ǿ�ٿlt��   �   �������j
�������Z�����H�x��:�f��oԲ��bb����5;��&lu�;����ܽ2�2������Ⱦ��	���2�y�]��<��G>���H���*���!����Vᢿ��������]�\�2������Ǿv����1��W۽Pl��nut��
�� ����b�X"���@��?;�:�y����������V���Z�
�B��   �   ~F9�V�5�� ,��N�><�uſaQ����l��*�|B�h���j�1�պɽ�o���F�iÆ�O9ݽ��1��~���e�����L}�8	:��U��Dj���w��9|��fw���i��ZT��D9���������_��K���Ҝ0�)s۽�r���D���m��(ɽ��1�D����Z���*��Em�����V�ſ�2￨�����@x,�6��   �   �c� `^��XQ��&>��K'����qU쿝{�������JQ����깾[}_�"����|�2����	�\Ld��Ƚ8� �u�k��`��o.;��������'���(�m0,�y�(�Z��gU�����w̾�g��h�i�.A�%�Žt�`�JO���
�hz�������^�����(��Y>Q�W��)����� ,�p�'���>�L�Q� �^��   �   ����y���y���`���C� &��	��ۿ�8���`v���*��|޾Y����b�k6����ҼHi'�-��$�#��ߟ�Qf���<�P`z��Y���I����˾)پ��ݾ��ؾ�˾􎵾a��� �x�);�������z ��~����|	μn���n����y�ݾD|*��v����|�ڿ�	��H&�NJD�Za� Mz�Ǣ���   �   ����u����,����q_���;�������G{������r�B�4Q��mP�� 7*�k;��̸��+�;��G<@��: u���`[�@~��&c�¡1�vuV�3�s�/��20��Pׂ��r�(fU�Dq0�\,��+��%W������0-;��R< *�;�w���Ù��N)�g������*B�A1��E�������~�;��_�״��4H��G���   �   �������{��
[���v�&�M�ܞ'�|���ο�N��"�U�R�����:=��&�����lD�<�g�<��<�S�<PP������t��_��%轻m�:l�j��,�����x����L�p�$w�� �a�TΑ<�z�<Rh= ��< �	}����;��E��B-���T�fҗ�NͿ\5�A'�4FM�V�v�e^�������ή��   �   �ٿ�$I��M)��)o�������Y���0��e���ؿ�u����a���#඾^yI������D��,��<�,=��<=Zm=O�<@�;\���̡#�6s�RƘ�����6M�������2_p��� �b����;���<tb"=��?=�.=H�<�l��qǲ��BH����}���`�ܟ�j�׿ ���	0�|Y�/I���P��"��L���   �   	Ͷ�ai��n���N����{�JAQ��o*�
���ѿ1����fY��Q�v�\�>�ߏ����E����<,vI=x`=�xK=�2=ܰ�< ��:P���B�B��d��xo�`gb�R�>���V�� 6;�@�<
|=�R=�g=�wP=��<��%��؟��;�s������\�W�Z�����Ͽz���Z)�^-P���z����*ƥ��c���   �   ���M����������v�NSM�0~'�ʀ��
ο�B��6mU�o���X���i:�
���h�G�4��<D�;=r�K=�s/=��<pu<�NA�f��Q�/��%꘽������ ���CK��4��(�#�`�6<X��<��6=f�R=��B=��<8(��b����7��r��ND�i�S�}����̿d��@�&�gL���u��֏��	���R���   �   ����ؕ���N���Ԇ���g�2B���������ÿ�m����I��� ���r�.����PgQ��@�<�=�d= ��<���:9ļ��R�������ѽV��������t�������ν�ٜ��J�$����U`;�e�<^�=<)=,b�<^3�ڳ����+��M��Gh��mH�����¿ë���h�ƪA���g��ن�Mo��]����   �   ����'���p���r�<aR���1�2)����೿(����7����
�����W�����o��:<�K�<P,�;0Jp�f�:�J�������.�#�`�F��0b�֬s�Ofy���r���`��D�8H!�9�󽊸��*�1���N�8[<��<�V<�
T��݄�7O�Ǫ��:c�6�6���h)����迬��6}1���R�v=s�����B^���   �   j��x�y�n8j���S�r9��g����Ͽ�z��i�o!�{�о�oz�z����r��H��p�����"��|��D��^���C.���h��'�������ھ���˾��Ͼ�˾Nɽ�P��Ė����e�RE+�]$�ڇ��H���Д��v%������&l�t��hx���ϾZ �(Sh�o.��A�Ͽ�/������9��^T��k�@`z��   �   ��U��XQ��XE��3��n��~��B࿩����>���E�}X��쭾��N�߽̑�PY��o޼D@ټ��B�so���z��Z����������~�3��4��:"�����C�����$���:����W�J��������;�,�̼XӼz T�ݽ��M�G����;`E��I��7���8�࿆��=�"�4�6;F���Q��   �   x\/���+�V�"�����$�R���D듿8�_��� �{�پ^b����#�@���V�L�*s&���i�5uǽ��#��x�5���c3�o����/�5xI���]��Rj��|n�3�i�Z�\�}&H��R.�3N����'���H�u�ub!�{�ý
5d���!���H��T�"�23����پq� �}D`�=r�������l�
��|��H�#�vu,��   �   ���Ng
�L����Lտ�-��������j�8�/������禾DHQ��������~NR���w���ƽjv$�;����=��"����(�	�Q��x�m���M嚿O��l���碿�,��ϟ���v��O�q'��l ����R�~�,�"��Ľ�Ht�4P��"���&�Q��a���|���0��Al�x���g��+�ֿ�Q����
�
��   �   n�ܿ'}ؿoKͿ)����饿�ߌ��]e��M2�<��;����q�������8Fm��m�ۋ�����2As�V@����ϒ3��g���� ��n+��HKο�ٿ!�ܿŀؿ�NͿR����쥿?⌿�ae�9Q2��������q�6�	����Gm���m�h������e;s�6<��N��<�3�}g����$(���GοOٿ�   �   -	���䢿})��
����v���O��m'��i �����
�~�ڲ"�eĽ�Ct��P�����o�����Q�>e��������0��El��z���j��k�ֿ^U����
���Ri
�N�D��,Oտ-0��ގ��"k��/�����ꦾLQ�P���;����LR���w�h�ƽ�q$�����9�����(���Q���x�����6⚿�K���   �   rwn��i�P�\��!H��N.��J���澑���K�u�d]!���ý�,d�$�!���H��R�"��5��u�پ�� ��G`�Mt������o����l��l�#��w,��^/� �+�j�"���^��&⿝���!퓿$�_��� ���پdd���#�L�����L��m&���i�cmǽ�#�s�x�E���9-龺��<�/�msI�z�]��Mj��   �   o6"�����?�i����羭��������W��������;��̼�SӼ�"T�xݽ��M�~I�����bE�LK��@������ �d?�0�4��=F�X�Q�(�U�8[Q��ZE���3�&p���&E�x���A@��>�E�Z���N��߽�PY�dh޼�0ټ��B��f���t�o�Z�X������X�<{�%���0��   �   6�Ͼ�˾rý��J�������e��>+�������h���u��2%����Z)l�4��,kx��Ͼ�[ �Uh��/��!�Ͽ�0�"��h�9��`T��k��bz�"���y��:j���S�9��h����Ͽ|��i��!�X�о8rz������r��C���\��@p"��o��;�����<.�\�h��"��&����Ծ���˾�   �   �]y�&�r���`���D��A!�3��i�����1� hN�p{<���<�%V<�
T�'߄��P�&���Se��6�6����*����迪��v~1�4�R�j?s������_��T���)���q���r��bR���1�*�C���᳿�(���7�����r��ί��X�o���:<�X�<�u�; p���:���������p�#�֟F��(b�D�s��   �   *{�@�������ν�ќ�p�J��t�� �`;�s�<p�=j,=�d�<�_3�*���M�+��N��i��nH�N����¿�����i���A�ʠg��چ�4p��U�������ǖ���O���Ն���g��2B�F�t���d�ÿn��]�I�k�������.������bQ��E�<.=�j=��<@Ѿ:� ļ�R�A���e�ѽB�����   �   �𞽢���]��6;K�&��p�#���6<���<��6=��R=�B=���<(��c��o�7��s���D� �S����3�̿¡���&��gL���u��֏�G
��6S��y���>N����?	��4�v��SM�t~'����(ο�B��|mU�����X��j:������|G�4��<|�;=��K=�w/=��<��<�2A��]��Q�?*��$嘽�   �   �xo�tgb�x�>����,W���6;�?�<�{=��R=Xg=xwP=���<��%�:ٟ�|�;�����#����W�}�����Ͽ���[)�z-P���z����4ƥ��c��	Ͷ�Yi��c���N��ֻ{�.AQ��o*����ʌѿ����fY��Q�3���>�P���h�E��<�vI=|x`=FyK=�2=x��<���:�O����&�B�Ζd��   �   �𞽳���n��F;K�(&����#���6< ��<�6=�R=��B=@��<@(�Bb��0�7��r�� D�$�S�L��W�̿4����&��fL�D�u�2֏�V	��0R��k���5M����m���v��RM��}'�j��G
οCB��zlU����W���h:�Q����tG����<f�;=
�K=�w/=p��<�<�2A�^��Q�J*��2嘽�   �   9{�L������ν�ќ�z�J�`t�� �`;�t�<J�=�-=�i�<�P3�'�����+��L���g��lH���=�¿���^h� �A�z�g�Lن�{n��p�������ޔ���M��Ԇ�t�g�1B���N�����ÿ�l��r�I���������.����� SQ��J�<� =�k=�<�ܾ:L ļ��R�D���q�ѽX���р��   �   �]y�@�r���`�ƃD��A!�<��a���T�1�peN�`�<���<�2V<h�S��ڄ��M������a�|�6�q���d(��������"|1�8�R��;s�����]��ɲ���&���o��$�r��_R�Z�1�0(�N��y߳�'��\�7�]�L	��!������@�o���:<(]�<���;�p�<�:�z�������x�#���F��(b�X�s��   �   D�Ͼ�˾�ý��J�������e��>+���u��,f��l�@�$�T���`l�P��>ex���Ͼ�X �<Qh�+-����Ͽ�.�v���9��\T�4k��]z������y� 6j���S��9�Ff����ϿAy���i��!���о;lz����\�r��6��0;���e"�dn�w;����<.�Y�h��"��.����Ծ�Ơ˾�   �   w6"�����?�p����羲��������W�����^�;�8�̼FӼ�T��ܽH�M��D��b�^E�BH��l�����*� <�.�4��8F�X�Q� �U�:VQ�,VE���3��l�}�n@࿞���0=����E��V�%ꭾ��N���߽�EY�Z޼�'ټ��B��e���t�N�Z�Q���ޒ��\�@{�,���0��   �   |wn��i�X�\��!H��N.��J���澊����u�]!�A�ýf(d�*�!���H��경��"��0����پ<� ��A`�_p��<���j�n�����4�#�8s,�(Z/���+�6�"����!�ѱ��3铿�_�� ���پ�_����#��}��|�L��f&���i��kǽ��#�4�x�5���2-龺��?�/�psI���]��Mj��   �   3	���䢿�)������v���O��m'��i �������~�D�"�^Ľ�<t�~�O�qO�����Q��^���x���0�V>l��u��e���ֿKN�����
�v��Fe
�.J�?���Hտ�*��?�����j��/�6���!䦾CQ��������AR���w�@�ƽ�p$������8�����(���Q���x�����9⚿�K���   �   s�ܿ+}ؿtKͿ.����饿�ߌ��]e��M2�6����v�q�
������<m�`�m�䀲�����5s�Z8������3�cg��썿���$��RDο�ٿ��ܿ�yؿ�GͿ��祿:݌�LYe�_J2�n�������q�.��
���9m���m�O�������:s�<��B��7�3�|g����'(���GοTٿ�   �   ���Pg
� L���� Lտ�-��������j�4�/����v禾�GQ����������AR���w��ƽ�l$�n����4��;���(�=�Q���x�Ā��3ߚ��H�����Yᢿo&��1�����v�Y�O��i'��f � �����~�c�"��Ľ�5t�\�O��s���R�Q��a���|��ۭ0��Al�x���g��-�ֿ�Q�����
��   �   x\/���+�X�"�����
$�T���E듿6�_��� �V�پb����#�ۀ����L�Zc&���i�eǽ��#�4�x�����`'�1���/��nI�o�]�@Hj�rn���i�4�\�!H��J.�G���澠�����u�uW!�m�ýPd���!��H��첽>�"��2����پf� �wD`�;r�������l�
��|��H�#�xu,��   �   ��U��XQ��XE��3��n��~��B࿫����>���E�qX��쭾��N��߽HY�8V޼�ټ.�B�^��o�+�Z���_����꾙w�/��s,�-2"�����;�������~�� ����W�ֺ�fꮽ8x;�ؘ̼�>Ӽ�T�M�ܽ��M��F����3`E��I��6���7�࿄��=�"�4�8;F���Q��   �   j��z�y�n8j���S�t9��g�� �Ͽ�z��i�h!�V�о\oz�v��8�r�,5��p���F"��b�k3��Iu�6.�B�h����ϫ���ξ���˾��ϾW˾����OE��3�����e��7+����v��8L���G� �$�h���& l�h��wgx�t�ϾZ �#Sh�n.��?�Ͽ�/������9��^T��k�@`z��   �   ����'���p�� �r�>aR���1�4)����೿(����7���
��Ȋ������o�(�:<�g�<p��;��o���:�J���������#���F�� b�כs�Uy���r���`�D|D�;!���󽵥����1�h4N�(�<���<�BV<��S�\ۄ�|N�����c�6�4���g)����迪��4}1���R�v=s�����C^���   �   ����ؕ���N���Ԇ���g�2B���������ÿ�m����I��������.����0UQ��M�<�#=�p= �<��:h	ļ6�R�=���]�ѽr���{��u��������ν\ɜ��J�\����a;|��<4�=2=o�<�K3�_�����+��M��>h��mH�����¿ë���h�ƪA���g��ن�Mo��^����   �   ���M����������v�PSM�.~'�ʀ��
ο�B��6mU�l���X���i:�U���hwG����<��;=B�K=4{/=��<h�<�A�rV�
�P��%��>����랽�������T2K����p�#���6<��<�6=&�R=�B=X �<�(�b��T�7��r��KD�h�S�}����̿d��>�&�gL���u��֏��	���R���   �   �@���`���|��������b� Q>���d��E��R�����E� ���^��nR&�j&���j��<=��`=8[v=2�b=�%3=8��<p(<��黸͸���J�,�F�5�z)�K����9��ȧW<���<j@=<�o=\��=��m=N3 = H�:��z���!�&���Z��*aC�� ���V��������=���a�3J��f]��\���   �   {����ƚ�3���̀��S^���:�Bv��=�����%*��IB�����^���"� Ձ�� ��U=�'T=�%c=^�H=��=���<�;غlʪ�|*�F�Q�^�s�~A~��3p���J�~��|����ٮ:�Z�<��=��U=�"p=a=|f=��:��t��R���d��l�?�����7���%�W���9�j�]������'���̚��   �   ������v���D�q�b�Q�f1�B��J4�G���g⃿�e7��ﾸ���=��q� �%�,��<ڬ,=E(=���<x�-<�S��+�B���xҮ�I>ҽ1�轓z���t~ν�����v��������d<�l=�X5=u9=�= �.:��b�E{�r����hz5�e���F��/�翶��}0��sQ���q���������   �   ��(���j�r�>�Z�� ?��S"�:�6qֿw�����p�)�&��ؾuπ�����~V��l��D�<�E�<��<�R���툽	�ҽ&��T�-�h�F���V���[�T�U�7�D���*�e�	�KX˽�L���L𼀎d�䎞<�g�<H*�< ����I�0h�Z�}��վ�K%��Qo�ƣ�*�տ���B"�e?���[�R�s�����   �    f��a�h�S�8@���(� 9�����������S�~���>��-]�z}彪�9�H���; �9�Ϫ��@_�Z~Ƚ[\��WM�r���Uf��GЪ�5u���1��櫵��[��w����}�C�H����C���HP�tƏ�`#N;��< M���'/���߽Z�#���o���S��T��d��E��j��*�)�NA���T�~�a��   �   j$B��5>�j�3�~$������4�Ϳ#o��Rx�?,3�(���$��p5��	���O"��ŀ��Ix�D������D���j@�Tu��#���x�ҾK���$�������kl�l�����Ͼsĩ�0ӂ�\�;��,��Qʋ����N�`R\�Ƶ��b3��0��j�%�2�`fx��ã��Vο����$
��.%���4���>��   �   be ��R���̗�)�8ϿĪ�K↿�.K�R��8þ�t�f��l)��4C��^�l�1�G�����(�[� ����Ѿԑ��T�7���I��2U�0�X��xT� 7H�BR5��~������ξ�Q��CJW�#
��Y���(��_׼L�ꕐ����=t��8þ�^���K���֫���пi����	������   �   �b��������W�ܿ�QÿT����T���xU�I
��9ྶq��8�6�4�Ͻ�c�L�n�=��ꣽ��Yic��z��٤�&�=�>�i�b��6����� N���Ǘ��͔�W������NK`�rY<�j#���T*����_��x�W5��V}8��l�Hqa�z�Ͻp+7�����j� �@W�dz��y���ſU�޿�^�t����   �   &@ʿ�kƿ4���t䫿t��G���0P�'.!������h:T��T��6���Z3��3����q �wJV�&���i+�X�"�&]R���������ca���5��&ǿ�Cʿoƿ_��_竿�v��bI���4P�/1!����a�� ?T��Z��o����3���3����n �%EV�]���O&��"�YR�(�����W^��|2���ǿ�   �   �ė��ʔ�����l���F`��U<�) ����a&���_��t�^0��~x8�dl��ua�Z�Ͻ|/7����o�� ��W��|�����ſ��޿eb�3����d�����j�𿆼ܿ�Tÿȇ���V���{U����=�at����6��Ͻ��c�����=�壽K���bc�cv��B�龫��>���b�B4��%���%K���   �   +�X��sT�Y2H��M5�8{�h����ξtM���CW�x�	��S��^�(��X׼6	���������At�+<þ�`���K�؊���ث�a�п�����	������rg ��T���z���:Ͽ0ƪ�䆿T1K�S��;þ��t����G+���B��T�(�1������0�[������Ѿl���P�� 7��I�.U��   �   ���h�Ǒ�`����Ͼo���ς�յ;��"��Ë���N��J\������B3��2���!�q�2�aix�sţ�Yο������j0%���4���>��&B��7>�b�3�:$� �a���G�Ϳ�p���Tx�:.3����&���5���P"�ܾ���-x�������9���c@��p��ڑ��U�Ҿi���j�����   �   �+��8���vV��7r���}���H�����9���9P�ܰ����N;�<�F��,*/��߽�Z�S������S�V���e��a�����)�A���T���a�Tf�2a�h�S��@�>�(�H:����.�������x�S�Ƥ�v@��D]��彄�9�@�� :�; #9h����0_��sȽ�U��OM�����Fa���ʪ�uo���   �   ��[��yU�܇D�H�*�t�	�$N˽}D���1��a����<xq�<H/�< ����I��i��}�شվM%��So�Cǣ���տ���&C"�vf?���[�B�s����Ä�0���B�r���Z�6"?��T"��rrֿn����p�1�&�MؾPЀ�����V��`����<�Q�< �<��������䈽Y�ҽ��e�-���F���V��   �   �pｃw�^uν1���T�v����p��`�d<Fs=�]5=�w9=@=�v.:d�b�x|�r��]�x{5����*��L��d��~0��tQ���q����d������ݞ��-���t�q�P�Q�1����#5�솳��⃿Af7���D���ʉ��q� r%�$��<°,=�J(=p�<p�-<h^S�n������ɮ��4ҽzw��   �   &8~��*p�F�J����İ�����:�d�<��=��U=�$p=<a=�f=��:��t����R���e���?�o���78��_&� X�b�9��]����
(��q͚���Uǚ�3���̀��S^�&�:��v��=����V*���B��������"�Ձ����.W=�)T=�(c=�H=R�=䠒<@i׺|���4"�X�Q��s��   �   D�5��)�FK�h���;����W<���< @=��o=-��=t�m=�2 =�1�:��z�<�!�g���ZZ��`aC�!���V��0�����=���a�@J��q]��\���@���`���|��������b��P>����d���D��1�����E�����^��R&��%���Q���=(�`=�[v=��b=�%3=��<�(<��黐͸����4�,��   �   H8~��*p�h�J����̰��@��:�d�<�=��U= %p=�a=�g=@*�:��t����Q��Gd��*�?�ӷ��k7��_%�\W���9���]�j���:'���̚����mƚ��2��3̀��R^�H�:��u��<��M���)���B���������~"��Ӂ�@��xX=�*T=.)c=\�H=��=��<@g׺h���B"�p�Q�2�s��   �   �p｝w�|uνG���f�v����H��@�d<�s=b^5=Xy9=�= Z/:��b�Nz�����쾼y5�챂����a��2�8}0�sQ�f�q�&��ý�����9��������q�F�Q��1����'3�Z����ჿzd7�ﾗ�������q��6%����<P�,=~K(=��< �-<�]S�T������ɮ�5ҽ�w��   �   ¾[��yU��D�V�*�}�	�'N˽rD��P1��a�(��<@u�<�5�< ߥ���I��f�M�}�x�վ�J%�_Po�$ţ���տ4��A"��c?�p�[�~�s�����������t�r���Z��?��R"�N��oֿ@�����p���&��ؾ�̀�����wV�7��L��<V�<�"�<���@��_䈽F�ҽ��j�-���F�ϰV��   �    ,��D����V��@r��(�}���H�����9��N9P�X���`�N;�<p��� /���߽b	Z�M���"��S��S���b��m��F��ƚ)�� A��T�H�a���e�� a�R�S�f@�H�(��7����瑾����y�S�ء�`<���]�Bx���9�p���Y�; �%9H����/_��sȽ�U��OM�����Ja���ʪ��o���   �   ���h�͑�l����Ͼv���ς�ŵ;��"��^�����N�01\�����鶽d3��.����+�2��cx������Tοu������,%���4���>�."B��3>�b�3��$��-����Ϳ=m���Nx��)3����["����4����E"�d���x�N��7���A9���c@��p��ԑ��R�Ҿl���m�����   �   2�X��sT�_2H�N5�<{�m����ξmM���CW�#�	�YR��L}(�L׼��א�����B9t��5þ�\���K�5���pԫ��пs��J�	�$�����Tc ��P�����	�I5Ͽ����`����+K���E5þ�t����N#��$8�<G�ƚ1��������[�v����Ѿh���P�� 7���I�.U��   �   �ė��ʔ�����o���F`��U<�, ����O&����_�<t�v.��Nr8��b��fa�"zϽB'7� ���f�t ��W�Sx�����ſ#�޿P[������`�>���e���ܿ�Nÿ�����R���tU�g��5�un��d�6�ӫϽt�c�|�r�=�㣽����bc�Cv��/�龤��>���b�B4��'���)K���   �   +@ʿ�kƿ7���w䫿t��"G���0P�'.!�������9T��R��p����3�f�3����2j ��?V�є���!��"�KUR�♁�6�f[��M/��gǿ�<ʿ[hƿ����q᫿Vq���D���,P��*!�������4T��K��?���3���3���(m ��DV�3���6&�	�"�YR�'�����X^��~2���ǿ�   �   �b��������Z�ܿ�QÿV����T���xU�G
��9྅q����6�ְϽ2�c�r���=�$ޣ�����\c�Or�����`���>��b��1��X���5H�������ǔ��������B`�gQ<���*�� "��n�_��o��(���k8��`�\ia��}Ͻ�*7�����j� �8W�bz��x���ſW�޿�^�w����   �   de ��R���Η�,�8ϿĪ�M↿�.K�L��8þ��t�o��6&��F9� A�(�1�a�z���[�9�����Ѿ(��M�X�6�H�I�)U�,�X��nT��-H��I5�Qw���
�ξ�H���<W� �	� K���s(�4B׼@����������<t��8þ�^���K�숇��֫���пh����	������   �   j$B��5>�l�3��$������7�Ϳ%o��	Rx�<,3���$���5�\���G"�䭀��x����󦒽E/��0]@��l��Ȍ��e�Ҿ�y��Æ�<��(���d�������Ͼ;����ʂ�ʮ;����h���h��x|N�H#\�­��붽�3�x0��H��2�Yfx��ã��Vο����$
��.%���4���>��   �    f��a�j�S�:@���(� 9�����������S�x���>���]��{彘�9�����x�; �,9����� _��iȽ�O�xHM���\\��mŪ��i��/&������
Q��:m��8|}�:�H����}/��<)P�\����@O;�,<����!/���߽jZ�����c���S��T��
d��D��h��*�)�NA���T�~�a��   �   ��(���j�r�>�Z�� ?��S"�<�8qֿy�����p�&�&��ؾEπ�G��\zV� 8�� ��<�_�<�1�<�9������ۈ��ҽ�����-���F� �V�̶[��qU�s�D�p�*�W�	��C˽�;��`��^�<��<0��<�<�<@�����I��g��}�вվ�K%��Qo�ƣ�(�տ���B"�e?���[�R�s�����   �   ������v���F�q�b�Q�h1�D��M4�I���h⃿�e7��ﾛ���҈�Bq�`?%�`��<D�,=4P(=��<�.<p3S�����������+ҽ�m�g��m�:lν�����v����XX�8�d<{=�c5=R}9=�=��/:2�b��z�S����ez5�d���E��-�翶��}0��sQ���q���������   �   |����ƚ�3���̀��S^���:�Bv��=�����%*��JB�����Q���"�zԁ� ���X=,T=:+c=`�H=��=��<��ֺ|���\�ГQ��s��.~��!p�~�J�z�� ����g�:�o�<��=��U=�'p=a=ri=�D�:Z�t���R���d��i�?� ����7���%�W���9�j�]������'���̚��   �   ���{���Tm|�,c��E�J�'��V
��:ݿ�	���+y�4�,���߾6˄����;� U1<�?7=Z}=/F�=B�~=�T=�= d�<���;�m��8���Xhʼ�ټ����`ف��T���
(<0�<�u.=��i=��=�n�=�ǉ=ZSM=h�<��#��]��4��̈́۾B�)���u�A��>�ڿ�%	�Ԃ&���D�
�b��;|�����   �   �������,w���^�6B�*�$�\�a�ٿh���t��W)��C۾�ց��2�$5��+0<VJ1=*�q=�D=�g=z6=<�<��5< <ƻ����2���$��j-�������������{����<N�	=6�K=��}=1��=I�=�G=Lƃ<J~�:��\�|�%׾d�&���q�OE��4u׿j����#��kA�>^��w����   �   8r}���w�\kh�x�Q���7��h��S���ο펞���g����}ξ��r�ֿ��J1$�0�(<�=
kN=2[J=��=T@�< �s:,���74�P���������z庽�g���x���4v�<�"����pD�;��<��5=<`=6�c=�3=�|<,�Z�齸ol�@wʾu��`e����94Ϳ�� ����t�7��
R��h��x��   �   ��d�4
`�οR��L?��B(����y���彿u/��%S�.��Ơ��.wX���ֽ��X5<��<�=2�<�<(��0�A�ࢽI�b��-$��2��^6��0�@?!���	�eVٽ�5����+��8=���e<��=X%=8y=x�]<�b��?ͽDGS�D���yL��ZQ�'A������N�����(���?��]S��t`��   �   �]H��GD�J9��)��X�������ӿ�m��B"��+9�;��<���7�CҲ�U���;���<6Q< Ȼ��A���:���eN*�*�X��0���p��K����۞�@���������}�\\S�jU$�ժ�	���P��������8�<���<� <�'ļ���� �3�h靾q&��J+8��t��=��0�ӿ�> �b�|�)��&:���D��   �   
�*��~'�n���-��� �SQܿr۵������Y����Ҿe��|'�希��5�� ��� �T��0��v�R�_�ȽJ���`��1��﴾�Ҿ�n꾲=��%������5��Ͼ����	���tIZ�0��TM����>��e��I;��;$���䆽$}�
3��hѾ���Y��V��[���s�ݿ���J:����0(��   �   ��[�� �I;�]�ֿqM��������l�h-1����vŦ�N�L������Q�������H���ԼL�r�����6��V���C��L��k
��{��/�mL:�ؓ=�݂9�!�.����AX��,�#w�����\91��*ٽ�b�������"��zHJ�-�ݽQ�K�J���������1��n�H����޸���ؿ0O����<���   �   ���1�Bvտnÿ$��������4o��F:���	�rT���az��/�yE��.a��������Z�o��,���=�n���Fɾ���c;&�WvF���b�V�x�Ae��B���d߂��w��p`�u�C��#������žR���?+9�<_ܽ��e��cټ�=��H��&����{�������
�h�;�W�q�UD��|j���Eſd�ֿo��   �   -����x���������7(����`��~5�<���_˾Jڊ�/�L#ǽʈI���Ҽ� ռ�[M�ކʽR�1�(�Tξ<x���7�7�c���������K��{+��@����{��q��+����*����`�T�5����c˾P݊�M/��(ǽ��I�`�Ҽ@�Լ�TM���ʽ��1�̾���ξOu�>�7��c�7�������H��n(���   �   �����܂��	w�Il`�b�C���#�˥��žΗ��$&9�&Xܽ��e��Zټl=��L���������{�b����
��<�X�q��F��/m���Hſ� ׿��J��%5�^yտ�pÿ����Դ��A8o��I:�&�	��W���fz��2��H���c�����$����o��$�V�=�>j���Aɾ����7&�rF��b�2�x��b���   �   [�=�{~9��|.�ݕ��T�5'�kr�������31��"ٽn�b��빼 	�4$��XMJ�	�ݽ8�K�.æ�����W�1��n�]���4ḿ��ؿOR��>������\��"�D>� �ֿ�O��l�����l��/1�`���Ǧ���L�o��b�Q�������H�0�Լh�r�ǫ���6��R���>��F�yh
��w���/��G:��   �   ���:��w/�'�ϾU�������&BZ�_��qD����>�(�d� ZI;`;x����憽��5��Y!Ѿ�����Y�;X��g���ۤݿ$���;�L��(���*���'���^/�ܟ ��SܿOݵ�W��s�Y����hҾ�f��z)�Ѻ���6�� 8���bS�����R��yȽ��V�`�-���鴾��Ҿh��6���   �   �֞�5���8���L�}��TS��N$����hХ�������E�<���<�<X,ļ����z�3�V띾?)��6-8�;w�;?���ӿ�? ����)�\(:�^�D�f_H�fID��K9�f)��Y�����V�ӿo��T#���,9�e=��������7�(Բ��V传�;��< TQ<��ǻ�{����������G*�&�X�X,��l��3����   �   wW6��0��8!���	��Kٽ�,����+�H=��f<��=�%=�{=��]<|g�}Bͽ�IS������M�&\Q�7B��
��EP�ܤ��(��?�_S�zv`���d��`�L�R� N?��C(�г�����潿S0��j&S�������xX�V�ֽ���:<���<v�=XA�< �< e��"�A��֢�=��6��l&$��2��   �   �ܺ��^��kp���%v� �"�D���P��;+�<��5=L@`=��c=F�3=P|<P���ql��xʾd���e�a��65Ϳ&� �z��V�7��R�H�h�Nx��s}�F�w�~lh�n�Q���7�.i�hT�T�ο������g�9��Nξ��r������1$���(<T�=�nN=0`J=n�=Q�< `v:���H)4�SH��E������   �   �b-����t�������@��<��	=��K=.�}=��=��=G=Ń<���;����|��%׾��&�v�q��E���u׿���L�#�dlA��>^�~w�x�������-w�<�^��B�t�$�����ٿ���Y�t�X)�D۾�ց��2��5��.0<�K1=
�q=VG=<�g=�6=`�<0�5<pƻ����<�\�$��   �    �ټė���ف�PV���	(<��<�u.=Z�i=���=�n�=bǉ=�RM= �<��#�$^�5���۾q�)���u�b��c�ڿ�%	��&���D� �b��;|�������v���Fm|�c��E�4�'��V
��:ݿc	��R+y��,�I�߾�ʄ�ȟ��;��W1<b@7=xZ}=]F�=��~=*T=V�=�d�<���;�l������<hʼ�   �   �b-��������䢒� ��<��	=��K=j�}=Q��=-�=.G=lȃ<B}��9����|��$׾*�&�^�q�E���t׿6����#��kA��=^�4w����C��e��8,w��^��B���$���Ńٿ���8�t�@W)��B۾ց��1�05�60<�L1=��q=�G=��g=�6=��<��5<ƻ����D�f�$��   �   �ܺ�_��~p���%v�6�"�\������;P+�<�5= A`=&�c=N�3= |<R���齎nl�hvʾ٥��e����3Ϳ� �,����7��	R��h��x��p}���w�jh�b�Q���7��g�NS���ο���^�g����ξ��r�Ӽ��x,$��)<��=pN=$aJ=�=�Q�<�pv:����<)4�PH��Q������   �   �W6�,�0��8!���	��Kٽ�,����+�X=��f<��=�%=T~=��]<�Y�"=ͽoES������K�:YQ�P@���
��TM����(�z�?�\S�"s`��d�~`�<�R�xK?��A(�������使^.��j#S����򞹾�tX���ֽH��M<ܖ�<��= D�<x�<�c����A�p֢�,��5��p&$��2��   �   �֞�?���B���[�}��TS��N$����J|��� a���I�<���<h<�ļ.񪽣�3��睾"$���)8��r�V<����ӿ�= �.��)�%:���D��[H��ED�TH9�n)�@W�M�����ӿ)l��� ��)9�08�����7��Ͳ�E�`?�;���<^Q<@�ǻ�z���������nG*�"�X�X,��l��9����   �   *���C���/�1�Ͼ_�������&BZ�P��#D��^�>�`�d���I;�_;H����߆�sz�01���Ѿ-����Y�U������=�ݿt���8���b(�,�*�}'����N,�*� ��Nܿaٵ����[�Y�����Ҿ�b��&$������#���p���]R�t��d�R�+yȽ���8�`�
-���鴾��Ҿh��6���   �   _�=�~9��|.����T�<'�or�������31��!ٽ:�b��乼������X?J�}�ݽz�K��������;�1�un�^���yܸ��ؿ3L����|��
�BY�>�18򿔌ֿ�J��l���5�l��*1�� ��`¦�ƊL�����Q�H���@�H��Լ��r��⽆�6��R���>���E�xh
��w���/��G:��   �   �����܂��	w�Ol`�f�C���#�̥��ž�����%9�"Wܽ
�e�xOټ�+��~>�
Ᵹf��l�{����A�
�g�;���q�B���g���BſD�ֿ'⿓�忌.�sտkÿy���G����0o�JC:�G�	��P��,\z�.+��>���U� 橼 �� �o�i#���=�j���Aɾ����7&�	rF��b�5�x��b���   �   0����x���������9(����`��~5�=���_˾.ڊ��/��!ǽ��I�pvҼ�Լ�IM��yʽ�1������ξ�r���7�Ґc�ڷ��+���E��j%����u�����׈���%��b�`�_{5�Q��*[˾�֊��
/�]ǽ(|I�DpҼ\�ԼOM��~ʽ�1������ξFu�7�7��c�6�������H��o(���   �   ���1�Gvտnÿ(��������4o��F:���	�]T���az��.�KC��0Z�0橼Ĵ�\�o�p�؇=��f��*=ɾ���!4&��mF�t�b�+�x��_��ߏ��ڂ��w��g`�&�C���#����&�ž쓌�/ 9�Oܽz�e��Cټ�'���@�a흽d���{�s�����
�_�;�S�q�RD��{j���Eſe�ֿq��   �   ��[�� �N;�`�ֿuM��������l�g-1����VŦ�ȎL����*�Q�p���8�H�d�Լ��r������6��N��:��7@�e
��s���/��C:��=�z9��x.����nQ�;!�rm������T-1��ٽD�b��ӹ����0��\BJ�5�ݽ��K����������1��n�E����޸���ؿ/O����<���   �   
�*��~'�p���-��� �UQܿt۵������Y����Ҿ�d���&�����l'���?�� Q���x�R�KpȽ����`��(��Z䴾��Ҿ�a��/��&���Z����(��Ͼ��������n:Z����:���>���d���I;��;t����ᆽ]|��2��DѾ��إY��V��X���q�ݿ���J:����2(��   �   �]H��GD�J9��)��X�������ӿ�m��D"��+9�;���X�7��в�J传C�;X��<�wQ< dǻVm����������@*�d�X��'��Bg��+����ў�*���k���o�}��LS�H$����捽���� ���X�<0��<�!<�ļ��k�3�<靾X&��C+8��t��=��/�ӿ�> �b�|�)��&:���D��   �   ��d�4
`�пR��L?��B(����|���彿w/��%S�,�������vX���ֽ��PM< ��<��=�Q�<��<�K����A�P͢����0���$��2�rP6�4�0� 2!���	��@ٽ##���}+�h�<��8f<Z=�%=��=@�]<�Z�>ͽ�FS�&���oL�zZQ�%A������N�����(���?��]S��t`��   �   8r}���w�Zkh�z�Q���7��h��S���ο���g����rξʧr�����.$��
)<��=�rN=TeJ=��=a�< �x:����4��@��0������Ժ�tV��Ah���v�z�"�pފ�@��;�;�<��5=�E`=��c=��3=8|<�����{ol�.wʾp��[e����84Ϳ�� ����r�7��
R��h��x��   �   �������,w���^�4B�,�$�\�c�ٿi���t��W)��C۾�ց�b2��5��30<M1=��q=�I=@�g=x6=t%�<�5<@�Ż������H�$�DZ-�z����������� ���<��	=��K=̭}=���=!�=|G=ʃ<�|��9��A�|��$׾`�&���q�PE��3u׿j����#��kA� >^��w����   �   8d�2f_��9R�r�>���'�\P�x3��H��i����TR��C�Z����T��'˽غȼ<�<�[=�`�=���=��=u=^C=ī=�ڪ<�< 6x9਻p�һ@^`�@bl;�f<���<N�)=^�d=�Ȍ=�=N��=�w�=d��=.[=8���9���L�����܇�.O��Ꮏ�T��V:��m��-'��v>��R�Xd_��   �   ,�_�P[�">N��a;�^�$�����;�N������lN�?m��n��,�O�M(Ž������<��V=�m�=�2�=�܂=��Z=R#=�K�<��&< h1�p�N�䡘�����tX���T���;�r�<�=j�D=�F=���=�E�=�B�=�{{=\�=ةt�Rz���EG�Gί���
�uK��q���D���x��$�g$�� ;�6N�@[��   �   �S�\�N���B���1�������m�ݿ ���骆�sC��2�����$A�����轟�h�<�'G=jjp=ʡl=��G=�-=�}�<�zs�`6{!�hV�0�v�£���o�b=H�^��`��@`n;�V�<0�.=�Gl=���=xG�=��i=ʣ=�A�����Ie9����N��-�@�xW��5U��ņܿ>��i���1�d/C�P�N��   �   �L@�t�<�d&2���"�����h����˿y����
v�b1����G����*�������h�`I�<�{*=p3;=�S=��< p?9�Լn|[�ҟ��Oս����@	�Ly�0(�O��mʽt\���=�t;����<�;�<l2@=z�\=�J=��<�������#��5��\���/��Qt�=��lL˿�T��F��#�6�2���<��   �   ��)��&����Ă�� �Bۿ���@���dX�N��}jоjj���\�(�t��{�D��<���<ܻ�<�2!<<����=L�v��XP�,++��N�j�6`{��H�� 0y��e��H�@$� ����ͣ�^*��(��3�<~
=JS=��<`�.�D�^�M	�^~�/ξX��I�W�W���"����ۿ#� �N;����'��   �   ���A�`�������ܿ����������s�r�6����0��P�Q���޽�2���r��Mp<(St< �߹�S�` ����D2�֢m�5���^>���J����;	�Ѿ�̾�ݾ�6奄^����>e�ܿ)�jg⽞�|�l������;��<<��<��s:$�!���׽��N�6���`�u�6���t�檛�u����޿���������   �   ���3ￅ��n�Ͽ΁��k7���F��TG�c���Ͼ*���wx�L�����开҉��h�;�Qڻ��������� �U����������P��y����T���*�,��L ��X�u{��]���D�M����1��L�������<��;��м!���Hs����Ͼp��O�H����4���v9��q`ѿe%�6���   �   ��Ŀ����'����Ѧ��ܒ�Ɗx�tI���\侵����bF�$:߽��M�PIv���̺80	����ſ��Z�N�f�����+ܾ��
�Q�&�N?��(R��!^��a�e$]�	WP��<�'�#��;�R�׾+��� `�0�����,���p�� �9؟d���L���4(H��8���s�Wq�p�K�}{�ކ��#w��r鷿�����   �   ky��Pl���/������ �`���<�����	����*m]�Fq��$����Ѽ 尻����kܼ֮�����(�a�����������?���c�����vQ��G��|���n��42��ք���`�b�<����2羖���\r]��t��)����Ѽ�ﰻ ���h_ܼ{���ļ�n�a�(����������?�L�c�8�N���
���   �   g�a��]��RP��<���#��8�Z}׾9���`�ĵ�؋���y��0 9�98�d���L�/���,H�:<���w�&t���K�*�{�8����y��=췿s����Ŀj���ܔ��Ԧ�ߒ���x�BwI�|��O侜����fF�|?߽��M�0Rv���̺�	����󸣽6U���f�Z��=&ܾ��
���&�.	?��$R��^��   �   s��'�������Rᾊv��P���؟M��������P���@Q�x�<��;��мF����v����Ͼ���E�H�଀�Y����;��%cѿO(�?����/�V���Ͽ���k9��J�>WG�w���ϾT���T{���������Ɖ����;@ڻ���������B�U�X�����������������   �   �Ѿ(�̾ؾ�$ꩾ滏�F7e���)�e]�@�|�Ā�� �;L�<���< Ks:ث!���׽��N�� ���b���6�}�t���������c"޿=���8��B��:�pC����\���_�ܿ����U���{�s���6�v���2��)�Q�.�޽:2�@�r��Wp<�ht< 5۹�:���R��B>2�Кm�����"9���D����;�   �   2D��y'y���e���H��$�����,ģ�
O*�P���D�<փ
=�V=��<@�.��^�2O	��~�q1ξ���s�W����%$����ۿ@� ��<�`��� '�h�)�r�&�������� ��Cۿ���+B���fX����tlо�k���^�n�t��~����<���<���<X!<Hᅼ�-L�!l��mJ�M$+��wN��j�{W{��   �   8s�:"��C�tcʽNS����<�D!�� (<�K�<h8@=h�\=$�J=8��<��W�����#�7��^�h�/��St�->���M˿�V��<��#�p�2��<�RN@���<��'2���"����Aj����˿r���Lv�&c1�H��X���m�*������h��K�<F~*=8;=�Z=�Ʒ< �J9\}Լ�k[�N����սZ���B	��   �   ���*�o�V/H�z���I����n;Xg�<��.=�Ll=�=�H�=��i=��=A������f9�����B�@�+X��V��̇ܿڄ��i�\�1�T0C�R�N��S�T�N���B�T�1�4��R��?�ݿɬ��l���3C�3�8���%A�����������<x)G=zmp=$�l=N�G=5=p��< �r�dֹ��m!�qV�:�v��   �   4���XJ��@:��B;\}�<��=R�D=�I=˼�=�F�=!C�=
|{=֛=x�t��{���FG��ί��
��uK�cr��SE��ly�J%��g$�$!;��6N��[���_��[��>N��a;���$����!<鿕������lN�qm�1o��n�O�~(Ž������<�V=�n�=�3�=ނ=� [=�#=V�<��&<�1���N�x����   �   `�һ _`� al;��f<(��<"�)=�d=hȌ=��=(��=lw�='��=�Z=ܑ�����ZL�ꇳ���A.O��Ꮏ�T��y:�n��-'��v>��R�^d_�8d�,f_��9R�b�>���'�JP�U3��H��K���mTR�eC��Y����T�@'˽(�ȼh=�<��[=�`�=ݬ�=,�=hu=�C=�=�ڪ<��< Lx9Pߨ��   �   L���|J��x:�`B;L}�<��=^�D=�I=伕=�F�=eC�=�|{=P�=@�t��y��ZEG�ί�P�
��tK��q���D��xx翴$��f$�N ;��5N��[���_��
[��=N�a;���$�N��!;����F���kN��l�/n���O��&Ž�ｼ(�<0�V=�n�=�3�=Kނ=� [=�#=\V�<X�&<  1���N������   �   ���<�o�r/H�����I�� �n;lg�<��.=Ml=È=4I�=��i=\�=pA�6���Bd9�:�����p�@��V���T����ܿ���|h�ʘ1��.C�Z�N��S�V�N���B���1�֙�,��Y�ݿ;���1���SC��1�L��#A����@���D�<�+G=�np=&�l=�G=�5=,��<��r�ֹ��m!�qV�@�v��   �   >s�D"��C�cʽWS����<� !��()<�L�<N9@=��\=��J=(��<��ﻫ���&�#�q4��rZ���/�Pt�<��BK˿�S��n��#��2���<��K@�"�<�&%2���"����g���˿J����v��`1�~����΂*�.󙽈�h�pT�<>�*=":;=�[=�ȷ< vK9H|Լ�k[�3����սU���C	��   �   8D���'y���e���H��$�����'ģ��N*�8���F�<��
=|Y=��< l.���^�K	�~�-ξ���v�W�-��!����ۿ� � :�����'�l�)���&�,�����x �@ۿ�񴿗?���bX�����gо�h��IZ�̽t�h_���<���<���<�^!<߅��,L��k��PJ�@$+��wN��j�W{��   �   
�Ѿ.�̾!ؾ�+ꩾ컏�E7e���)�E]⽠�|��~��+�;��<ܣ�<�Lu:��!���׽R�N����^_�m�6��t�I��������޿���\��:��"�j@����#�����ܿ����������s��6�"���-��a�Q���޽��1� dr��np<xxt< �ٹX7�v�����>2���m�����9���D����;�   �   w��$'�������Rᾏv��Q���ʟM�x��h���T��� �ﺐ�<�^;D�м"��o�;톾t�ϾZ����H�f���7���'7���]ѿ�"�:����.	￠�⿿�Ͽ`��I5��C��QG���Ͼ򆾈t�N���8�开������;0�ٻ,�� ��D���U�B��v��������������   �   j�a��]��RP��<���#��8�\}׾5����`�����@s���Ÿ� !�9�}d�x�L�}���#H��5��}o��n�7�K�0y{������t���淿�����Ŀ����b���	Ϧ��ڒ���x��pI�����V����]F��2߽�}M� !v���˺(	��������T�|�f�?��'&ܾ��
���&�+	?��$R��^��   �   ly��Sl���/�������`���<�����	������l]��p��#��p�ѼЫ��б���KܼP��������a��������
��]�?�-�c��끿eL������v���i��--��0�����`�,�<�������&g]��l����(�Ѽ����฾�,Uܼŧ��7���a�	����������?�H�c�8�N���
���   �   ��Ŀ����)����Ѧ��ܒ�ʊx�tI���U価���`bF��8߽��M�`0v���˺���������rP���f�O���-!ܾ��
��&�)?�$ R�c^���a�3]�KNP�ئ<���#��5�x׾��f	`����򃚽�`������ ��90�d��L���ཾ'H��8��ds�Nq�i�K�}{�܆��"w��s鷿�����   �   ���6ￇ��r�Ͽҁ��n7���F��TG�a���Ͼ����w�����x���҈� ǰ; �ٻ������d����U�6���
����徢��8�#�����S#��������L�hq������M�"��t򖽨���@��<�k;l�мL����r�Tv�Ͼe��F�H����2���t9��p`ѿf%�8���   �   ���A�b������!�ܿ����������s�s�6����0���Q�w�޽��1� �r��sp<X�t< ,ֹ,!��������72��m����4��H?���;�Ѿ?�̾{Ҿ��䩾J���R/e��)��R��|��e��@r�;8�<|��< Mu:��!��׽�N����`�m�6���t�㪛�r����޿���������   �   ��)��&����Ƃ�� �	Bۿ���@���dX�M��pjоIj���\��t�(h�虥<\��<���<�!<0ȅ�L�{b���D��+�XpN��j��N{��?���y���e���H��$����P����>*�����Y�<b�
=�]=d�<�r.���^��L	�~��.ξO��B�W�T��"����ۿ"� �N;���� '��   �    M@�t�<�d&2���"�����h����˿z����
v�b1����5���τ*�������h�T�<�*=�=;=�a=�ط< �U9LbԼ�[[�	���Hս���R	�.m�I��8��Xʽ�I��|�<�l��hV<�^�<@@=��\=��J=���<���鐌�^�#�s5���[���/��Qt�=��iL˿�T��F��#�6�2���<��   �   �S�\�N���B���1�������n�ݿ!���ꪆ�tC��2�{���$A����`���4
�<|,G="qp=��l=
�G=0<=���<`1r�,����`!�cV���v����d|o�8!H�\��$2�� �o; y�<R�.=�Rl=8ň=�J�=��i=D�=PA�����e9����H��'�@�vW��5U��Æܿ>��i���1�d/C�P�N��   �   ,�_�P[�">N��a;�^�$�����;�M������lN�?m��n���O��'Ž����<F�V=lo�=�4�={߂=�[=�	#=�_�<��&<��0� �N�����ܝ��,<����`�;�<��=��D=�M=c��=�G�=@D�="~{=�=H�t��y���EG�>ί��
�uK��q���D���x��$�g$�� ;�6N�@[��   �   ��8�^s5���+�����
�֓�KĿE̛��7l���)�1澱����,��������=��x=���=x�=�(�=��=�e=$9=��=���<���<x`q<8�i<pO�<�q�<<'=�I7=�k=�R�=�I�=��=���=���=o
�=:�O=�<�=]��$��w��Hv�,'�K&i��;����¿�N�2N
�h����+�Rt5��   �   4�5��:2���(�0�Xo���鿜������^�g�N�&�_ᾐ͌�Hv�~[��@�G��/=u=��=�P�=^��=Qx=��J=�B=\��<X~<� <��^; �4;�c�;H;U<���<�?=L�J=���=O�=�.�=&M�=��=ߋ�=�O=hx"<r)T�04�i����۾��#�u
e�[���������迀�l��(�HE2��   �   
>,��
)�� ���@���޿*H��i#��'_[�`5�e�Ӿ�Z��X�%g� ��9o=��h=P�=Ty�=��g=��5=�)�<��]<�>���y�|�м
(�"�`�Ц� ����8<l�<�F/=�;q=��=���=,-�=�ȑ=~�K=سK<�5:����}�hϾu��Y�����\��3wݿv������; �~,)��   �   ���L�ڭ���"̿|!������G��n�f^���`i�]��|K:�@�;hx=�\R=�^_=��E=�l=p�<�����漨�L�a��������X����½�������|�|�:�%��b���.�;4�<L�H=�=%�=���=V�D=���<����|}a�a���|��HF��������h̿��  ��[�BV��   �   �B�	�X����￢DԿVC��1̔�l�i���.�s��uw��B}D�>uȽ ��hL*<��=��.=ƛ=�<`�+;�ϼԙi�`y���������2(0�L�=�d�A�RQ;���*�40�-�潼4��rw8��]O�X<{=��P=�]=�x6=,�<P�Ƽ������>�	��8����@.�L�i�i����ɵ�b$տ��pH�:7
��   �   )�P��7U��`ο�f��-<��x�}���E���`h;EW���^��������9u<,T�<xU�<�h�<&��d )��{���6�� 4�~c�w���r��X���c���퟾�`���؂���Y�TP)��G�𷐽L�qj;�I�<��!=��=���<�F��w�����$���̾�����F���~��.��ʢ��y�Ͽ⿯V��   �   M�ɿ�ƿ􌻿Zm������&��@{O�ё ���� ���L���g>� ˖��y�<��<(�J<��G��K� �ɽ�j ��b���������UӾu�꾮;����������M�羡2Ͼ9�������a�W���f���$��to���< -�<N�<�.P��4���߽��L������w�!��RQ�����g���ڬ�-���6�ƿ�   �   ���➿�5���و���o���I�{I"�gG���!���'p�r �� ��@#�����;���<�A<x�,�R}G��<ѽ�
.��������}ݾ��������)��3���6���2��(�á����r�׾�h���lv�;L%�r���R�,��C����<TO�<�
<����-���LH���s����������$��pL���r��:��*O���~���   �   Guy��Jt��[f�a�P�(�5�@���0��i��i�V�#��$���W��=��H�}<h�r<��Q�8_�'��"Z)�f��K���,!���u�G�8�6S�NRh��]u��yy�dOt�`f�;�P�� 6�.���5�m��O���#��*���_�@ʥ�p�}<��r<`NQ�bV�T ��hU)�8��)������r���8�5{S��Mh�+Yu��   �   ��6���2��(�q�����p�׾zd��cfv�0G%������,� ��@�<P�<(�
<𧴼>���L�;�s�Fĵ�i����$�<tL�}�r��<���Q��$�������䞿J8��܈���o���I�)L"��K���$���,p���+���-�� ��;���<8�A<i,�rG�5ѽw.���!���4ݾ}��j����)��3��   �   5���d���\��6-Ͼn���q�����W����%崽��$�`�n�(�<�1�<(M�<�Q�^4�G�߽̳L������!��UQ�����i���ܬ�����ñƿ��ɿDƿT����o��� �����~O�� ���뾬����L����l>����z�<t�<�K< ]G��K�b~ɽEe ���b�H�������RPӾc��T5���   �   �^��韾%\���Ԃ�8�Y��I)�s=ｈ���@e�@k;0W�<��!=6�=l��<0�F�O{�����'����̾���0�F���~��0��Ҥ����Ͽ��4Y+�̩�W�cο�h���=��7�}��E�����j;Y��6a��
���œ�@8u<,X�<l^�<w�<p�����(��r��P1�B4�_vc�$������0S���   �   �A�&J;�6�*��)�,��H+���g8�+O��><P�=��P=��]=Ry6=P
�<8�Ƽ7���j�>��������B.���i�����W˵�@&տ��I�h8
�8��h�	�l����_FԿ�D��p͔�n�i�*�.�gu��y��sD��wȽ����I*<.�=*�.=�=��< �,;dxϼ`�i��o������F��L!0��=��   �   ��½���[���8�|���%�`H�����;�&�<>�H=,�=��=h��=n�D=p��<<�����a��������IF����&ç��̿���� ��\�DW����6��������#̿"��׺��T�G��o��_��Lbi�����M:����;4y=_R=�b_=�E=�s=H��<1�� ��БL�����﫽�N���   �   j���� ���PW�� _<!�<�M/=LAq=�
�=���=5.�=ɑ=H�K=�K<�8:�<���}��Ͼ\��IY�����]��9xݿ������< �B-)��>,��)�b �N��ĸ��޿�H���#��`[��5�F�Ӿf[����&g� ��9�o=��h=cQ�={�=��g=��5=�8�<��]<@��h�y���м~��   �   `�4;`��;�QU<0�<XD=:�J=F��=��=�/�=�M�=	�=��=*O=�s"<|+T��4��i����۾Z�#�*e�ʢ��3���������F�(��E2���5�J;2��(�`0��o�	������ ����g���&�j_��͌��v��[���G�t0=u=���=�Q�=���=Tx=d�J=G=0��<�(~<8 < ._;�   �   H�i<`O�<�q�<'=TI7=lk=gR�=vI�=��=���=���=8
�=��O=8�<�>]�%��w���v�W'�{&i��;����¿�N�>N
�t����+�Xt5���8�Zs5�|�+����v�
����KĿ*̛��7l���)���{������������>�=&�x=㤕=Ex�=�(�=��=R�e=H$9=��=��<ؒ�<�`q<�   �   ��4;p��;�QU<(�<XD=8�J=O��=��=0�=N�=P�=j��=bO=�{"<�(T��3��h����۾��#�
e�!���d���$��F�&���(��D2�ʟ5�|:2�2�(��/� o�	�����O����g���&�6^��̌�Wu�Z����G��1=&u=!��=+R�=θ�=vTx=��J=FG=���<h)~<� < ._;�   �   `����0����W��(_<!�<�M/=|Aq=�
�=���=�.�=�ɑ=��K=ؼK<�2:� ���}��Ͼ���HY�f���[��bvݿ���j��<; ��+)�F=,�
)�� �
�����޿BG���"���][�m4���Ӿ�Y����� g� ��9xr=��h= R�=�{�=p�g=j�5=�9�<P�]< ��h�y�H�мp��   �   ��½���g���H�|��%�<H�����;�'�<��H=��=��=~��=�D=줂<V���潐{a�	�������FF��������9̿���2���Z�FU����R ������%!̿F �����t�G�Xm��\���]i�q��nE:��,�;D}=�aR=�d_=��E=u=�<�*�����d�L�a�����N���   �   �A�,J;�>�*�*�8��G+���g8�*O��@<D�=h�P=P�]=f}6=��<D�Ƽ2���L�>�o���}��P?.�S�i�0���=ȵ��"տ��\G�6
��}��	�6�����BԿ�A���ʔ��i���.�?p��Yu��,zD��pȽκ�Pe*<=��.=��=$#�< �,;,vϼ��i�1o��\���0��B!0��=��   �   �^��韾(\���Ԃ�>�Y��I)�f=�f���$d��k;�Z�<��!=��=0��<�eF��s��L�� #����̾����F���~�I-��堷�X�Ͽ(}�4T&�̤��R῱^ο�d��b:��j�}�\�E���\e;U���[���������Vu<�b�<�e�<�|�<����.�(�hr��1�4�>vc�������0S���   �   7���g���a��9-Ͼt���r�����W�����䴽��$� �n���<�:�<([�<�fN��4��߽�L�s���B�5�!��OQ����e��Sج�ʸ����ƿ��ɿ7 ƿ����k���������/xO�Q� �������s�L�f���\>�����t��<<!�<�K<XRG��K��}ɽ�d ���b�/�������FPӾ_��R5���   �   ��6���2��(�u�����r�׾xd��Xfv�G%�����<�,�0����'�<�]�<��
<0����񓽐D���s�X���p���O�$��mL���r��8���L��B|����� ����3���׈��o��I��F"��B�����H"p�8��=������>�;���<�B<�Z,��oG�4ѽ.��
�����ݾu��e����)��3��   �   Kuy��Jt��[f�f�P�,�5�A���0��i��R�$�#�$��pU� ����}<��r< �P��K�c���P)�.��<������o�<�8�RwS��Ih��Tu��py�yFt��Wf�g�P���5�(���+�e���
�N�#���L�@��ج}<P�r<`Q�S�0��U)���
������{r���8�2{S��Mh�+Yu��   �   ���➿6���و���o���I�|I"�gG���!���'p�& �����h���#�;��<�B<�B,��eG��,ѽ2 .����閭�ݾ�����Q�)�F�3�	�6��2�C(������,�׾`��G_v��A%�X���j�,�ศ�01�<�`�< �
<p��������G���s�����������$��pL���r��:��)O���~���   �   M�ɿ�ƿ����\m������*��B{O�ґ ���� ����L�3��>d>�@���t��<�$�<�-K<�2G���J��uɽ�_ ��b����䆵��JӾh��/��ɬ�����V�羧'Ͼ}���+�����W�ݗ��۴��$�@5n��#�<�A�<�\�< �N�4���߽U�L�����m�!��RQ�����g���ڬ�.���7�ƿ�   �   )�T��8U��`ο�f��0<��z�}���E���Xh;0W��~^����ظ��(Pu<�d�<�l�<���<�{����(�+j���+��4��nc�ⱆ���NN���Y��4䟾zW��8Ђ���Y�ZC)�W2�o����G� �k;�i�<��!=<�=���<XoF�Uv������$����̾�����F���~��.��ɢ��y�Ͽ⿱V��   �   �B�	�X����￤DԿYC��2̔�l�i���.�s��jw��}D�ntȽR��H]*<,=��.=�=�0�< H-;�]ϼyi��e��a������u0���=���A��B;�X�*��#�أ�j!��W8���N��k<^�=,Q=�]=&6=`�< �Ƽ����Z�>����#����@.�E�i�g����ɵ�a$տ��pH�:7
��   �   ���L�ܭ���"̿}!������G��n�^^��d`i�����I:���;�|=RcR=�g_=d�E=�{=x�<pԯ����&�L�Ė���嫽�D����½���Մ����|��%��,�� ��;�:�<T�H=��=��=���=
�D=H��<P����:}a�I���r���GF��������g̿�� ��[�BV��   �   
>,��
)�� ���B���޿,H��j#��)_[�_5�b�Ӿ�Z��.��#g� ��9�q=$�h=S�=}�=��g=��5=xG�<(�]< ��`�y���м������P�������`�<�2�<"U/=�Gq=]�=���=0�=�ʑ=��K=P�K<D4:�����}�YϾo��Y�����\��2wݿv������; ��,)��   �   4�5��:2���(�0�Xo���鿞������`�g�N�&�_ᾋ͌�4v�;[����G�b1=(u=y��=�R�=���=�Vx=��J=K=���<�=~<�5 <��_;@C5;���;�hU<�<DI=��J=+��=A�=X1�=O�=�==O=�|"<�(T�4�i����۾��#�s
e�Z���������迂�n��(�HE2��   �   �<����l'	��S���|޿���%����u��n8�"� {��wyT���ݽ����F<2,5=��=�y�=˯�=hޕ=E��=yw=��W=��9=�; =ƒ=��=�	=Q=\�1=`�T=RZ~=�Õ=��=Jſ=�!�=0��=���=ti�=7Ӌ=Z�	=�씼�J���F�8���, ���5�^s�i���,����ݿ	��x	����   �   :��z1����/ ��M�ڿ�̺�j��*[q�.�4�Jj �P����-O�h}ֽܔ��DY<d%6=���=ߐ�=���=�G�=Y�=b=�>=��=4�<l4�<��<���<��<Z=��2=��_=�[�=^��=U�=���=X�=���=�7�=�[�=~�=�������\9A�1���l]��\p2�po�r�����LKڿ;�������9��   �   �	��,��5 �y����Ͽ/e��z��Ofd��*�q�񾅢��(�?�����x꼼І<l8=�}y=k��=���=.5v=j5O=s =��<�ہ<�9�; �}��뚻� �%����;�̕<�*=�>=2�{=r��=�ί=!�= �=;j�=���=�5=PG<��/���73�+B����j�(���b�Dΐ�S���l�Ͽ�vS ��C��   �   2���������Pؿv���n������"&P����پt����'�4���U���¬<j :=tj= s=�\=�20=��<`�:<@�Ȼ���P��\5E�r�^�:!b�
�N�T�%�̎Ӽ� �XD<0m=�vP=���=���=�o�=�[�=#�=z�=���H����d��)���B־���P*O� Ȅ�����B��Ozؿ�M�?����   �   �]ῥ<ݿ��ѿ��h���ߏ�7jj��g6�!��|����}q�j�	�$�t�����@7�<2�7=�Q=<GB=�<=(��<�������c��Ĥ��1ѽ�<������ ��g�{N��jg��r���3�诀<"�=XBi=n<�=�	�=�t~=�(=�S�;��K������k������1��76���j�_J�����j���>pҿީݿ�   �   Z���(>���*�������֐���t��xF�mQ�ee�˙���@��Cн�� v�;��<D�.=��+=�-�<(D-<<����K��|�����L$�Q�D��<^��m�
r��Kj��;W���:��~�޽�4��P��@��:��<vWD=��l=�g=�J/=8�j<h ��;ƽ �=��0��Χ������G�Ӆv��ȑ����l��Ế��   �   CӠ�~���Z���Ї�n�G/H�	� �}2�����l�m�������@��<P�=
�=�T�<��<( ���V}��F޽��#���Z��䇾]������r��2s���^��O������ځ�H�L�������$�>���� v�<�(=|�E=��.=���<P�P��\�����o��O��f���ɪ"��AJ��Tp�U숿R����/���   �   $ ���{���l���V�LH;��O�C������4��z*��ٻ�|���T};l#�<�s=D��<Ќ7<௥��x���N�8�:�����O`����˾�\�e��w�
��A�Z�	��/����[Hƾ�!���Nv��-��Qٽ�^V���$����<ܣ=
�$=1�<�=�;0�½�/�&n��pn��PR��b���=��/Y�Q�n�<�{��   �   �)C���>�Y�3�&%"��G�y��i���Z����G5�z�׽]E�@��XI�<D�=�<=<��< �0���`��}�Ͻ>�T����.��WZ�|��cz$��K5���?��-C�L�>�Ó3�E("�QJ�2��M���rą��L5���׽(gE��M���A�<�=�==��<`�0��`��v�ȸ>�󊾻*��bU���(w$�
H5���?��   �   �>�A�	��,�O�群Cƾ����Gv���-�~Iٽ�RV�l$��<ʦ=��$=-�<��;(���½�	/� q��#r���V��(��F�=�83Y�/�n�B�{�,"���{���l�,�V�]K;�'R����������6��b*�`߻�����};��<�t=D��<��7<8����r��F򽮾:����\����˾GW�h��T�
��   �   n���Y��TJ��&����ց���L�"������>����`��<R(=��E=��.=t��<�P�&a��O����o��R��X���=�"��DJ��Wp�5W����1��cՠ�����Q���҇�Tn�2H�Q� �!6��ꓱ���m����	��\������<8�=$�=�]�<(�<����H}��=޽T�#�¾Z������X��ƪ��[���   �   r�Dj�(4W�8�:���A�޽5,���}��?�:���<]D=f�l=l�g=�I/=�j< �h@ƽH�=�!3�������s�G���v�Qʑ�񕥿g��񼾿l���.@���,��}���ؐ�A u��zF�:S�(h�͙���@��Gнr� a�;l�<��.=�+=�8�<8d-<�m���K�t������,	$�n�D�85^�@�m��   �   .�� ��\�qD��|^�����2��Ā<D�=�Hi=�>�=�
�=xu~=��(=�:�;@�K�����k�Ë��K3��96�F�j��K��]�����rҿīݿ�_῁>ݿF�ѿ*���oi��#᏿Clj��i6�c��Y�����q�6�	���t�����5�<�7=r�Q=ZKB=�B=h��<�����k���c�㻤��'ѽ�1�����   �   �b� �N��%��rӼ� ��JD<Pv=`~P=���=۝�=q�=�\�=A�=H�=p%��Ą���f�+���D־����+O��Ȅ�Ы��MC���{ؿ3O������3��O���T�뿥ؿ����q������x'P�%��e�پ�u���'��5���Y����<� :=�uj=�s=l�\=t80=��<h�:<��Ȼ캼���%E�V�^��   �   ����#�p5�;�ޕ<�2=��>=��{=Ι�=yЯ=r"�= �=�j�=ⱉ=b4=�P<��1��293�9C�����`�(�(�b��ΐ�+���`�Ͽ�T ��D���	�"-�6 �k�꿓�Ͽ�e���z��6gd���*�u��<����?����� 꼼φ<Zl8=�~y=^��=��=�8v=H:O=�x =0��<,�<���; g{�@����   �   ���<̙�<�^=��2=��_=5]�=���=5V�=ˡ�=�X�=;��=�7�={[�=��=�������M:A�ڒ��P^���p2�'o��r�����Kڿ�������,:�����1����� ����ڿ�̺�]j���[q�w�4�|j ������-O��}ֽ2���DY<�%6=��=_��=� �=�H�=���=$b=>=x�='�<�=�<��<�   �   �	=Q=N�1=B�T=2Z~=�Õ=��=2ſ=x!�=��=���=Hi�=Ӌ=̺	= eK��2F�n���, ��5�K^s�����,���ݿ�	��~	�����<����f'	��S���|޿����$����u�fn8����z��"yT�/�ݽV�� �F<�,5=��=�y�=诚=�ޕ=b��=:yw=ЮW=�9=�; =֒=̥=�   �   ܍�<ܙ�<�^=��2=��_=@]�=̣�=HV�=��=�X�=r��=08�=	\�=.�=���"���8A�푤�]��p2�o�Ar��F���Jڿ����L���9����(1�6�������ڿ̺��i��mZq���4��i �����u,O��{ֽn���LY< '6=���=ʑ�=� �=�H�=���=�b=x>=��=�'�<<>�<��<�   �   𚘻 #��5�;�ޕ<�2=�>=�{=뙙=�Я=�"�=p�=Mk�=벉=�7= ><��.���63�qA���쾾�(��b��͐�������Ͽ#��R �^C�V�	��+�5 �h����ϿSd��Wy��ed��*���a���z�?�3�����0׆<o8=��y=/��=�=:v=0;O=�y =���<(�<��;�S{�p����   �   �b��N�
�%��rӼ�� �(KD<|v=�~P=���==��=�q�=�]�=��=��=P����hc��(��:A־���)O�0Ǆ������@��yؿ8L쿱���}0��$���Q���ؿ&���F������$P�����پs��x�'��0��(K���ˬ<�:=�xj=6s=8�\=�90=���<��:<`�Ȼ�꺼����%E��^��   �   $�� ��\�rD���^������2�Hŀ<Ԍ=RIi==?�=��=�x~=@�(=�y�;��K����C�k������0�66���j�*I��k��Զ���nҿ�ݿ�[῿:ݿ��ѿ��uf���ޏ��gj�f6����0����zq���	�v�t��[��0B�<��7=��Q=NB=�D=��<`����h���c�{���T'ѽ�1�����   �   r��Cj�*4W�9�:���3�޽,��B}� R�:���<�^D=�l=*�g=�O/=`�j<� �i7ƽ��=��.��
����ńG�#�v�Ǒ�W�������ܸ��F���<���(��ᔤ��Ԑ���t�vF�fO�2bྡș�@�@�A>н��p��; �<��.=��+=�>�<�m-<�i��l�K�Ns�������$�D�D�5^�-�m��   �   	n���Y��UJ��'����ց���L������.�>��������<�(=z�E=f�.=��<�lP�X����Ȃo��L��������"�?J�_Qp��ꈿ\����-��(Ѡ�e���X��χ��n�S,H��� �q.��񍱾��m�N�� ��(݇���<:�=J=�e�<0�< ���F}�	=޽��#�v�Z������X������R���   �   �>�B�	��,�S�群Cƾ����Gv���-�?Iٽ�QV�Pf$�̯�<��=6�$=>�<�y�;�
���½�/�pk���j���M�������=�(,Y���n�@�{�����z�	�l�%�V�E;��L�����J���1���*��һ���� �};�2�<T{=0��<��7<�����q��-E�J�:�󢁾�[����˾5W�d��R�
��   �   �)C���>�[�3�'%"��G�{��h���T����G5��׽�[E����P�<��=`D=Ȫ�< �0�t�`��n�г>���&���P���� t$��D5�H�?�&C��>�ی3��!"��D�{��=�������~B5�;�׽bPE�ȼ��Y�<Ĥ="D=,��<Ƚ0���`��u�`�>��򊾖*��EU���!w$�H5���?��   �   $ ���{���l���V�OH;��O�D�������3��S*�Eٻ����@�};�,�<�z=$��< �7<@����k��l=�,�:������W����˾�Q�u��9�
�|;�!�	��)�Π羺>ƾq���@v��-�U@ٽTDV�?$���<��=��$=<�<p]�;@���½P/��m��Kn��1R��V���=��/Y�N�n�;�{��   �   GӠ����]���Ї�#n�I/H�
� �{2�����Q�m��������釼짉< �=x=�l�<��<����:}��4޽��#��Z��܇�8T������K���h���T��}E���|���ҁ���L�\�������>�@k�����<@(=��E=>�.=��<�|P��[�������o��O��I�����"��AJ��Tp�S숿R����/���   �   [���)>���*�������֐���t��xF�nQ�be�˙���@�&Cн��P��;��<�.=T�+=�G�< �-<�U��\yK�k������$���D��-^�d�m��q�$<j��,W�L�:������޽#���n����:�	�<
eD=�l=p�g=�O/=0�j<� ��:ƽ��=��0����������G�ͅv��ȑ����l��⺾��   �   �]ῧ<ݿ��ѿ��h���ߏ�:jj��g6�!��w����}q�5�	���t�`z��p>�<��7=��Q=fQB= J=�<`c��hP���c�����jѽ�&�$��E�� �wQ�,:��HU�����H�2��ۀ<��=Pi=�A�=z�=�z~=:�(=`k�;��K�*����k�{����1��76���j�]J�����k���?pҿ�ݿ�   �   2���������Qؿw���o������$&P���޺پwt����'��3��TR���Ǭ<6:=|yj=ls=��\=,?0=<��<0�:<�4ȻҺ����zE��^�p b�ĢN��w%��UӼ�s �pxD<�=��P==���=qs�=�^�=:�=z�=���������d��)���B־���J*O��Ǆ�����B��Nzؿ�M�A����   �   �	��,��5 �{����Ͽ1e��z��Ofd��*�o�񾁢���?�m���\	�Ԇ<zn8=R�y=؉�=⚇=:=v=v?O=6 =��<���<0��; �x�pH��0I�� � ����;�<�:=Z�>=R�{=���=�ү=V$�=��=l�=Q��=�7=�A<��/���73�B����e�(��b�Cΐ�R���l�Ͽ�vS ��C��   �   :��z1����1 ��O�ڿ�̺�j��,[q�/�4�Ij �N���w-O�N}ֽX��HY<�&6=���=	��=X�=�I�=���=b=�>=n�=�/�<LG�<���<���<���<zc=\�2=��_=
_�=S��=�W�=���=�Y�=��=�8�=N\�=p�=`���h��F9A�(���f]��Zp2�no�~r�����LKڿ<�������9��   �   )F�q>��Կ��¿!����ő�ϕm��9��@	�9?��ѿz��5�sČ�H<y�t�<
�7=�p=C��=l�=*�=t�}=,�l=p�[=��L=@�B=�>=�@=�yK=">^= �x=7�=�ϟ=q��=���=T��=���=��=���=��=�Q�=�_g=P]s<�53������)j�������o
7���k��/���L�� f¿��Կ6D��   �   u��zܿi	ѿ�@��ﳨ��2���Ai���5�Q��� �� �t���Oۆ�rY���<��9=�xo= ��=?�=�P�=�iq=��\=.FH=�96="�(=�"=>(#=�-=�@=��[=8�~=ޅ�=\ը=���=��=��=���=0=�=�=Ŭ=�?i=��<D�)�њ����d��Ե�v
��3� �g�!���$j���(���ѿɇܿ�   �   Yaտ3�ѿ��ƿ����h��Z���Э\�k+��!��i/��H^c�t��uk��f�����<�2?=4m=$y}=��x=�>f=��J=��+=Ф=���<߳<૗<�$�<P��<�W�<L�=v�+=��[=JƇ=�R�=Hu�=R��=���=�'�=? �=��=84n=���<T�Yg��U�u�������)�u�[�Jm�����������ƿ�ѿ�   �   }Ŀ5}��FV�����M�����w��I�t���]�p���+GH���޽�=6� [U:���<��E=�f=xj=6W=*z4=��=R�<x�< 6�8�=������� �����s�0ӹ�p��;���<��=F�a=NN�=ﱪ=�)�=W��=��=��=��t=x�<�N˼�c���<��\���}���r�H�4x�D͒��馿���ʹ���   �   "��辪�U����a��(b���$Z�q0�}Z�Gžp��P�%������漘69<��=�-K=ؒZ=0K=�}#=��<(�<�)�(�2�=�J�{���l��顽oڕ�Ը{��s7���ȼ�R����<j,=��x=���=�o�="��=�=�=��y=
a=��H��ڕ�����l��ëþ~4�`T0���Z�6ⁿ��:���
���   �   ?锿C��/���L{���[��Q8�����Dᾙġ��)W�����on�x9#�8��<�t+=��K=��D=0=\Y�< /:��ɼ��U�~����~۽ң����v|"�8w$�bY�����':����j�X�Լ@||;�w�<[T=�$�=�j�=�}�=�i{=0=�	�:xqO����j�U�3,��ӛ������9�/7]�]�|�/����]���   �   u�1p��qb�aM���2������.����z��P �㍮�L����<n
=~�==�dD=d�"=�'�<@0غB��S���	ݽ���L�?�r�b�
�}�S1���I���@�t���U���.��� ����g8�������<z]:=�fv=!څ=~�v=�33=�s<������#��N�R��W����!�4� 8O�v�c���p��   �   �EA�=�S�1�U� �y�
���q볾����_�3�O�սV A��w���<H`2=�0I=��2=���<@-$;V�;ݘ�1����6�hp�)ē��T���~��rf˾A�ξ3fɾa�������ؔ��M_�`9$�Ũ׽�ad�XVb�dɜ<D-=FRa=�mi=�C=�1�<��λ�V��彍�<�n����K�����r��"��m3���=��   �   JS�����|��̾[����]�<55�,��p�f�(�C��a�<��+=z�R=0VK=�#=@M<�?��Z5���� ���C��䆾�T��N�Ҿs�������-V�������]��υ̾����c�:5���佶�f���C��V�<��+=�R=�VK=\&=0,M<80���/��֋ ���C��ᆾ�P����Ҿs��`������   �   X�ξgaɾ֋������.����F_�04$�s�׽�Td�8/b��ל<-=�Ta=�ni=��C=+�<�ϻ��V�N&���<�=���^O��T��{u���"��p3���=�IA�'=�K�1�� ���
�ك��l�����3���սX)A� w�@��<j^2=�0I=��2=��<@�$;����֘����D�6��o�k����P���y���a˾�   �   �E���ꄾ��t�ԠU���.�������Y8����ƶ<dc:=�jv=ۅ=��v=23=s< �㼫��(#�GS�U����<���4��:O���c�L�p��u�| p�ub��cM�(�2������1���z��S �����0Y����<
=��==�eD=p�"=�1�<@?׺�������ݽ���C�?���b���}�j-���   �   q$�YS�/��5��0��~�j�@�Լ`,};��<�aT='�=<l�=>~�=li{==���:>xO�
���U��.���⾱����9��9]�M�|�Ú���_���ꔿ�������{��[��S8�����G��ơ�-W�`����un��J#�4~�<�s+=x�K= �D=�3=�d�< 1:̠ɼ~�U������u۽���6��hv"��   �   �ߡ�rѕ���{��c7�Tsȼ@�
�D��<�&,=��x=<��=Tq�=1��=T>�=��y=�^=X�H�ޕ�[��5n����þ�5�)V0��Z�nみH󓿮��O�����a��������b��Lc���&Z�0��[�@ž���l�%����l�� -9<��=�-K=>�Z=�K=�#=��<`�<`�P�D�=���{�攽�c���   �   ����P�s�Ps��P�;�ʴ<V�=��a=MQ�=T��=P+�=���=В�=	�=Ąt=4�<LV˼bf���<�^����^����H�
x�KΒ��ꦿS�������Ŀp~��mW��-���<��� x�!I����|_侟����HH��޽�@6� �T:���<��E=��f=Pj=$W=Z~4=B=`�<��<���(�=��x������   �   �ϟ<�g�<��=��+=�[=ɇ=*U�=3w�=���=��=�(�=� �=��=R3n=���<J��i�t
U����������)���[��m��Z��|�����ƿ�ѿCbտ�ѿ��ƿV�����綇���\��k+��"��40��j_c�<��$wk��p��H��<�2?=�m=Xz}=��x=�Af=� K=t�+=0�=,��<�<��<�4�<�   �   �-=~@=d�[=��~=a��=�֨=���=���=���=z��=�=�=�=�Ĭ=�>i=P�<2�)�@�����d�?յ��
���3���g������j��
)��5ѿG�ܿ�u�N{ܿ�	ѿA��<����2�� Bi�J�5����>!��r�t�c���ۆ��sY���<��9=:yo=T��=��=�Q�=Zkq=��\=�HH=�<6=��(=`"=(,#=�   �   �yK=$>^= �x=/�=�ϟ=b��=���=D��=���=֮�=t��=��=�Q�=l_g=�Zs<h63�S���*j�*������
7��k��/���L��.f¿��Կ:D�)F�k>�ܟԿ��¿����ő���m��9�y@	�?��z�z��5�Č��9y�T�<`�7=.p=[��=��=D�=��}=`�l=��[=�L=\�B=�>=&�@=�   �   �-=�@=��[=��~=m��=�֨=���=���=���=���=�=�=j�=\Ŭ=D@i=4�<^�)�2����d�@Ե�>
���3���g�Ⰾ��i��8(��QѿV�ܿ�t�[zܿ�ѿI@��|���&2���@i�g�5�ق�1 ���t�F��
چ�(jY�@��<�9=lzo=���=4�=R�=lq=��\=tIH=:=6=��(=�"=`,#=�   �   4П<,h�<�=��+=*�[=ɇ=7U�=Rw�= ��=V��=�(�=6!�=��=�5n=���<���e཮U�������K�)���[��l�����븵���ƿ;�ѿp`տH�ѿȝƿ�������������\�j+�9 ��7.��z\c����pk�0L��@��<x5?=m=R|}=d�x=Cf=�K=��+=B�=���<��<��<�5�<�   �   ���� �s��q����;�ʴ<��=ƪa=oQ�=���=�+�=��=���=8
�=N�t=�"�< G˼�`��*�<�y[��(|���&�H��x�Y̒��覿��������9Ŀ�{��U������A�����w�>I�,���[������DH��޽>86��vV:���<��E= �f=j=�W=t�4=(=lc�<��<���@�=�@w������   �   �ߡ�Kѕ���{��c7�sȼ@�
����<',="�x=���=�q�=��=�?�=&�y=e=��H��ו�Ŗ�k��ʩþ83��R0��Z�ၿ�����T	�����d���ߓ��R`���`���"Z��0��X��ž�
����%�����Ȗ��K9<��=|2K=�Z=,K=��#=��<��<`�����ޱ=�z�{��唽Yc���   �   �p$�FS�$��%�0��N�j�̔Լ�1};��<vbT=�'�=Bm�=��=(n{= =�ø: jO�����U�*��������9��4]���|�����a\���甿�������W{��[�2O8�����A�¡��%W����8fn�P#� ��<fz+=��K=8�D=l7=k�< �1:��ɼR�U������t۽@�����?v"��   �   �E���ꄾ��t�РU���.�����𯽂Y8��~��Ƕ<�d:=�lv=�܅=|�v=,93=�.s<�㼞��L#�(J�9O���������4�$5O�W�c���p� u��p��nb�^M���2���.���+����z��L �	����9����<�"
=��==*kD=��"=�8�<@�ֺ6}�Y��s
ݽ5����?�V�b�g�}�V-���   �   N�ξ`aɾԋ������,����F_�$4$�O�׽fTd�,b� ڜ<-=Xa=^si=��C=�>�<`�λ��V�C�6�<�����dH����꾑p�K�"��j3���=��BA��=�G�1��� ���
�b{��糾ǀ����3��սA� �v����<�f2=7I=��2=��<��$; ���՘����6���o�@���lP���y���a˾�   �   FS�����}��̾Y����]�.55����̴f���C��e�<Ј+=ƩR=�\K=�,=�KM<����)��և ���C��ކ�M���Ҿ��󾭶�
��eP�0��R��q���|̾t���XW��/5����@�f�x�C��r�<
�+=��R=�\K=+=x;M<�)��q.��@� ��C��ᆾ�P����ҾX��W������   �   �EA�=�T�1�U� �y�
���o볾����J�3��սfA��w���<d2=D6I=� 3=0�<`#%;����Ϙ����ۇ6���o�����SL��Nu���\˾g�ξ�\ɾ1���:���[���(@_��.$�W�׽NFd�� b��<�"-=�[a=�ti=@�C=:�<@�λ*�V���
�<�6����K������r���"��m3���=��   �   �u�2p��qb�aM���2������.����z��P ������I����<�
=<�==�kD=��"=|A�< ֺ�s�y���ݽS���?���b��}�x)���A���愾V�t���U���.����x篽�J8��O��ٶ<`k:=�qv=ޅ=x�v=N83=�#s<t�㼯��@#�<N��Q��2�����4��7O�q�c���p��   �   @锿C��0���L{���[��Q8�����Dᾒġ��)W�z���*nn�83#�4��<�x+=v�K=��D=�:=(u�<��3:��ɼ��U������k۽!��Z��Bp"��j$�.M�R��T��'��r�j�LxԼ��};؜�<�iT=i*�=o�=ր�=�n{=�	= e�:<oO�)���
�U�
,����⾼����9�)7]�Z�|�/����]���   �   $��辪�V����a��*b���$Z�q0�}Z�Fžj��8�%�y��P��0>9<��=�1K=ؘZ=TK=��#=l#�<h�<x��L�鼂�=�H�{�Rݔ�vZ���֡�Dȕ�,�{��S7�Vȼ`�	�dɨ<"0,=L�x=a��=�s�=~��=|@�=Z�y=�c=�H��ٕ����fl����þr4�WT0���Z�4ⁿ��:���
���   �   Ŀ7}��GV�� ���O�����w��I�w���]�l���GH�f�޽�<6� �U:Ј�<��E=f�f=`j=�W=&�4=,	=@p�<h�< ���|=��_��ꬼ0�����s���`b�;pߴ<��=��a=�T�=%��=�-�=���=���=�
�=^�t=� �<�K˼�b����<��\���}���k�H�0x�B͒��馿���δ���   �   Zaտ6�ѿ��ƿ����g��[���ѭ\�k+��!��i/��@^c�`���tk��_��,��<�4?=
m=}}=��x=REf=�K=��+=,�=���<���<�ʗ<LE�<8��<,x�<��=��+=�\=̇=�W�=py�=���=���=�)�=�!�=,�=�5n=D��<P��f཯U�e�������)�r�[�Hm�����������ƿ�ѿ�   �   u��zܿk	ѿ�@����2���Ai���5�Q��� ���t���1ۆ�xpY�4��<r�9=4zo=���=y�=�R�=zmq=j�\=�KH=�?6= �(=4"=0#=�-=� @=D�[=8�~=��=(ب=ꞽ=��=���=P��=:>�=��=�Ŭ=|@i=�<��)�����w�d��Ե�r
���3��g� ���#j���(���ѿʇܿ�   �   4��{���"���,����|��"U�,�(��g¾Mԅ�8�*��(���Y)������a�<�=&h.=P|<=g?=�<=�!9=��6=�~7=��;=��C=b�P=��a=�w=��=&P�=�`�=�l�=\u�=XK�=��=���=���=��=��=ؽ�=yΜ=.;3= )��5H��\i���y������Y�^�*��5T��s|�V��w!������   �   �C��j3��L^�����dx��.Q��(����e�h���t&��>��P$��V*�@]�<�O=(0=�1<=j�<=��7=X�1=*p,=�(*=�+=vL1=>�;=�K=�`=<�z=�'�=Jߞ=@ϱ=���=���=�e�=0��=���=���=���=��=�@�=�6= ו��x��z�6t��ַ�p����b'��`P���w�:���%f���=���   �   �����ƛ�RS���/��Vk�r�E��&��]��a汾�s�z��&��Bw�@c3;���<PS=p�4=�:=��4=.�(=��=�6=�=���<$��<HH�<Nd=�=�}4=^V=��}=���=\�=�{�=4��=,��=�#�=�?�=|g�=���=�P�=�,@=�`�;��Y����c�������..��?E��k��D���s���ݛ��   �   �Z��▎�����D!u�:XV��3�%5�%Mܾ#��k�V��;������=��0�3<���<d�)=�9=��5=�%=dC=���<��<0'd<��<��; �S;#�;��;8�i<4<�<�=�ZD=�|=�.�=˘�=[��=l�=6��=p��=u�=&F�=�N=77<x+�=���J�>b��|Dھk���3���V���u�����ξ���   �   N��J�{�(nm���W���;��������ӽ� a��{2��vн�y=� �û��<��=D59=ƛ<=8+=�x
=���<��><�&� �K����,�ܤ����ZL�8��xe�� ��� �D<Pv�<�wE=�n�=T�=

�=A�=>��=1/�=b'�=��]=��<X�Qɶ�.�*�G���䈽�<J��[��6�<��}X�G6n��|��   �   ��Y�%xU��I�6�� �0[�x�Ͼ�����?Y�ͷ	��[���ż`�%<� =\D7=H�F="�9=6g=0��<�_�;�.����D�H�o׈�����[���ɮȽ`6ǽҢ��Ƞ���7p���� �L� �C<��=@vc=�c�=���=��=�0�=�ۜ=ll=�U�<�jF�H󅽖���Z�Ki���Ҿ@����zw7�J.J��V��   �   .�1�V�-�HI#��@�pG��uѾ������o���!�z���L#'��e��i�<�#3=~R=��N=x.=Щ�<�/< 9g�j>&������ǽ�N��"����)�|
4��]5�0J-��N�~��r�˽ڔ��z���G� �<*E=[��={��=)ǡ=�b�=tv= �=`�R;�I)�x|ǽ��(���x�ˊ��!Y־e��%�_�$�w.��   �   >S
���O������$¾�˝��vq�v�*���ֽ&�V�p�'�藮<=.=�G]=*Kg=h9O=��= �<��&���-�����o"��#���J���m��O���h��fH����}���]�T�5��$
��ﺽ�oK��I��$�<��2=V�w= ��=M �=��y=��2=��<tG��������:��M��(⤾�SȾ��y9 �W���   �   ѱ̾�3Ǿjt��7���%�����\���"�".ֽ4�d���n�Į�<x,=��h=�^�=��t=��E=���<�t@:��מ��k�D�7�6#p��2��e1��-佾xɾ �̾8Ǿjx������b ����\�1�"��5ֽ��d���n�P��<�z,=��h=^�=h�t=��E=��< �A:t���ў�fh���7��p��/���-��&ཾ�sɾ�   �   �D��[����}���]���5��
�躽&cK�P�I�l4�<��2=~�w=n��=� �=p�y=�2=�<�S��������:�/P��J夾.WȾ��羾; �����U
�;���������¾ϝ��{q���*�A�ֽ�V���'�P��<`9.=�E]=ZJg= :O=��=�<м&��-�������M#�i�J�Ǹm�9L��`e���   �   �W5�dD-��H�l��b�˽���Z���G�@�<�E=���=1��=$ȡ=�b�=�v=��=��R;�P)�T�ǽ�(� y������\־yg��'�ʫ$��y.���1�ؿ-��K#��B�BK��^xѾj�����o��!������*'�@��La�<:!3=<R=��N=by.=���<C<�g�5&����f�ǽ%F��&���)��4��   �   1-ǽș��'����'p����pQL� &D<0�=(}c=�f�=~��=S�=L1�=�ۜ=8l=lP�< }F�������P�Z��k��ÂҾ������y7��0J�V�B�Y��zU�!I��6��"��\� �Ͼ�����BY�L�	�a_����ż��%<=�B7=ȽF=��9= i=��<���;��-�������H��Ј��{��䏽�ӥȽ�   �   �>���xK���A���E<4��<�E==r�=�V�=�=�B�=4��=�/�=I'�=@�]=p��<�!⼺̶���*�藅�����L������<��X��8n�<|�@O����{�Opm���W�r�;�B�����ս��b��G}2�Yzн�~=���û ��<N�=�49= �<=\+=B{
= Ŀ<X�><�s�@jK�𢼼��>�����   �   �;��i<�N�< 
=�bD=��|=�1�=3��=H��=��=@��=��=?u�=�E�=rN=�,7<�"+�>��;�J��c��YFھ���j�3��V�P�u�����ɿ���[��֗�������"u��YV�9�3�$6��NܾT$��@�V�:=������C����3<���<��)=��9=��5=%=�E=���<���<�>d<�<P4�;�PT;Pn�;�   �   &=ȃ4=FV= �}=��=��=j}�=���=f��=�$�=R@�=�g�=���=FP�=b+@=�O�;��Y�8�v�c�Ƴ��
�/��@E��k�\E��;t��<ޛ�L���@Ǜ��S��]0��Wk�I�E�='��^��3籾%s�{��'��(y��L3;���<�R=J�4=d�:=��4=��(=��=�9=�=���<T��<�S�<Tj=�   �   (�`=:�z=)�=���=pб=���=���=zf�=ƽ�= ��=��=���=��=�@�=�6= ���x�@{�<t�D׷�G���c'��aP�6�w������f���=��QD���3���^��a���zdx�M/Q�[�(�����񽾩����&�!?��
%�@_*��\�<jO="0=*2<=��<=� 8=��1=�q,=�**=B�+=O1=�;=�K=�   �   �w=��=(P�=�`�=�l�=Ou�=LK�=��=���=���=ʙ�=ډ�=���=FΜ=�:3=�=���H���i�׳y�ڮ���Y�z�*��5T��s|�`��}!�����4��w���"���,����|��"U��,���:¾&ԅ���*��(��Y)�@����b�<L�=\h.=x|<=Bg?=:�<=�!9=��6=�~7=�;=��C=x�P=��a=�   �   v�`=x�z=2)�=���=|б=���=���=�f�=ؽ�=��=0��=���=(�=*A�=��6= r���x�(z��t�Cַ�����Fb'��`P��w������e��==���C��3���]������Rcx�M.Q���(�2����ڭ���&�O=��:"��:*�D`�<Q=�0=�3<=,�<=�8=��1=�r,=�+*= �+=�O1=��;=N�K=�   �   �&=>�4=�V=`�}='��=��=~}�=؜�=���=�$�=�@�=Ph�=p��=HQ�=R.@=�q�;��Y� ���c�ڱ����-��>E��k�%D���r���ܛ�㸞��ś��R��!/��"k�a�E��%�<\��3屾s��x�\$���s�@�3;���<�U=(�4=�:=�4=��(=��=�;=R=���<���<hU�<k=�   �   p�;��i<|O�<r
=�bD=(�|=�1�=X��=x��=&�=���=���=2v�=ZG�=�N= D7<(+�p��A�J�a���Bھl����3��V��u�����۽���Y��蕎�˼��|u��VV���3��3�2Kܾ�!���V�:�ڶ���4����3<��<��)=�9=26=l%=I=���<�Ʀ<Hd<��<PA�;@eT;Pv�;�   �   �=����J��?���E<���<�E=jr�=W�=o�=C�=���=�0�=�(�=8�]=���<p⼼Ŷ���*�������G����z�<��{X�!4n��|��L���{��km���W���;�!�̈́���ѽ�T_��>x2��rн�r=�p\û��<V�=�99=��<=�+=L
=�˿<@�>< ��P_K�h�����Ė�����   �   �,ǽr���ꗝ�B'p�^��0PL�8'D<��=�}c=�f�=��=&�=�2�=�ݜ=�l=`�< QF�2���|�Z�g��?}Ҿ�����Tu7��+J�
V�(�Y��uU�HI�=6���kY���Ͼ8����;Y�ִ	�W��X�żx�%<�%=nI7=��F=�9=�m=��<p��;�-������H�jψ��z�����6�Ƚ�   �   �W5�;D-��H�X��G�˽�
��@�F�0�<�E=a��=
��=sɡ=�d�=<v=��=@SS;8A)��vǽ<�(�F�x�
����U־�c��#���$��t.���1�Ⱥ-��F#�?>�bC���qѾʠ����o�Ϋ!�����'� u���u�<l)3=R=��N=�~.=X��<�T<�g�H1&�����ǽ�D�������)�l4��   �   �D��I����}�v�]���5��
��纽�bK�P�I��5�<��2=*�w=���=��=�y=ܗ2=��<6��,����x�J:��J���ޤ��OȾV��47 �����P
�s�����f��S¾�ȝ�qq���*���ֽ��V��'����<RC.=�M]=�Pg=�?O=�=T�<��&�"�-�2���Q�#���J�O�m�L��=e���   �   ��̾�3Ǿct��1���!�����\���"� .ֽ��d�p�n����<��,=��h=�`�=��t=��E=��< �C: ��C˞�cd���7��p�9,���)��ܽ��oɾp�̾�/ǾIp��i��������\���"��%ֽ�d��cn����<~�,=��h=�a�=��t=@�E=h�<��B:��� О��g��7�p�R/���-��ཾ�sɾ�   �   8S
���K������ ¾�˝��vq�j�*���ֽ��V��'����<�>.=�J]=�Og=�?O=��=��<H�&�N�-���Z�F#���J�R�m��H���a��A�������}��]��5��
�xߺ�UK�8[I�G�<r�2=�w=I��=��=@�y=��2=��<@������~��:�RM���᤾MSȾX��l9 �N���   �   *�1�T�-�GI#��@�oG��uѾ����x�o���!�B����"'�@C��Hl�<8&3=8R=��N=r.=��<8e<h�f��(&�~����ǽ�<��֝�N�)���3��Q5�b>-�@C����˽����2��`EF��'�<�E=!�=��=�ʡ=�e�="v=��=@S;�F)�{ǽ#�(�,�x������X־le��%�V�$�
w.��   �   ��Y�&xU��I��6�� �.[�v�Ͼ�����?Y���	�m[��d�żX�%<�"=ZG7=��F=2�9=\o=���<��;�-�����,�H��Ȉ�ms��φ��^�Ƚ�#ǽY���'����p�����L�xSD<��=�c=�i�=D��=��=�3�="ޜ=Fl=t\�<_F��
��h�Z�i���Ҿ-��ި�qw7�D.J��V��   �   N��M�{�)nm���W���;��������ӽ�a���z2��vнy=���û �<*�=�89=l�<=~+=.�
=�ѿ<��>< ��?K�H�����v�����,0����<0��pܙ�0JE<|��<��E=�u�=�Y�=��=�D�=,��=�1�=;)�=��]=��<��Yȶ���*��������J��N��-�<��}X�F6n��|��   �   �Z��㖎�����F!u�<XV��3�$5�#Mܾ#��`�V��;����p<��p�3<܍�<Π)=\�9=~6=�%=K=��<TϦ<�]d<8�<�~�;��T;��;�i�;0#j<b�<*=�jD=4�|=�4�=ꝳ=���=��=��=���=�v�=G�=
N=@>7<�+����ҍJ�b��bDھ`���3���V���u�����Ͼ���   �   �����ƛ�SS���/��Wk�q�E��&��]��^汾�s�z�a&���v��m3;���<�T=��4=�:=��4=.�(=��=L>=�=���<\��<D`�<�p=�,=J�4=� V=��}=���=��={�=���=��=�%�=rA�=�h�=���=dQ�=�-@=pj�;��Y�����c�������(.��?E��k��D���s���ݛ��   �   �C��l3��O^�����dx��.Q��(����d�g���p&��>�� $�@Q*�<^�<`P=20=h3<=N�<=L8=l�1=�s,=L-*=�+=�Q1=�;=�K=`�`=f�z=�*�=�=�ѱ=���=���=hg�=���=���=���=P��=e�=GA�=��6= ���rx�hz�!t��ַ�j����b'��`P���w�:���&f���=���   �   j�q��l�Z�_���J���0������뾺ݳ�(��Bn1�>sངb�������[;��< ;,<��(<��!<�)<��L<Ģ�<���<���<�x=4�:=�
`=Y�=�i�=��=�Q�=��=��=��=�w�=�>k�>F�>���=��= ľ=#��=�P=�{[�ꔽ�7�ݤq��ϭ�TM�s���?0���J�r�_�!�l��   �   �&m�v�h�p[�		G��Y-����"�󯾊!~�\�,���ؽ��s�p�޼��׻C�;Pa)<��?<(�6<�C)<@�)<�C<@�z<|B�<pH�<�u=`�,=,�P=��u=��=0��=�v�=���=���=X9�=��=x>�>��>�!�=���="��=�q�=,&
=|@�.����^��Hl�S=������k�,�Z�F�g~[���h��   �   �n`��
\�T{O�2<�x�#�0K��پӗ���2l�����5ý60Q�0����hi�`V"<��l<H�u<�D]<��<<�F&<h�%<8N?<�Lr<8�<���<��=<!=��C=�i=)��=b��=���=Q�=R��=��=6��=���=l-�=	�=h�=2�=���=��=@\�����I�,�\����־���(w#�`,<���O��/\��   �   ΐL��sH��<���*�$A�>J���2þP撾r:P�<��� ���C�����<�Q�<��<腢<��<؇Q<x�<���;��;PC�;�B�;pU<��Y<p��<���<�= �:=�h=���=�'�=,F�=n��=�,�=d�=��=��=ܶ�=j}�=�,�=H�$= �q�	S�T��HE�:��)0¾Dy������[+�6F=�ϷH��   �   Y3���/�;#%���� ���Ծ�|����x���,��ڽ�Bk�x��� �;��<l��<H��<�F�<(*�<�/X<���; P�� �˻h�0�xc���w���i���3�0X���lb;ȫl<���<P5+=�h=���=X��=3|�=v3�=N%�=8��=p)�=��=�F�=
46=�:
<~��Hr½]'�a5x�ڙ��*�־���V���%��0��   �   ���9��Vw
����C1־��K���iF�
�����xC� ����+�<��=�=^I=��<A�<��>< <i9��;����vw��-��]H�x7W��W��8F��3$�X伨KI����;��<x�1=��y=�(�=���=�w�=XR�=]��=>��=d��=��F=�ʌ<�P��#���F��;L��2��vó�-2ھm��B��8��   �   �%��1�0�ݾ�Kƾ����È��O�����_����1��� �<�<*�=l�5=�9>=N�.=$
=xR�<�\�;�� ��/伒�=�_���%��Q���{ӽϜ۽�m׽�tƽ�j���:���'�4�� k<�}=�yU=�Ҍ=DB�=$��=�(�=\ߨ=&�=v�R=���<�����N��u̽���n�^�j᏾�`��qY˾�G�f��   �   ~���9���c���0����z��EF����ݼ���E�P^=����<��=�wP=0�f=(b=TE=�=$�<����D˼�O�Mힽ}Xֽ&��b���+���4�x5�FL,�D���l� rɽ�l�� �0���x��<l:=\$=���=���=�=�=^1W=���<�g;̨��E.���콦;(�ʓ[�p���<T���K��ƹ���   �   N���QA���no��P��*���z�� �:�XB/��<��'=��g=n}�=�+�=�'=\�R=�=��T<�
c�f�8�̛����8��&�C���c��|�����c ��ZD��qto�l�P���*���耭�J�:�pf/��ٖ<F�'=��g=�{�=�*�=b&=�R=�=��T<��b��8�I�����y����C�t�c�B�|������   �   F5�$G,�\��hh�	jɽ�e��$�𯂻d¼<�:=d)=�Õ= �=��=v�=1W=h��<��f;p���2��:��?(��[����+W���N��/������N=���f���3���z�JF����)㼽�F�@}=�h��<�=&tP=t�f=4&b=dE=*�=��<@���l˼��N�r螽TRֽ`"�r^���+���4��   �   �e׽�lƽ�b���3����'����ؒ<��=R�U=�Ռ=bD�=���=�)�=�==&�=��R= ��<����N�z̽���=�^��㏾bc���\˾K�	ﾀ)�q5��ݾ�Nƾs��Gƈ��O�����d����1�� � 2�<F�=Z�5=H7>=��.=�	=�S�<l�;p� ��$��=�����;�������|sӽ��۽�   �   j+F��&$�0���I�`�;�1�<|�1=x�y=�+�=ӕ�=�y�=�S�=1��=���=L��=>�F=�Ō<�Y��h������ >L��4���ų�5ھHp�����9����
��y
����4־I����M���lF��������I� }��$�<t�=��=�G=��<�@�<��>< zk9P�;�����<p��-�XSH��+W��W��   �   p	���	c;��l<���<z=+=�h=ά�=꼬=T~�=,5�=�&�=(��=*�=J��=�F�=�26=�/
<ڣ�}u½T_'�V8x�����t�־����X�%��0��Z3�Y�/��$%��R� �%վV~��v�x�ּ,�[ڽtHk�P��� �;�<���<���<$D�<�(�<�0X<��; ��@p˻�}0�x�b���w�؛i���3��   �   ���<��=҆:=H�h=���=9*�=nH�=P��=.�=��=Ύ�=@�=2��=p}�=�,�=$= ����S�.��<E�����1¾={��ά��\+��G=�B�H�D�L�3uH�r�<���*�3B�	L��4þ|璾I<P�����"��xG�����<�M�<@�<`��<D�<H�Q<��<���;� �;P_�;�f�;�j< �Y<���<�   �   ��C="i=Z��=t��=���=��=���=F��=.��=\��=�-�=`	�=��="�=c��=8�=`m绚���K���\����־���x#�S-<���O��0\��o`��\�F|O�<�8�#��K��پ�����3l�~��7ý�2Q������i��P"<��l<P�u<PB]<��<<�G&<�%<`T?<�Ur<��<`��<��=�!=�   �   �u=��=D��=�w�=���=���=:�=���=�>�>��>�!�=|��=���=�q�=B%
=��@�6���@_��Il��=��ѿ�����,���F��~[���h�-'m���h��p[�t	G�
Z-�`���"�d�"~�,�L�ؽ��s�(�޼ �׻@=�;�^)<h�?<��6<0C)<��)<��C<��z<�D�<TK�<rw=T�,=R�P=�   �   g�=�i�=��=�Q�=��=���=��=�w�=�>g�><�>���=���=�þ=�=2P=X~[�]ꔽ8�#�q��ϭ�~M辆���?0���J�}�_�&�l�j�q��l�L�_�p�J���0������뾓ݳ��'��n1��r�b�������[; �<X;,<�(<0�!<x�)<h�L<$��<��<��<�x=T�:=�
`=�   �   ��u=�=j��=�w�=���=���=$:�=���=�> >�>�!�=���=f��=$r�=�&
=Hx@�����(^�VHl��<���������,���F��}[�x�h�&m��h��o[�~G�0Y-�����!�f򯾀 ~���,�\�ؽ��s��޼��׻N�;�f)<`�?<`�6<�J)< �)<x�C<��z<pG�<�M�<rx="�,=��P=�   �   �C=�i=���=���=���=�=���=f��=X��=���=<.�=�	�=�=��=���=n�=�I绂����H���\��퟾~�־D��iv#��+<�̰O��.\��m`��	\�IzO�8<���#�jJ�rپ�����0l�&��Z3ý�,Q�(寮��h�x`"< �l<��u<Q]<�<<PU&<�%< `?<�_r<X�<(��<T�=�!=�   �   ���<�=��:=��h=���=r*�=�H�=|��=D.�=��=&��=��=���=�~�=+.�=B�$=  7�ZS�W��bE����.¾ww�����VZ+��D=�d�H�Z�L�TrH���<�Q�*��?�-H���0þ�䒾"8P�h�����?������<�X�<�%�<荢<�'�<8�Q<ȱ<@��; A�; |�;p�;Pu<��Y<��<�   �   `����c;H�l<���<�=+=&h=���=��=�~�=~5�='�=¬�=�*�=���=�H�=�76=�M
<|���n½�Z'�h2x������־b�����%�20�XW3��/��!%���� ���Ծ�z��A�x��,��ڽ<k�,�����;�#�<H��<|��<�P�<(5�<�HX<���; j�I˻xl0���b���w� �i�ؘ3��   �   �)F�D%$�h��I���;t2�<��1=��y=�+�=(��=1z�=GT�=.��=��=i��=4�F=֌<�B��З������7L��0��	���X/ھ�i�����46���Y���u
��	��J.־[����I��fF�*��B���;� ���6�<��=$ =�N=`!�<LN�<��>< �q9@�;���k��-�
PH�)W��W��   �   �d׽	lƽ5b��E3���'����x�<d�=ȀU=�Ռ=�D�=n��=�*�=��=n(�=��R=��<x��X�N��o̽,��7�^��ޏ��]��5V˾Dᾰ��!�.��ݾaHƾ���V�����O����Z����1�� � I�<�=��5= ?>=(�.=�=<a�<��;P� �L�ĕ=�1���E���ـ��+rӽ��۽�   �   �5��F,�-��Ch��iɽ`e��������`ü<h:=B*=|ĕ=
�=q�=��=7W=b =��g;����(���콊7(��[��~��&Q��LH��@���nz��X6��`��z-��2�z��@F����<ּ���E�:=��΍<B�=�}P=��f=�-b=v!E=�=��<�ʩ�l˼�N��垽Pֽr!��]�B�+�#�4��   �   *���4A���no��P��*����y����:��@/�(�<��'=*�g=R~�=-�=�+=��R=Z=0U<��b��8�����b������C���c�4�|�f������&>���ho���P��*�R��r����:�X/����<��'=��g=5��=s.�=x-=��R==0U<��b���8�Ô�����|��ژC���c���|�^����   �   �}���9��rc���0����z�tEF�����ܼ�^�E�0\=���<��=hyP=��f=�+b= E=��=���<�{����ʼ��N��ួgJֽ���Y���+�$�4��
5��A,�.���c�laɽ^��:��X��tԼ<F:=�/=�ƕ=��=��=3��=>7W=h =�jg;�����+��콮:(��[�����S��qK�������   �   �%�1�(�ݾ�Kƾ����È��O�����_����1�X� ��=�<t�=P�5=d<>=V�.=�=�a�<��;h� ��� �=���������Cz���jӽ��۽q\׽�cƽZ���+��@�'�p��P�<&�=��U=�،=*G�=0��=I,�=b�=�(�=v�R= ��<���f�N��s̽�����^�᏾V`��<Y˾sG�K��   �   ���4��Sw
����A1־ꊯ��K���iF�������C� ����-�<�=V�=�L=��<XM�< �>< �s9�;�@㺼�d�t-�FH��W�|�V��F�,$�����H� >�;�E�<N�1=��y=�.�=���=|�=�U�=8��=���=���=��F=�Ҍ<�I��p������^:L�c2��6ó��1ھ�l��5��8��   �   Y3���/�;#%���� ���Ծ�|����x���,��ڽ�Bk�|��� �;,�<���<8��<�M�<t3�<�HX<��; ^��.˻�Y0���b�H�w�@pi�t3���� �c;��l<�<NF+=�h=7��=俬=ڀ�=T7�=z(�=ޭ�=�+�=��=�H�=:76=�F
<����p½�\'��4x�������־���I���%��0��   �   ΐL��sH� �<���*�$A�>J���2þM撾j:P�0��� ���C��� �<$T�<"�<Ԋ�<�%�<��Q<�<���;�Q�;���; ��;`�<�Z<谜< ��<ڰ=X�:=T�h=�Ì=-�=�J�=z��=�/�=<�=<��=��=���=�~�=..�=��$= `O� S�h���E���0¾&y������[+�2F=�ηH��   �   �n`��
\�U{O�3<�z�#�0K��پї���2l����x5ý�/Q����� Gi��Y"<H�l<p�u<�M]<H�<<XU&<�%<�d?<gr<8�<@��<��=�!!=(�C=8i=ȝ�=���=���=��=p��=���=j��=p��=�.�=D
�=z�=�=���=�=�Q�i����I���\�pm�־���"w#�[,<���O��/\��   �   �&m�w�h�p[�
	G��Y-����"�󯾇!~�W�,���ؽ��s��޼��׻�E�;hc)<h�?<P�6< I)<��)<��C<H�z<�H�<�O�<�y=��,=ҘP=��u=�=s��=�x�=���=���=�:�=X��=>@ >/�>4"�=��=���==r�=�&
=`y@�ए�l^��Hl�H=��
����j�,�Y�F�g~[���h��   �   f�!�pU���yZ�j��x��1h��2f��c&�e��*��� :O��1����&����h�3���F��N���F���-�2���ۡ�x���A7<@��<�t1=�o=HB�=���=���=4�=���=T��=v�>�>��	>Qw>8�>���=0��=��=�u=�8�<$r���1��e	�h�S��Ւ�zz���羁#���A]��   �   ɂ�mE���Ѫ����hZ��c󔾃�`�I�!�]޽o����!D�x�����Q���}�~�*��o>��*G���@�4�)����(������PK!<���<B;(=b�d=���=	�=�(�=���= ��=p��=�>#�>��>�`>P�>��=���=�^�=\6v=(t�<����������6O�\Џ�J���M�⾔����HT��   �   ɂ�Kc���	�Q�����վ�g���슾PPP��L�%IȽ�����#�T߼�d���IƼ�����<-&��2��(0�~��$:��pc��p���E�;0i�<��=��D=6N{=$��=83�=��=��=�\�=0;�=�>�>P>Z >J��=�K�=���=L�x=���<K��%�\�����A����SѮ�*�վY��/�	�T���   �   ́�Q��*���o�߾�2���ʝ�{�v�*�6��������G��Ἄk����D�a������Ѽ ��v���q�Ĵ���������/Z�@���<<��<.1=�?=zms=��=vY�=g��=��=���=v{�=��=���=���=Ly�=�t�=&a�=��{= =�=ػ6�W�R�۽��-�.s��	��~X���������&���   �   -�뾩,��`׾����褾\<����N�m����Ƚ
�r�����c?� 
���m�: �%���л@/a�dԬ� j޼�-��s������m����(�x��ݻ ;<;��^<Tz�<B(=��P=�{�=5��=�=>��=h��=��= ��=h �=���=���=V�=h�{=T�= ����~)�{U��v���mR��'��|&��2�þ8�پ\P��   �   �,ľb���	��s��%A���uW�{E"���*����pw ��C�;Еv<���<h�d<@Q�;������'��ę�P�ԼR� �����p��t����d��� �v�@��� <<@��<Z�=��Z=�G�=��=x8�=Ea�=�j�=�\�=�t�=��=���=$�v=��=�"�;d���m��A���n.�,ud��R��x������V����   �   �����ږ�̗����u�M�Ey ��t�-������!���H<���<R=41=�,�<���<�3< ��8,G��/��b�
�v91�΍Q�>Uj�΁y��|�P�r�Y�x_0��󼐏\� E�;�ٿ< 	+=�o=�ؔ=H
�=�>�=^��=j��=!9�=��=vij=��=xs/<ĳ���S`����l�
��6��`�����*�5����   �   �i��`�Q&M��Y1������ս
H��ک��9ǻ��<j=Ҏ7=�$J=ZF=~�/=�A	=l��<�j�;��
��Lʼʀ(���j��|���꯽��Ž�ӽ��ֽ�<Ͻ�)��ET���'o�,K�8�V���#<JV =>jK=s3�=�z�=��=�G�=Ҙ=d��=zkT=�=�tP<P�I�`&�iU���սt(���+�|G�,I\��1h��   �   ��#�B��_�	��4彫��He�0Sݼ �Ѹ��<F+=(ta=Z��=�~�=��=�b=��3=�+�<xs=<�Z
�����4�[�g�D4Ͻ �������"���$��#�j��d�	�\<�\"���Se�Hgݼ ����<L+=oa=(��=�|�=��=�b=��3=h(�<Xq=<XW
����Ծ[�"�/Ͻ����h������$��   �   �5Ͻ�"��sM��Bo��?���V���#<�] =�pK=!6�=�|�=��=bI�=yӘ=��=mT=Z=XsP<��I��&�LX���ս+���+��G�tM\��6h���i���`��*M��]1�L���ս�M��
���vǻ ��<�=
�7=P J=>VF=}/=�>	=��< _�;��
��Jʼ�}(���j�ky���毽Q~Ž~ӽ�ֽ�   �   �Y�T0�X��e\�0��;��<f+=h�o=K۔=��=t@�=���=���=>:�=��=^jj=��=�n/<8���>X`�=����
��6���`�۱���󐾲������4ݖ�2�����u�
M��| ��z��1�����<��nH<ش�<�z= -=d%�<���<��2< ��1G��/����
�@61�؈Q��Nj�|yy�d�|��xr��   �   �v�����X_<��<�=j�Z=�J�=B�=�:�="c�=>l�=^�=�u�=��=2��=h�v=��=p�; ��������bq.�Pxd��T��.z��\�������{/ľ������Ou��C��6yW�HH"��������P� ���;8�v<���<�d<04�;��P�'�8ș��Լ�� �H�6�����P�h��������   �   ��^<Ї�<�.=��P=�~�=ݸ�=h�=D��="��=H�=X��=^�=D��=$��=��=H�{=V�= ���R�)�!X��M���oR�)��H(��B�þz�پ�R羘��/�c׾)����ꤾ�=���N����7�Ƚ��r������t?�@������: �&�pѻ@<a�ڬ��n޼`0��`s�<����i�X����x��qݻ �<;�   �   �5=��?=8rs=�
�=�[�=T��=�
�=B��=�|�=��=V��=���=�y�=$u�=:a�= �{=���<�Nػ��W���۽<�-�T�s�@��Z��m������)��ӂ�P��
���#�߾4���˝���v��6�P���h����G�8�,r��x�D�X�a�����̊Ѽ������6s������������'Z� j���<���<�   �   ��D=HQ{=���=�4�=q��=��=^�=&<�=>Z�>�>� >���=L�=w��=��x=���<@K��(�N�����A�x��UҮ�W�վ�����	������d�R�	�������վlh��|튾~QP��M��JȽ
�� �#��߼|i��NƼ\�����0/&�D2��)0�*��X:��@b������S�;�m�<\�=�   �   �d=k��=�	�=C)�=V��=���=���=A�>V�>˗>�`>f�>6��=���={^�=�5v=�r�<`���頌�T�T7O��Џ�ⴹ������H��T�-���E�i�������Z�����`���!��]޽����"D�����@T���~���*��p>��+G�R�@���)���(������O!<���<�<(=�   �   �o=ZB�=��=���=4�=���=N��=x�>�>��	>Mw>/�>���=��==|u=�7�<Ts��62��8e	���S��Ւ��z���羌#���F]�f�!�lU���mZ��i��x��h��f��c&�#�������9O��1����&����~�3���F��N��F���-���ۡ�@v���B7<���<�t1=�   �   ��d=���=
�=p)�=x��=Ծ�=��=J�>b�>՗>a>y�>r��=���=�^�=$7v=�u�<��Z���M� 6O�Џ�೹�ˊ�G�����S�b��E����n��ܡ��Y���򔾙�`���!��[޽n����D�������N��|�̩*�n>��(G���@���)�����#���q��8U!<t��<�=(=�   �   �D=nR{=��=5�=���= 	�=,^�=L<�=3>n�>�>� >���=�L�=X��= �x=8��<P	K��"�^���d�A����hЮ�վ����	�������b��	�����|�վnf���늾�NP�zK�GȽ���j�#��߼L_���CƼ��|��)&��2��$0�6��41��4Z����� k�;tr�<>�=�   �   �7=Z�?=hss=c�=�[�=���=�
�=z��=�|�=<�=���=��=fz�=�u�=ib�=z�{=� =�ػ8�W�B�۽��-��|s�����V���������"���F��)�����߾�0��ɝ���v��6�
���7���H�G���Ἔc���D��na�~���{Ѽ$�����k��������h���Z�`)��<蹱<�   �   �_<���<N0=��P= �=+��=��=���=f��=��=���=��=���=$��=�=N�{=��= `��Nx)��Q�����jR��%���$���þ�پ�M羬��2*�s^׾�����椾�:����N������ȽR�r�����O?�@p����: z$�p�л`a��Ǭ��\޼���6k�(����\����h�x��Rݻ �<;�   �   p�v�����He<(	�<��=�Z=(K�=��=�:�=sc�=�l�=�^�=�v�=��=Ɩ�=��v=��=`V�;D����������k.��qd��P���u��t�������2*ľ���	���p��	?��,rW�SB"�Ӥ�����B	�H^ �0q�;8�v<X��<�e< ��;�����u'�����,�Լ� �"����z������,����   �   	Y�R0�T��Pa\�`��;<�<�+=��o=�۔=��=�@�=���=���=^;�=%�=�nj==H�/<����I`����
��6��}`�`��������ҥ�� ؖ�=�����u��M��u ��n罾'���������H<���<��=�6=�8�<���<�3< ��h	G������
�.1���Q�BHj�8ty�"�|�8ur��   �   �4Ͻ"���L��@o��>��V��#<:^ =qK=i6�=K}�=d�=#J�=�Ԙ=��=pqT=\%=��P<��I�F&��O��Bս�$�^�+�lwG�AD\��,h��i��~`�z!M�"U1������ս�A�������ƻ��<�=��7=.*J=�_F=��/=0H	=(��<p��;Ƞ
�88ʼLu(��j��u���㯽�{Ž�ӽn�ֽ�   �   6�#�ڂ��	��4�V��zGe�PRݼ �и���<�+=�ta=ܧ�=e�=��=�"b=��3=�6�<�=<�3
�ď��f�[��螽�(Ͻ����&��z�L�$��#��~� �	��,�c��,;e�=ݼ ྸ	�<*+=Fza=*��=m��=��=�%b=`�3=<:�<�=<�4
�P����[��랽�,Ͻ����P���F�$��   �   ��i���`�&M�oY1�t��m�ս�G��|��`6ǻ��<=��7=�%J=�[F=��/=E	=��<p��;��
��6ʼs(�Ȟj��r��e߯��vŽ�
ӽڵֽ�-Ͻ����E��2o��2��dV� �#<0f =�wK=?9�=��=l�=�K�=֘=P��=ZsT=�&=(�P<؋I� &�
R���ս'�p�+�{G�pH\�W1h��   �   a����ږ�����i�u�M�.y ��t��,��L��( ���H<,��<N�=�2=�0�<���<83< ��G������
�v+1�*}Q�Bj�^ly���|��jr���X��F0����X6\���;���<�+=��o=iޔ=I�=�B�=H��=��=�<�=�=*pj=�=��/<𦡼�M`���+�
�Ԗ6�(�`�b����������   �   �,ľN���	��s��A���uW�jE"������F��u �@H�;��v<ఋ< �d<�c�;@#��H�'������Լ� ���8��0��j����\��� ^v�pY����< �<��=.�Z=MN�=<�=F=�=ne�=Ln�=�_�=�w�=��=z��=��v=��=�M�;,���������m.�Qtd��R���w������.����   �   �뾜,��`׾����褾T<��{�N�^����Ƚ��r�x����a?�@������: f%���лx%a��ͬ�ta޼P"���k������Y�l��� �x��*ݻ�)=;�_<���<�6=T�P=��==�=���=2��=	�=��=��=���=ޞ�=��=��{=��= ����z)��S������lR�7'��:&����þ�پCP��   �   ȁ�N��(���l�߾�2���ʝ�w�v�"�6�k���������G���ἰj��P�D��{a������Ѽ���V���m��������0��pZ�@��<���<$<=��?=xs=��=^�=���=��=��=<~�=d�=���=���={�=zv�=�b�=��{=( =�%ػh�W��۽��-��~s��	��RX������������   �   Ȃ�Kc���	�O�����վ�g���슾KPP��L�IȽ���P�#��߼d��pHƼP���~��+&��2�"&0�@��,2���Y�����v�;Dv�<��=��D=HU{=���=y6�=��=h
�=V_�=V=�=�>΃>�>� >h��= M�=���=L�x=���<�K�$�����G�A�~��0Ѯ��վF��(�	�P���   �   Ȃ�lE���Ъ����iZ��a󔾂�`�I�!�]޽e���f!D�P�L��`Q��:}���*�"o>��)G�j�@���)���$��@p��0W!<���<�>(=�d=b��=�
�=*�=$��=z��=���=��>��>�>,a>��>���=��=_�=X7v=v�< 􅼚�����\6O�HЏ�<���A�⾐����GT��   �   ��ɾEž����cy��+���bCi���7����ٚѽ�0���焽�e}�W���!?����Ž�n�~N�e����F��K�|�ὲӲ�Z {������lٕ<h*=x�~=�G�=���=�:�=��=�>e>�>;�>�>f>�  >��=���='A�=�0]=�< �p��o�A�ݽ
P&�̴_���������gw��H+ž�   �   �[ž��������ա�.���d�c���2�����Vʽ嵙�@�}���q�����	ҝ��
���⽧{ ��+��2�ې��W ��ݽOq���)w��C
�`���?�<�%=��x=�٠=B�=Ψ�=H1�=�} >Ō>�H
>v�>�x
>j>0.�=��=n��=�W�=��\=�l�<@�b�ԁi���ؽ��"��[�t舾Y������6"���   �   �U��J���;��SF��Q>����R���$��9��~5��ۆ�ڔZ��O���e��"������̽���� �(��K�����Ͻ/��:�l�x�� ��Xs<�s=��e=�E�=�D�=���=���=�I�=� >�J>*>^.>`>Ȑ�=�=�S�=�a�=$aZ=��<�<�OW�D�ʽ ����M�-���渗��䩾*}���   �   [��������|���؆���d�8,9�-x��ѽ����R��M#����TD.��[�<苽2���q�Ƚ
,޽[r�Q�彵�ֽr��ڽ��*Z_�g��:�X�<�w�<؅C=ҿ�=9:�=�
�=���=H��=H9�=���=a�>Ly>�*�=���=0&�=~��=���=h�T=���<h��=��n��|�	�R�9�$th��/:��˂���   �   �h��[I��f"��4d�Ī?��i��X�e^���oS���������¦���μ�7��H�����Ou��� �����Z!½MƸ�����	犽[U�ڄ�\ �����:�Ԗ<R�=P=��=Ԫ�=�&�=��=Ҍ�=RH�=>��=V�=ا�=�=�=���=uر=�0�=R�H=L��<�T��� ����tq!�A�I��Cm��|������   �   Vk���b��UP��5�m�����x5����Q��"�H�>���0� Cu� D����r��R༢�(��[_��Q��Dʕ�6���߿���ᐽXh����U�ԙ#�pTټ`�J���;p݋< =�^?=]y=Ǒ�=�I�=���=�>�=���=�@�=���=W��=�8�=l�=hǀ=p�3=���<@ ��q��&��#�ɽ��
�(��`E�	k[��zh��   �   �}6�[�-�(����fdԽ�ՙ��B�xU����@�0�2<0��<xѠ< �{<С�;�X��p���2�f�1���X��s�`��������y���g���L���*�'��a�����=�;��<�= UW=Z�=�̞=E��=�6�=��=ʪ�=�d�=��=�@�=t�X=\:=�'�<�hû̪����c��\��=W޽]������-��\6��   �   ���c�����׽���"��0�� rv�0c�;|m�<�	=&�!=fj$=P=l�<�܇<@�l;��#��5��&%��:�0\���u� ���g������A7����m�DK���H�ļ�6���<���<^\.=�Yg=���=���=Ȧ�=�2�=(Ҕ=g6�=0�Z=��"=�3�<���;hk:�����h$M�䕎��^�׽`��Pn��K��   �   P��q՛�}� �4��QǼ ���P�z<�1=Bp;=�:a=t=,t=*�b=�A=��=��< �< a˻���`���J��5~�7?���W��"���ˊ��x��������ڛ��}�2�4�ldǼ�Ѓ���z< +=Xj;=�5a=t=Ht=T�b=*�A=��=4�<H�<�˻`�� ���J�24~�t=��=U����k��������   �   ~�J���<�ļ����<�<�b.=l_g=Y�=�=	��=�4�=EԔ={8�=8�Z=ξ"=�:�<0��;pd:������%M�j�������݇׽̺��p��N����������׽+��j��R��p�v��*�;�`�<�	=Ư!=e$=�J=da�<�ч< Vl;�
$��?��4)�|:��\�l�u�-������(����3����m��   �   �S�����y�;�'�<��=[W=�\�=Ϟ=���=�8�=���=���=�f�=��=�B�=\�X=�<=�*�<�cû@����c�_��^Z޽._�;��h�-�`6�$�6���-�[�z���iԽ�ڙ��B�d���XA���2<��<�Ơ<0�{<pt�;P���l������1���X��s���������:�y��g�P�L���*�� ��   �   �1;��<�=hd?=|by=@��=.L�=���=�@�=V��=|B�=���=�=:�=��=lȀ=�3=@��<�"���r��(����ɽ۝�D�(�@cE�n[�>~h��k��b��XP��5���j�潐9����Q�(/��>��:1� �v��o��8�r��^���(��a_��T���̕�z�������㐽�h���U���#��Mټ��J��   �   Lܖ<n�=jP=� �=次=�(�=���=f��=�I�=���=VW�=���=�>�=���=Nٱ=61�="�H=p��<P\��� ��򜽈�6s!�s�I�NFm�~��0��<j���J���#���6d�?�?�l�`\佖a��*uS�¢�lɸ�H̦���μ�<���H�m���=x���#�������#½,ȸ������犽2[U��������$�:�   �   �|�<��C=W��=�;�=K�=���=���=p:�=���=��>�y>�+�=���=�&�=��=���=��T=��<P��V=�fp����	���9�vh�����p;�������������>~��چ�� e�.9��y�2ѽ:���R��Q#�����H.���[��ꋽ������Ƚ�.޽�t�e��f�ֽ��������Z_��f��:�h�<�   �   Fu=��e=�F�=�E�=���=���=�J�=!>/K>w>�.>H`>>��=t�="T�=�a�=aZ=��<�<�QW���ʽ���M�케������婾&~���V��@���<��$G��?��� S��$��;��7���܆���Z��O���e��$�����w�̽���� �����c����Ͻ�����l�L�� ��`
s<�   �   �%=֞x=hڠ=�B�=P��=�1�=�} >�>I
>��>y
>/j>b.�=��=|��=�W�=F�\=�k�<؊b��i���ؽ@�"��[��舾�Y������"��?\žT ��q����ա�������c�_�2�R��OWʽ������}�z�q�Ɛ���ҝ�~����(| �.,�3�B���W �|ݽ�q���)w��C
�М�\A�<�   �   �*=��~=H�=���=�:�=
��=�>h>
�>8�>�>f>�  >���=���=A�=�0]=@
�<��p���o���ݽ4P&���_���������rw��N+ž��ɾ@ž����Ty�����>Ci���7������ѽ�0���焽�e}�_���8?����Ž�n齆N�j����>��
K�b�ὌӲ��{����0���ٕ<�   �   � %=��x=�ڠ=�B�=|��=�1�=�} >��>)I
>��>"y
>Bj>�.�=��=Ќ�=,X�=��\=o�<�b�N�i���ؽ�"�2[�舾�X������!��*[žD���n����ԡ�������c��2�>��nUʽ𴙽��}�f�q�*���9ѝ��	����{ �+��1�1���V ��ݽ�o���&w�\A
�p��dD�<�   �   �w=B�e=�G�=&F�=���=���=�J�=!>CK>�>�.>f`>���=��=�T�=�b�=vcZ=$�<��;��KW�?�ʽ���j�M�d�������㩾%|���T��;���:��]E��u=���R���$��7���3��]ن���Z��O���e�^!��E����̽��꽾 ��������{�Ͻ���d�l�Լ�����s<�   �   ��<&�C=?=p<�=��=\��=���=�:�= ��=��>�y>�+�=���=t'�=貽=*��=��T=ĭ�<����=��k����	�J�9��qh���8��[���渦�5����{���׆�A�d�**9�av��ѽC��(R�BI#�j���?.�v�[��勽y�s�Ƚ�(޽�n�����ֽ���M���@S_�``���9�p�<�   �   ��<J�=�P=�!�=x��=6)�=5��=���=J�=ֶ�=�W�=^��=�?�=���=[ڱ=�2�=�H=��<$���� �휽_��n!�n�I��@m��z���
���f���G��� ���0d��?��g�oT佽Z��.iS� ��8���P���{μ2���H�,����q���������½����6����⊽`RU�V|������:�   �   @r;��<0=f?=�cy=���=�L�==��="A�=���=�B�=l��=V��=�:�=��=ʀ=V�3=觯<0卻�h�T"����ɽ8��ޓ(�$]E�fg[�2wh��k���b�RP���5�x��x���0����Q���`h>���0� �s� ��x�r�E�"�(��S_�4M���ŕ�D���κ���ܐ�c����U���#��@ټ��J��   �   �K����軠��;4+�<�=\W==]�=UϞ=п�=�8�=L��=��=3g�=\�=�C�=��X=6A=�6�<0%û8���`�c�AW��Q޽�Y�$����-�
Y6��y6���-���0��h^ԽyЙ�>
B�,E���~@���2<L��<pݠ<��{<���;���������1���X��s�ܫ��S����y�@�g�<�L�H�*����   �   ��J�����ļh���<��<�c.=�_g=��=\�=[��=i5�=�Ԕ=H9�=z�Z=��"=<C�<���;�F:������M�����촽�}׽E��j�H��������׽0��������Nv�`��;l{�<$	=.�!=Xp$=:V=Dy�<@�<�,m;��#�#�����:��\�r�u�צ�����N����0����m��   �   �}��!ԛ�*}���4��OǼ������z<:2=�p;=p;a=�t=�t=4�b=|�A=��=X��<��<P7˻��������J�`(~�27���N���鶽v��~���Tx���Λ�^�|�\�4��<Ǽ�A����z<9=�v;=�@a=�t=�t=�b=Z�A=r�=��<��<�˻\���|���J�T)~��8��Q�������M����   �   ���C�����׽���B��v���ov��f�;\n�<0	=��!=k$=�P=�n�<p��< �l;h�#��,��<��:��\���u�7���i��ܸ��}-���m��J��	���ļ���<�<pj.=fg=U�=��=���=�7�=�֔=e;�=��Z=��"=�J�< ��;�=:�ļ��M�+����ˀ׽h��m��J��   �   >}6���-���E��dԽ�ՙ�"B��T�� �@���2<��<�Ҡ<�{< ��;M��x���j���1���X���s�h���,���"�y���g��L���*���t>��P]�0��;�9�<=dbW=`�=�ў=&°=�:�=B��=�=i�=�=uE�=��X=�C=�:�<�ûX����c��X���S޽�[������-�"\6��   �   �k�d�b�UUP�³5�N��}��N5��J�Q�"� �>� �0��%u��?����r��P�
�(��Y_�&P��Pȕ���������ސ��c��B�U��#�|:ټx�J���;���<�=�k?=&iy=D��=�N�=X��=
C�=d��=nD�=���=͎�=H<�=��=.ˀ=F�3=l��<�⍻�i��#���ɽ����(��_E�Jj[�dzh��   �   |h��@I��R"���3d���?��i��X�D^��HoS�`��4�������Ԅμ7�*�H�����|t�����o���t½�ø������㊽�RU��{������:��<0�=�P=�#�=���=(+�=  �=R��=�K�=0��=�X�=���=�@�=���=X۱=�3�=b�H=l��<�%��F� �o~�jp!�b�I�Cm�N|��n���   �   A��������|���؆���d�,,9�"x�~ѽ�����R�nM#�j��D.���[��狽������ȽG+޽Rq�����ֽX��V���ZT_�x`���9���<(��<��C=�Ã=�=�=:�=���= ��=�;�=��=x�>Uz>�,�=���=:(�=���=ï�=ȰT=h��<h��=��l����	���9��sh��:�������   �   �U��A���;��MF��O>����R��$��9��p5��ۆ�Z��O���e��"�����Z�̽��꽢 �Ԃ����
�ｵ�Ͻ�����l�<������s<�x=ʋe=bH�=G�=���=���=�K�=�!>�K>�>
/>�`>��=d�=:U�=c�=�cZ=l$�<��;�zLW��ʽ���V�M� ��������䩾}���   �   �[ž��������ա�,���a�c���2�����Vʽٵ��0�}��q�珄��ѝ�n
���⽑{ ��+�d2����>W �[ݽ�p���'w��A
�0��D�<T!%=^�x=!۠=4C�=��=N2�=~ >,�>VI
>ͧ>Fy
>fj>�.�=<�=��=eX�=�\=�o�<��b���i��ؽf�"��[�^舾�X������-"���   �   ʎc��^�ʨN�r�7��C�" ���ͽ�^��|���e����=���˽�"�$��3H�>}j�Tg��/ǌ�U���Ì���h��A�|�}�ս���\���f8<:F)=��=E�=�~�=���=��>z]>&&>�W>�>(e><>.��=���=F��=9��=tMN=���<����0�t��6{���(�4��N��^��   �   2W^�t�X�I�I���2�����U����ƽ=Ϡ�����x[������O�ĽN>������C���d�a��������������XT���2c��=��
�vfѽNz���؇9<��'=��=�e�=\�=ظ�=ޙ >h;>�>�4>��
>�$>� >�2�=���=�)�=/��=K=��<0=������)���޽��� 1��I��*Y��   �   oSO��I�<�:�0�$��!�0L��̱�k����s�fyp�/���%�����LO�@B4�C�T�=o�ލ������=����p�cU��2�L��Ž��j�l{���s9<�h"=D��=ʒ�=���=���=2=�=��>��>�>�K>Y>���=��=��=�h�=g��=p@=�e�<�泻�k��D���zѽ�g	�?&���<�)�J��   �   �C8��.2� �#��]�Ӄ�I���1��d_�:���7���Y��Z��[a��[^���"�;�BT�#e���k��g��}X��T@��X!��p��-���V��ȝ��.<�L=�t=�&�=�R�=x��=�B�=h��=��>B�>�>���=���=���=D��=�Ȣ=4�~=&�,=��<`�λ�(�^���0���������"T)��95��   �   ������6�+@�-$��Ws��,O�������Xݼ�G�rUK�.̑���ƽ����U���1�0�A���H�nF��:��&�8�� �ݽr��<A��ʕ��=<X1=�X=#�=�!�=�W�=(��=zH�=��=���=��=���=B9�=Ze�=���=EN�=f�X=��=��^<0"�h<��0o��ʪ�8�ڽ����w��   �   F����|�	�νDU��wn��27����(�j������ջ��V�Nؼj�9�}�������y����X����"��D"�(��D��S?������Dg3�t����H;d}�<D�/= �t=�e�=�{�=�4�=t&�=��= ��=r>�=��=(Ͻ=���={!�=��c= �"=���<��;��u���DOa�m���h伽�4۽	�����   �   �d���v��Oƍ���Y�*f��8��`wH���<x`q<p�y<�/<����Ҕ�<<���r�����ɽҀ潨����������3���ƽ!~���`���43�l�ʼ bƻ��C<���<�7=��r=�=Ob�=��=H]�=�Կ=Pm�=Jo�=�s�=�Z�=lyT=��=���<��;H` �L�м�&��4b�md��ܣ�aص�����vg½�   �   ��V��' ��|¼������;Tf�<���<f�=*�=�I=��<��<p���ۼS9�`f~��|���{��7=��!ϻ�m���\��,=���'z�\�E��t��C����.<,��<��%=��Z=�T�=iL�=�>�=��=��=݈=Dih=��4=���<@bi<@u��t����~�:�)�
T�@�w������g���$����������   �   ��L�׼0�F���?;�'�<�=03=6�V=��j=(�l=��\=��;=8=�2�<��R;�\�����Y1�&J`�o���<댽3d��$����ׄ���n�2�K����׼�	G���?;4�<$�=�3=нV=��j=��l=�\=�~;=�1=�$�<�MR;0!\��Ｒa1�jQ`������팽�e��ꐒ��퍽�ք�P�n�N}K��   �    ;��0ś��/<P��<�%=��Z=LW�=�N�=�@�=o��=>�=�߈=�nh=��4=D��< }i<���������s�z�)��T�x�w�����xh���&��t!������������V�@/ ���¼ ,��P��; Z�<���<��=~�=D=�<�<0���-ۼ\9��o~�n������A��\һ����:^���=��\'z�<�E�Lq��   �   0Hƻ0�C<T��<z�7=�r=9�=ld�=�=V_�=�ֿ=po�=�q�='v�=X]�=�~T=�=\�< ��;xO ��м"�&��4b�e���ݣ��ڵ�����
k½�h���z��bʍ���Y��m��F����H���<xIq<0�y<@<@��`ᔼXD��r�]���ɽͅ�r���O��������6��ƽ]��;a���33�}ʼ�   �   ��H;��<��/=��t=�g�=�}�=J6�=$(�=P�=���=4@�=���=ѽ=���=�#�=Ȫc=��"=��< �;@�u�(�Pa�����Y漽87۽\�����^���ۀ�'�ν6Y��r���7����8�j���� �ջ��V�$[ؼ��9�����*���P�p������"��F"�*��F�eV�dA�����xg3�8���   �   �B<:3=l�X=W$�=#�=*Y�=���=�I�=f��=8��=,!�=T��=�:�=�f�=E��=�O�=0�X=ڜ=`�^<8��<�.2o�s̪�Z�ڽ|�����y�~����� 8��C轑'��qv���!O����ἬݼJM�z[K��ϑ�t�ƽ��������1���A���H�;pF��:���&�����ݽ�����=A�ʕ��   �   8.<,N=Rt=�'�=�S�=p��=�C�=b��=�>��>2>µ�=���=���=X��=�ɢ=��~=��,=D�<��λX)��^��#2��� �����U)��;5�4E8�Z02���#�<_���K���3��hh_�>
:� �7��Y�K]��0d���a���$�;�PT�8e���k��g�dX��U@��Y!��r��;���V�ɝ��   �   �t9<�i"=Ύ�=d��=:��=���=�=�=�>��>c�>KL>RY>T��=��=ľ�=<i�=嬋=�p@=df�<0鳻�l��E���{ѽ�h	� @&���<�]�J��TO��I�h�:�D�$��"��M�α�󴍽v!s�r|p�ܷ�������P��C4���T��>o�����nჾ���0�p�(dU���2��L�QŽ��j��{���   �   @�9<,�'=��=Nf�=l\�=(��=	� >�;>�>�4>��
>%>A� >
3�="��=(*�=_��=0K=��< @�����*���޽h��!1���I��+Y��W^��X��I�d�2�+��dV����ƽ�Ϡ�F���R\������\�Ľ�?��C���C���d�ra�����	������T��l3c�|�=�/��fѽ�z�����   �    h8<|F)=6��=E�=�~�=���=��>�]>(&>�W>�>#e>8>(��=���=0��=��=0MN=���<`õ������o{���>�4�N��^�ʎc��^���N�b�7��C�" �l�ͽ�^��|���n����=��8�˽�"�2$��3H�Z}j�]g��7ǌ�X���Ì�
��� h���A�_�L�ս����[���   �   8�9<��'=^ �=�f�=�\�=Z��=� >�;>�>�4>��
>#%>R� >:3�=\��=~*�=ς�=XK=��<�0��N���(���޽X�Q 1�\�I�*Y�rV^���X���I�%�2�	��TT��ΚƽPΠ������Z��ڵ����Ľj=����=C��d��`��0���4�������S��2c�:�=�
�eѽ�z�h���   �   h�9<l"=���=��=���=���=>�=5�>�>x�>_L>mY>���=��=1��=�i�=���=�r@=8l�<p˳��g��B��~xѽ�f	��=&�~�<���J��QO�q�I���:���$�� �J��ʱ�����Xs�Pvp�������(��AN�A4���T��;o�����߃�d��@�p�zaU���2��J��Ž�j� s���   �   �.<�Q=�t=�(�=^T�=���=FD�=���=6�>ի>M>��="��=J��=���=dʢ=N�~=��,=\�<0�λ�"��Z��S-��������$R)��75�zA8��,2�8�#��[����(F���.��X__��:�l�7��Y�cX���^��^[��!�0;�,T��e�d�k��}g�X{X�BR@�vV!��l�����V�,����   �   (Y<z7=��X=�%�=�#�=�Y�=���=J�=���=v��=t!�=���=(;�=ig�= ��=�P�=��X=��=�_<`��4��(o��ƪ���ڽ�����du�������3��;�S ���o���O�ԇ������ܼpB��OK��ȑ� �ƽ��������1�}�A���H�&kF��:�)�&���� �ݽ��4A�Ļ���   �   �%I;4��<��/="�t=�h�=`~�=�6�=�(�=��=���=~@�=J��=�ѽ=��=a$�= �c=��"=��<+�;@�u����Ea�g}��%߼�/۽~����ȸ��]w�	�ν�P��=j���7�̃��j��R��Vջ��V�Aؼ0�9�n���#���h
� ��\��}�"�rA"��$��A��M�+:��x����]3������   �    ƻ�C<X��<�7=��r=��=�d�=`�=�_�=׿=�o�=�q�=�v�=�]�=R�T=0�=��<���; : �Dwм��&�"*b��^��J֣��ҵ�ň���a½1_��q��%���<xY��]�@)���H���<Hyq<йy<�H<@���Ô��3���r�Y��L�ɽ�z�4���Q}��v���:-⽕�ƽx��$[���)3�Pmʼ�   �   D/��`���8"/<(��<ʨ%=4�Z=�W�=)O�=MA�=���=��=�߈=�oh=·4=t��<��i<@B��𫁼di��)��T�v�w�´���a�����������_@�V�� �<j¼ ����;Lt�<p��<v�=:�=:P=P(�<H�<P��d
ۼ�H9� [~��v��ru���6���Ȼ����2V���6���z���E��i��   �   ̒�0�׼(�F��@;+�<D�=3=��V=��j=��l=0�\=.�;=�8=�4�<`�R;��[����\V1��E`������猽�_�������獽�Є���n��qK�:��ԗ׼�F��y@;�7�<V�=� 3=P�V=Ȼj=��l=��\=�;=?=`B�<�QS;��[����nN1�>`�.����䌽�]�������獽nф���n�|vK��   �   �񀽚�V�% �,y¼ ���p��;�g�<���<ܘ=��=~J=�<p�<����ۼ|Q9�.d~�^{���y���:���˻��
��X���7���z�"�E��f��&��z���7/<@��<8�%=t�Z=JZ�=�Q�=�C�=��=��=��=<uh=��4=��<��i<�j��𞁼T]��z)��T��w�i���-b��9 ��I�������   �   c��(u��Bō�<�Y�e�H7��@mH���<0bq<�y<`1<���є��;��r����(�ɽ�����ځ��m���0�	�ƽ�y���[��~)3��iʼ� ƻ��C<���<r�7=L�r=�=g�=x�=�a�=ٿ=�q�=t�=�x�=o`�=��T=��=L�<��;( ��oм�&�()b�-_���ף��Ե�����
e½�   �   ͼ���{�?�ν�T��n���7���༐�j�p�@�ջx�V�\Mؼ�9�8���X�����������"��C"�'��C��P�,<������r^3������?I;��<��/=h�t==j�=��=|8�=3*�=F�=���=8B�=��=jӽ='��=y&�=F�c=�"=l�<�D�;��u�x��Ea�8~���༽�1۽���8���   �    ������5��?��#��s���O�>�����ݼ�G�&UK�̑�y�ƽv���#����1���A��H�lmF�+�:��&���K�ݽ`�>6A�`��� \<�8=��X=�&�=/%�=[�=<��=dK�=���=���=�"�=��=�<�=�h�=���=fR�=
 Y=J�=P
_<� ��4�^)o��Ǫ�|�ڽ��)��.w��   �   $C8�d.2���#��]�����H��1���c_��:���7�T�Y��Z��;a��8^���"��;�T��e�m�k��g�"}X��S@��W!�o�� ���V�����(.<pR=0t=�)�=6U�=���=2E�=���=��>R�>�>��=8��=l��=��=�ˢ=v�~=r�,=�<�λ�"�|[��b.����������S)�n95��   �   5SO���I��:��$��!�L��̱�[���js�Dyp�&���������BO�1B4�0�T��<o�̍����������p��bU���2�rK�'Ž��j��t��P�9<Xl"=
��=���=?��=r��=�>�=��>W�>Ƶ>�L>�Y>B��=��=���=�j�=n��=t@=�m�< ȳ�h�NC��Myѽ g	��>&�y�<���J��   �   W^�a�X�?�I���2����zU��қƽ7Ϡ�u���q[������M�ĽF>������C���d�a����������{���BT���2c���=��
��eѽ�z������9<z�'=p �=�f�=�\�=���==� >�;>>�4>	�
>O%>�� >�3�=���=�*�=5��=K=��<.��8��)��=޽��� 1�ڗI��*Y��   �   �"սK�νo���3��S8���ar���[���c����׶��$����+���b�����)���6ʾ���%�����Q��ǫ��kɾ���b`����S���*'�� r� �<�A3=.�=�H�=�Y�=���=z�>1)
>.v>�
>�p>� >h�=|��=4��=IR�=�ԇ=|F=h
�<`��;�w���`�p�Ӟ��gO��<�ν�   �   Z=Ͻv�Ƚ�������D����f���P�z%X���~��W7��)'�*(]�8N��1^����ž�Dܾ�����ﾟ���9ܾ�mž����T���:O�*��8�������[<`4=5��=d�=��=�=��>�	>�9
>M�>��>�=)�= ��=p]�=�
�=�у=vr?=h��<�'�;��|�,���-m��t��	����ɽ�   �   M^��̴��~˥�]	��h�m���E��0�&�6��b��1���-ݽ����L�D���\_�����g�ξ��ܾ���#ݾ�cϾ`鹾 ʞ�Ko��4iB��)�sӝ�|�h 3<"6=<M�=���=�	�=�'�=E>D�>�u>}`>��=���=,"�=���=? �=s�=��n=�{)=�h�< (b;�'�����80c�!����ӫ��Ӻ��   �   �ڤ�'R������T~f�	8����ܘ��^���*�~&z�-���(�T�3���g��?������,��|Ǿ-�˾��Ǿ)����&�������g�X/� �Ǌ�(�ļ�]<�7=�\�=b�=��=�x�=��=�" >* >��=B.�=R��=D��=0�=�I�=&�=�6C=x:=`�v< ���M��,����V��R��r��������   �   ���Ɗs�N�M��� �H���]����l��2���Ƽ^o*���� �ѽ�^�q�A�*q��K��������S���3��4���R���hy�b\I�����Yν�]i������<�v4=���=@B�=%��=>|�=�N�=J��=�[�=���=�C�=��=���=��=
�u=Tn<=�=�;�<�R&;�B�ܳӼ�&���M�04s�<ͅ�E6���   �   ��K��}+����t������ (��`�y;`�M; ���e��b�,��'����ݽ0t��q@�MJf�(���5��ߦ��?���SK���]s�\;P�:O(��H��\����H>���Q��(�<>�*=��=�,�=��=���=T��=h��=���=��=4��=7T�=OS�=(�U=ւ=4;<�_<�0u�����l�ڼ�����5��O�Xm`�?f�t�_��   �   ��� h˼�;Y� 3���6<d��<蚼<���<���<���;`/w�$~&�u����jֽ- ��J.�PI���[��d�*�b�XW�v�B�c'��.�ͽ�"���D��#"��w<V3=T�b=O�=�T�=��=���=��=
Ƶ=2 �=_�=��h=Z(*=x�<8x<��ѻ�a��d����(��1E�2X�Z�a���b��h[�D2K���1��   �   x鼼� � )o;���<���<.�=�,=&�.=�=x=�<�C<��Ʊ��������!Y�j%�����(�,�)��"��/���^�ֽ�����ig���Ho(�8�*<pK�<�9=��p= l�=��=\`�=.�=��=�x= �@=���<0�?<������ټ�~2�:1l�񇋽�ؘ�!��\���ɓ�P_���i��`@�l���   �   h�o�`�
;8#�<t= �6=V]=n�t=^e{=��n= N=$�=���< �������?��/��gʴ�pYӽ����Z6� �۽��Ľ*���{��hvI�dy��o�@�
; �<(p=ތ6=�\=��t=�`{=��n=LN=|�=8w�< ���&!?��5���д��_ӽ/���`��;�m�۽&�Ľ�,���|��^wI��x��   �   �k(���*<�P�<H�9=X�p=�m�= �=vb�=��=/�=�y=��@=���<��?<@���Ъټ�s2�`&l����� Ԙ�������Ǔ��]����i�a@�>��X＼�� � �n;ȏ�<\��<t�=,= �.=(=�0�<��B<H��j����������_�)����&)���)�#��2�����ֽ���lg�&��   �   $"�X�w<25=��b=��=&V�=��=R��=��=Fȵ=�"�=6�=.�h=�/*=P)�<0�<�Nѻ�P����@�(��+E�T�W��a�@�b��h[��3K���1�����p˼�NY��϶��"<d��<���<�<y�<�ȋ;HMw�ֆ&��Ƒ��pֽw�ZN.�.I���[��d���b��W�m�B�oe'�����ͽU$��<F��   �   ��Q�t)�<h�*=��=�-�=��=��=҇�=��=���=�=���=�V�=7V�=l�U=r�=�ھ<Xz<`�t��z����ڼ���0�5���O�xn`��Af��_���K�x�+����t����� ƀ�`Ly; SM;P䌻�q����,�,����ݽw��t@��Mf����7��਑�*���M���`s��=P�6Q(��K��L����J>��   �   H�����<�w4=��=C�=��=F}�=�O�=���=*]�=|��=�E�=��=���=�=�u=ds<=�=�D�< �&;x�B�H�Ӽ&���M��5s��΅�8�����R�s�
�M�z� ����g���l��E�4�Ƽ6u*�����ѽFa�.B�-q�~M�������«��T���5��ܽ�����*ky�R^I�(���[ν�_i��   �   \�ļx]< 7=�\�=��=���=�y�=t�=$# >� >��=�/�=���=��=��=�K�=��=:C=t==��v<`���K��D����V��S������T����ܤ�)T������Z�f�
8�n������T��d�*�f+z���L*�W�3��g�A��u����-��Ǿ��˾"�Ǿ����(��"���4�g��/���Ȋ��   �   �3<P6=M�=Z��=�	�=4(�=�>��>v>�`>���=���=2#�=���=V!�=��=��n=\})=Tk�<�4b;,'����>1c������ԫ�պ��_��J��� ͥ��
��B�m���E��0��6�&�b�~3���/ݽق���L�$�]`��6�����ξ��ܾ2��%ݾ�dϾE깾�ʞ��o��jB�,*�9ԝ��   �   ����[<�4=^��=Rd�=��=H�=	�>�	>�9
>~�>��>��=�)�=x��=�]�=l�=�у=*s?=`��<)�;X�|����x.m�<u�����D�ɽ>Ͻ?�Ƚ�������D��(�f�.�P�'X��������8���)'�)]��N���^��w�žZEܾk��^��3��d:ܾ4nž��������O�n�������   �   �q���<B3=L�=�H�=�Y�=���=}�>4)
>2v>�
>�p>� >\�=n��=(��=8R�=�ԇ=�{F=�	�<���;w�t����p�����O��T�ν�"սN�νo���3��N8���ar���[���c����?׶��$����+�+�b����)���6ʾ���0�����N�ﾾ���kɾ���L`��ʀS�����&���   �   L��Pc< 4=ޑ�=�d�=4�=~�=�>�	>�9
>��>��>��=�)�=���=(^�=��=Y҃=(t?=���< 6�;X�|�>���+m��s������v�ɽJ<Ͻg�Ƚ������C���f�6�P�$X�W ������6���('��']��M���]��b�ž,Dܾ.�������;9ܾ%mž���΍��PO�^��ݤ���   �   d� .3<6=uN�=��=v
�=�(�=�>��>*v>�`> ��=ބ�=j#�=��=�!�=�=D�n=L)=Lp�<�fb;x��z���+c������ѫ��Ѻ�.\�������ɥ����
�m��E��0�R�6�.�b�$0���+ݽ�����L������^��(���S�ξf�ܾ��᾿"ݾ�bϾA蹾�Ȟ�`n���gB�*(�ѝ��   �   �ļ�!]<�#7=X^�=��=b��=z�=��=I# >� >�=�/�=
��=+��=O�=L�=��=<C= @=��v< Q�<A�������V��O��K����~���פ�GO��C���Lyf�n8�:������b����*�"z����'���3���g��>�����}*���Ǿ��˾��Ǿ����W%������ �g� /�0�BĊ��   �   @����<|4=���=4D�=��=�}�=P�=��=j]�=���=�E�=(�=(��=��=`�u=4u<=Z�=K�<��&;ȗB���Ӽt���M�,s�EɅ�a2�������s���M��� ����hS����l����Ƽ�i*�� ��^�ѽ�\���A�'q�J��N���(���Q���1��B���|��Wey�WYI���)UνrUi��   �   ��Q��6�<T�*=O�=�.�=��=���=J��=b��=ҥ�=F�=Μ�=$W�=�V�=��U=�=�޾<��<��t��q��H�ڼ��� �5��O��c`��5f���_�.�K��u+�@�����������~���y; �M; ����X��|�,��#���ݽjq�Zn@��Ff�.����2���������5I���Ys��7P��K(��B��"���\?>��   �   h "�P�w<::=\�b=�=W�=*�=ʂ�=��=�ȵ= #�=�=��h=b0*=�+�<�<@>ѻ(K�������(��%E�`�W�̻a���b�
^[�(K��1���� W˼ Y��M���P<���<���<8�<x��<0�;�w��u&�����eֽ���G.�LI�k�[���d���b�W�W�B�&_'�����ͽ���:��   �   �I(��+<lZ�<��9=��p=�n�=� �=�b�=��=x�=ty=J�@=��<��?< ����ټr2��#l����Ҙ�*�����+Ó�/Y��x�i��U@�T���ּ��� ���o;(��<���<V�=�,=��.=�=8J�<1C<0��L�����F�R�!����C�(���)���"��+��
�T�ֽ����D^g�&��   �   @�o��;�+�<Fw=H�6=�]=��t=4f{=n�n=�N=��=���< F������?��.���ɴ�TXӽd��Y�'4��۽1�Ľ&���v��JlI��n�0�o�@D;x2�<�z=H�6=,	]= �t=�j{=^�n=&#N=�=�< ���轼d
?�)��Pô��Qӽ��S.�^�۽o�ĽH#��4u���jI��n��   �   �ۼ�p� � fo;P��<���<��=�,=��.=X=x>�<XC<0��R��Z��)����X�%������(�b�)� �"��.�8�ضֽ����ag�<�H(��+<_�<��9=0�p=�p�=��=�d�=�=��=	y=��@=���<(@<�O���ټ\g2�l��{��͘�������W���SW����i��U@�����   �   L��\_˼�.Y��鵺�<<���<���<���<���<���;�-w��}&�D����jֽ ��J.�I�U�[���d���b��W�q�B��a'�����ͽ���<��"���w<�;=|�b=O�=�X�=��=���=��=�ʵ=`%�=5��=�h=d7*=�:�<h�<��л�9������(�0E���W���a���b��][�()K���1��   �   "�K�Xz+�&��ؚ����� �� �y;@�M;@���ld���,��'����ݽt�lq@�*Jf�����4���������K��]s�b:P�N(�F��t���NB>�p�Q�\6�<�*= �=�/�=�=���=���=��=���==	�=��=�Y�=xY�=��U=��=��<@�<`-t� f����ڼ ����5�@�O�td`��7f���_��   �   ���0�s�z�M�p� �\�缐\����l�01�`�Ƽ"o*������ѽ�^�b�A��)q��K����������R���3��������hy��[I�����Wν�Xi����4 �<$|4=��=�D�=���=�~�=&Q�=��=�^�=F��=�G�=&�=^��=���=z�u=jz<=t�=�T�<@';�B�ԞӼ@���M�^-s�sʅ�4���   �   �٤�?Q��V���h}f�d8���8��� ����*�\&z����(�I�3���g��?��􀦾�+��qǾ�˾~�Ǿ����&��ۑ����g��/�w��Ŋ��ļ�]<�#7=�^�=B�=���=�z�=��=�# >E >:�=1�=x��=Ƣ�=��=�M�=��=�?C=xC=P�v<�-�\>��n��
�V��P��z�������   �   �]��?���˥�	�� �m���E��0���6��b��1���-ݽ����L�A���Y_�����a�ξ��ܾ����#ݾ�cϾA鹾�ɞ�o���hB�)�eҝ����)3<�6=zN�=9��=�
�=�(�=�>��>}v>Na>���=΅�=t$�=A��=�"�=L�=��n=n�)=�s�< }b;���D��v,c�����oҫ��Һ��   �   �<Ͻ2�Ƚ��������C����f���P�d%X�� ��y��V7��)'�$(]�4N��.^����ž�Dܾ��꾼�ﾗ���9ܾ�mž����>���O�������z��h`<�4=͑�=�d�=J�=��=1�>�	>:
>��> �>��=0*�=8��=�^�=S�=�҃=Lu?=���<�<�;0�|�
���+m��s��n ���ɽ�   �   8#ҼH�Ǽ����"���̓��`��b=��^�N����	��H�a���X��i�pZ
�
d�-0��;�z�>�m ;�40���	�I㾠���ł���/�S�ʽ�2�(�/<�J=�g�=+��=���=v^ >t�>�8>\�>�>�8�=���=:��=���=[u�=��=�0v=lB=2=�*�<pf<�i8���N�숣� nǼ�   �   ��Ǽܠ���f���9��<	������$���LUS�����F����C�3������be����N��,�9�7��3;�*�7�L�,�b��e�޾�r�����9�+��Ž|��(�A<>;L=���=�O�=���=T�=�>��>}�>�
�=&[�=�e�=���=��=�Ϥ=~F�=8|i=�6=r=��<��;�Jl���Q�0���h���   �   t���-���o��77��
%�xZ]�кü��2�� ��AF��4���|����.�Ӿ�K���\�Y#�TO-�.�0��j-�XD#�'n�����Ҿ~$���p����u����; �H�s<�R=�=���=0@�=���=>e>�=xP�=���=��=�n�=�|�=ہ�=��q=4qB=��=���<�hY<@:>;��̻Љ_�ܚ���r���   �   �߁���@� v��0���l�`cl��T����t�4�ͽf4�Ɵ_�Xƕ�[R��2}��k�(��Nj�}� ����Bm����zP�GW���?��4�W�� �ț�R���W�<�Y=���=m��=0��=@��=�N�=B��=���=|��=���=@E�=��=�ƅ=��Z=(�+=��<,��<�2< H;�̯���<�\5��`���Ҕ��   �   �9,��k����;���;h-<��< !�:�Tt�T�%�p�������:��M~��H���Ǿ���l� ��I	�#d�7�	�������&�ɾ�����q��N9����{��h��C�<d�`=�ʟ=���=l��=�-�=h��=
r�=���=TԽ=Jv�=�0�=��`=h)=|��<軆<�4�;@�,�X"��5u��P��X+������(���5���   �   0�ɻ��H;(vA<(s�<G�<��<��<�vd;�Z���JM��������OK�Bބ��ϣ�㿾�{־�^�2�j���{پ�ľ�ਾ�C���VU�@�Y��ZH;�P{����<��c=�h�=k�=~��=��=���=d��=䑮=��=f'm=N�*=���<�< ���h\����� ���
?"����W���8z����u��   �   �ك�Xy<�ϧ<x��<$V=�=|�	=l}�<���;$�����g�LʽM�t�J�)�~��ꖾ���>Ŷ��������p����l���v��]?]���)���P%�������cd;��=na=S�=��=�z�=4+�=f��=�R�=o��=�C=l��<���;8DY�t*�z�M�{���"{��\�����������I�����c��A3�p���|���   �   �է� H<���<�!=��C=t:S=�xL=�y,=@��<���;���	i��Ž�Z�P�7���^��8~��艾B����(��7���Jq�?�O��b)�L1�XR���R��Y����<�.=��U=9_�=eX�=�y�=���=(v�=�Ag=6�=t=�<���v�
��w� ����ؽ���������b����O?ѽ�`��ꃽ<�4�tZż�   �   �g$��L<p�=Z�@=^�m=c�=&,�=0�v=�#J=�=f"<3��L�I�5m������D�/��EB�0xK�s�J��@A�i�/�ף�����N^��Z�����a$�`�L<h�=~�@=Ȅm=~a�=,*�=~�v=<J=�=hD"<PG��Z�I�>t������!�0��JB�}K�"K�@EA�6�/�������%b�������   �   T^��x�<�.=��U=9`�=�Y�=�{�=͈�=�x�=�Gg=��=$O�<�Z�`�
�4�v�o����ؽ�{������i_����:ѽ�\��烽^�4�pVżpѧ�H|H<��<|�!=��C=�6S=|tL=�t,=���<��;L��$i�xŽ�^���7���^�*>~��뉾	����+������iNq���O��e)��3��U��`�R��   �   ܞ��`Kd;|�=a=��=	�=@|�=�,�=���=�U�=���=@C=��<�9�;�Y��b�M�̡���t�����߂�����J���طc��=3��������`݃��s<P˧<ȯ�<�R=�=�	=�r�<`Ô;�ʳ���g��Qʽ�P���J��~�^햾~��6ȶ�����������<o���x���B]��)�X��'���   �   �K;��������<�c=bi�=�k�=���={��=���=���=~��=��=z.m=f�*=���<��<����G��P��j�����7"�<���S�p��w��ȍu�@�ɻ��H;�kA<�l�< @�<0��<���<�"d;dg���RM����v���RK�Y���$ң��忾i~־�a�2�N�澕~پ ľ�⨾4E��>YU�B��[���   �   `{��h�B�<L�`=˟=:��=H��=�.�=���=�s�=���=�ֽ=y�=4�=��`=�&)=���<pˆ<pq�;@g,��	�@!u� I���%����������`6��x?,�p|����;`��;-<ء<���:0ht�0�%��s��������:��P~��J��Ǿ���� �_K	��e���	�в�%���ɾ���s���O9�����   �   �ɛ��U��V�<�Y=.��=���=���=��=�O�=v��=���=0��=���=�G�=b�=nɅ=2�Z=��+=t��<԰�<`2< ~;���P|<�4������Ԕ��⁼��@��� E0���m���l��#T�D'���t�C�ͽL6�"�_��Ǖ�T��!��l�N��k��� ����Qn����R羜X���@��ȟW���   �   |����< ���s<�R=<�=���=�@�=P��=�>de>�=�Q�=Ι�=X��=p�=�~�=���=H�q=ttB=��=���<�pY<�P>;��̻H�_������t������00���o��?7� %��c]���ü��2�����H�d�4���|�2���t�ӾTM���]�0#�4P-��0��k-�E#��n�����Ҿ;%���p�x���   �   Ž����A<R;L=���=�O�="��=��=�>��>��>h�=�[�=tf�=���=^�=UФ=GG�=�}i=b�6=�=$�<��;�Gl�h�Q�聠�Di��<�Ǽ�����h���;�����(������WS�Е�����رC�������� f�W��"O���,���7�E4;���7���,���I���޾Ps������+��   �   ��ʽ22��/<VJ=�g�=D��=���=�^ >z�>�8>`�>��>�8�=���=2��=���=Qu�=��=�0v=�kB=�=@*�<Pe<�m8�x�N�X���tnǼd#Ҽx�Ǽ����"���̓��`���=�h�^�bN����	�S�H�����w���澀Z
�d�-0�;�z�>�k ;�,0����	��H���eł���/��   �   DŽ6����A<�<L=8��=;P�=d��=��=(�>��>��>x�=�[�=�f�=���=��=�Ф=�G�=f~i=D�6=�=��<@�;�)l�H�Q��}���d��t�Ǽ�����c���6�����4�������TS��������C�輇�����dᾥ��YN���,��7�]3;���7���,�������޾^r��P��Z�+��   �   ����7 ���s<ZR=0�=���=A�=���=�>ye>0�=�Q�=���=���=Qp�=�~�=���=@�q=�uB=^�=ܽ�<�zY<@�>;�̻�y_�L����k����&�� o�-7�� %��P]�ܵü��2�f����D��4�n�|�J���,�Ӿ�J��\��#��N-�U�0�j-��C#�^m�|����Ҿj#���p�9���   �   �ě��G��p`�<��Y=���=���=t��=���=�O�=���=,��=\��=Ć�=�G�=��=�Ʌ=0�Z=�+=��<D��<�)2<�;���Xi<�X)��(��HȔ��Ձ���@��T���/�� l��+l�PT�d����t���ͽ�2�ҝ_�"ŕ��P��z{��j���(i�O� �[��l�����N羐U��[>��ěW�����   �   �{�xh��N�<Ғ`=�̟=Z��=��="/�=.��=�s�=.��=�ֽ=Dy�=T4�=x�`=�')=@��<�Ά<���;�<,�(���u�4?�����į���s���'��� ,�0>���%;p��;@,-<��<���:�At���%��l������|�:��J~�G���Ǿ.��"� ��H	��b���	�2��Y��ֻɾ|���p��!K9�N���   �   �?;��@��X��<� d=$k�=!m�=|��=��=���=���=�=��=�.m=�*=��<@�<���(D����弒|����F3"��{�XM���h���mu�lɻ I;�A<~�<0Q�<��<��< �d;�N���CM�c�������KK�S܄�zͣ��࿾�x־�[�!�Z���xپ�ľ6ި�PA���RU��<��S���   �   ą����d;v�=(#a=⁓=T
�= }�=�-�=���=�U�=ه�=�C=��<�=�;8Y�2�(�M�����ps�������������������c��63�0���\���@���h�<�ܧ<(��<�[==ȸ	=���<@)�;H����g��Fʽ�I���J���~�!薾����<¶��񻾮��u���j��^t���:]���)������   �   4F���<�5=мU=�a�=�Z�=z|�=a��=y�=8Hg= �=P�<�W�ڲ
���v�����ؽ{��+��l ��^���ｕ7ѽ�Y���ヽ�4��Fż �����H<��<�!=4�C=�?S= ~L=v,=���<��;l���n�h�y�Ľ�V���7���^�p3~��剾R���&��c���Dq�\�O�8^)�x-��K���~R��   �   �;$�`M<��=̎@=��m=9d�=�,�=@�v=�$J=D=�g"<82���I�m��g��W��/�~EB��wK���J�3@A�|�/�������S[�������C$� M<0�=T�@=ʌm=�e�=�.�=��v=�)J=�!=І"<d���|I�Xf������h�/��@B��rK�!�J��;A��}/�N��f���W�������   �    ���P�H<\��<Ĝ!=n�C=d<S=$zL=�z,=���<`��;���i��Ž�Z�3�7�|�^��8~��艾����(��ꁅ�AIq�K�O�va)�0�|O��܃R�\L���<d5=��U=�b�=*\�=~�=J��=j{�=�Mg=��=�`�<p�Z�
�h�v�����ؽ�r����r���Z�
��
2ѽ�U�������}4��Aż�   �   �����<�ا<��<hX=h=��	=�~�<@��;X�����g��Kʽ�L�a�J��~��ꖾ���%Ŷ��������2����l���v��u>]�|�)�5ｿ"������`�d;��=f#a=k��=>�=`~�=,/�=�=HX�=���=�C=���< ��;X�X� �@�M�N����l��O���6{����Q�����c��13�P��������   �   prɻ�I;��A<Tx�<�J�<� �<L�<@�d;�Y���JM�����z��OK�<ބ��ϣ�㿾z{־�^��K�澹{پ_ľnਾ+C���UU�2?�W���C;�`V�����<� d=jk�=�m�=n��=U��=���=���="��=��=�5m=��*=���<��<�P��D/�� �强r�����+"��u��H�8��(e�� lu��   �   H%,�@M����;���;�-<X�<�4�:�Rt�
�%��o��j���ٟ:��M~��H���Ǿ���j� ��I	�d�.�	�~������ɾC����q��WM9���ｎ{�ȃh�<K�<&�`=�̟=���=���=0�=`��=�u�=��=ٽ=�{�=Z7�=8�`=�.)=���<dކ<��;��+����P�t�D6��������r��@(���   �   �؁���@��f⻀0���l��Xl��T�\����t��ͽ^4���_�Sƕ�XR��/}��k�&��Kj�{� ����9m����YP�W���?����W�l ��ƛ�M��]�<��Y=r��=���=���=(��=�P�=���=���=��=���=�I�=
�=q̅=��Z=��+=��<���<<2< �;0���ha<�L'������ɔ��   �   �𪼬)���o�X47�P%��X]�8�üX�2�� ��2F��4���|����-�Ӿ�K���\�X#�UO-�-�0��j-�TD#� n������Ҿ`$��Ip�`������(: ���s<�R=
�=���=FA�=��=3>�e>�=�R�=8��=��=�q�=���=���=��q=ByB=��=���<��Y<��>;Р̻xw_�\����l���   �   ��Ǽ���|e���8�����D�������0US�����D����C�0������ae����N��,�9�7��3;�)�7�J�,�_���Z�޾�r������+�RŽ���h�A<<L=��=6P�=t��=��=E�>"�>��>��=|\�=:g�=���=`�=nѤ=sH�=,�i=��6==P�<$�;� l��Q��}��e���   �   �-�<��<8�<辘<P�<���V+�
�������S�aq���Ծ*X
�{B,��WM�n�j�������S7��=�����גj���L� +�����kξ_��� <�,�̽ �8ҙ<4,l=�̯=
��=���=��=�� >:��=]�=��=4�=C�=zò=WM�=�y�=nO{=��[=�?=�%=T�=�q�<x�<�0�< T�<�   �   �o�<���<���<8��<��3< L��jk�%W������N�C�����ϾI��r�(���I���f���}��3��?��5��p�}��cf���H���'����aPʾz���7��Kƽ�����l�<�ln=�=��=���= 6�=n��=�H�=P��=֭�=���=��=��=��=��=�]h=D�I=0o.=�z=�`=8�<�A�<d�<0b�<�   �   \��<0�<���<��<(L|< ��8μh'�����r?�_ጾ��¾�D���h��p>�{.Z�e(p��M~�z����j~�Mp�r9Z��;>�6�����Ao������_�*��]���aϼ���<�t=l��=T�=���=�^�=Bn�=v��=��=�V�=�l�=`-�=>Ύ=��t=VCO=�V.=�W=��<���<�+�<�~�<ྣ<���<ٳ<�   �   �,�<�"�<hF�<�I�<�?�<p�<@sj��OI�P�Ƚ��&��Pz�tƮ�0q�{���"-���F��[��?h�	�l��~h�d�[��3G��l-�xx�N�8��e4p�|���֘�\e��t��<�(}=�M�=��=���=���=���=R,�=.��=,d�=�e�=��r=,q@= =���<pL�<�G<��<p?�;���;���;�*<H�f<�<�   �   �ߪ<X��<�= h=��<�
�< ��L� �W����zqR�}i���ƾy6���-�M.�]@��.L�`hP�l�L�kA�O	/���������Ǿh┾3sM�2J���vm�P�ƻ.�=�ق=h�=���=d��=�b�=/��=拴=��=�y=Z�8=lQ�<�`< <z9�?.�|����*�� <ż�9���蔼��E��S��@{x;�qL<�   �   tb�<��<rp=�}$=�x =�W =�v<Ћ7�0H�
qʽ�p%�-�q������оR����K��#"�gt,��80�-�JA#����<, ��=Ծ-զ�!Zv�\�&��SĽz#��h�;�#=υ=@O�=�)�=��=�'�=�]�=�K�=|�K=l�<Л<��C�� � vD��w�xꋽ{���= �������V�>�#���ռ�6>�`�-;�   �   ���;X��<�!=��8=�'C=�1=���<�"<⮼1���	�1V6���}������ɾ���j���������S��W�Qﾮ Ͼ;���W)��HB�U �Z5��db��<߂<�+8=L8�=�1�=��=*��=��=�Rt=�%=��<���@���+�����߅⽢� ����~�	��#�_��ɽ�����c��B���C��   �    ^��<2�<XL=�;F=�a=��_=�?=t[�<��;`�漈3������:v6���s��˗�e岾	�Ⱦ�"׾�ܾYUپ	�̾��
�������29J���T&��`44�p꺻���<B�E=�=�&�=�@�=���=4\]=j=(l<8x���j�z������5&��A��vT��c]���[���O�(�;�Hg �$��G��(
~�P{��   �   �8�����;�<=j�J=b�w=k��=z=z�L=p��<I�;���6����^���$��iT�]�����˜��ʡ�����9����􇾘�i�&->����ɽ��m��/��0�;�==0�J=��w= ��=<z=X�L=���<��;�������f���$�koT�\c�>��>Ϝ��Ρ�j���l���������i�F1>���
ɽ��m��   �   �94������<��E=��=�'�=YB�=���=b]=$=0�<�`���j�*������0&�_�A��pT��]]�·[�x�O�V{;�"c �� �yB��~��u��A���5�<�L= ;F=�a=��_=��?= P�<��;L�漅9��d����z6�$�s��Η��貾ԳȾ�&׾�ܾ6Yپ��̾Z��ۤ��>ゾ�<J�ʎ�q*���   �   z8��`j���ڂ<4+8=�8�=X2�=D�=��=5�=�Xt=�%=@��<������#��q����|�Ҧ � ��ڤ	�>����}ɽ(��(~c��<���C�P��;8��<x!=��8=z%C=ķ1=|}�< �"<x�+���c"�*Z6���}������ɾ���o���������U��Y��TﾴϾ¨��[+��`B�� ��   �   WĽ� #��T�; �#=%υ=�O�=�*�=]�=�)�=`�=7O�=f�K=4�<��<@TC�T{ ��gD��w�㋽H}����������V��#�8�ռ�$>�@.;Xe�<���<�o=|$=v =NT =��v<��7��	H�vʽ�s%�,�q� ����о�����M��%"��v,��:0�-�7C#�b���- �<@Ծ7צ�B]v�� '��   �   4M���zm� �ƻ
�=�ق=��=���=���=�d�=6��=j��=��=Z�y=��8=Td�<H�`< ��9�.�(���,��|(ż`(��,ڔ��mE��/����x;�xL<�<���<�=\f=ܲ�<��< ��ܓ ��r�vtR�]k��XǾ89���/� .��^@��0L�WjP�T�L�2A��
/������x�Ǿ�㔾XuM��   �   ���xؘ�Ti��l��<P(}=&N�=z�=z��=��=��=&.�=i��=�f�=�h�=b s=�x@=�=`��<(\�<�8G<�<po�;���;`�;8*<�f<(�<-�<�!�<8D�<hF�<P;�<��<��j�\TI�e�Ƚ��&�Sz�Ȯ�.s澩��B$-��F��[�ZAh���l�z�h��[�5G�(n-�sy��O�m��)6p��   �   6�*�_��(dϼT��<�t=���=��=4��=�_�=>o�=���=���=yX�=�n�=�/�=�Ў=޸t=\HO=�[.=x\=p��<���<�1�<���<P£<���<ڳ<D��<�.�<���<x��< E|< |�8�μ,)���� ?�Z⌾��¾HF���i��q>��/Z��)p�O~�����k~�&Np�d:Z�S<>����2���p��(����   �   O�7�Lƽ\����l�<�ln=4�=X��=��=�6�=���=.I�=��=���=���=��=��=�=�=�_h=��I="q.=D|=6b=,:�<�B�<$��<db�<<o�<���<l��<���<��3<`V��m�;X�������N�������Ͼ�����(�:�I�R�f�8�}��3���� 6����}�df�a�H��'�����Pʾ���   �   � <�ǅ̽~�ә<�,l=�̯=,��=���=��=�� >H��=(]�=��=>�=C�=vò=RM�=�y�=VO{=��[=^?=�%=�=dq�<$�<|0�<�S�<x-�<d�<�ߺ<���<(�<@�ﻼ+�W���6��;�S��q���ԾCX
��B,��WM���j��������T7��<��� ��Ȓj���L��+�����kξ:���   �   �7�;Jƽ���Hp�<nn=��=���=L��=�6�=��=@I�=��=Į�=���=��=��=+�=8�=Z`h=�I=�q.=}=@c=�<�<tE�<��<\e�<Tr�<0��<���<L��<��3<`D��lj��V�����2�N�������Ͼ��!�(�B�I�=�f��}�E3�������5��Ӓ}��bf�p�H�L�'�+���Oʾ���   �   ڣ*��[�� Zϼlž<l�t=l��=L�=���=`�=lo�=���=���=�X�=�n�=�/�=�Ў=P�t=�HO=�\.=|]=��<��<�5�<$��<Lǣ<��<�߳<p��<d5�<d��<�ž<�T|<  �8�μ&����a?�������¾�C��h�&p>��-Z�V'p��L~�䜁��i~��Kp�_8Z��:>�Y������n�������   �   p���Ә�h[��h��<�+}=dO�=N�=��=t��=L��=X.�=���=�f�=�h�=� s=�x@=X	=���<D^�<X>G<0�<���;���;p�;�$*<8�f<@��<�5�<�*�<�M�<LP�<�E�<  <xej��KI���Ƚ��&�uNz�!Ů��o�x��!-�F�F�u[�>h�g�l�@}h�ӄ[�K2G��k-�Ow�L徛���1p��   �   XE���nm� Uƻ�=�ۂ=8�=� �=1��=�d�=���=���=5��=��y=�8=e�<X�`< �9�.��������P$ż4#���Ӕ�`_E�P����x;P�L<X�<���<F=Jl=Ŀ�<��<���H� �<���&��nR��g���ƾ4���,��.�M[@�-L�lfP�{�L��A��/������C�Ǿ����$pM��   �   �NĽ#����;��#={х=dQ�=�+�=�=@*�=n`�=yO�=��K=��< �<�RC��z ��fD��w�V⋽k|��y����6�V��#�8�ռ@>��l.;�p�<@��<�u=��$=<} =Z\ =��v<�t7�>�G��lʽ�m%���q�T���f�о/����I��!"�Wr,��60��
-�C?#�����* ��:Ծ�Ҧ�Vv��&��   �   �/���P����<�18=�:�=�3�=a�=ř�=��=�Yt=j�%=��<���2���#��3���=|⽖� ����n�	���A���ɽ1���yc��7���C��&�;4��<�'=J�8=�,C=�1=4��<�"<lӮ��}��D�R6�+�}�Z���a�ɾ\��q��p�g���Q��U�EM�C�ξ@����&��	B�� ��   �   t)4�0���<��<��E=��=.)�=jC�=���=c]=�$= �<`����j������m0&�:�A�hpT��]]�`�[���O��z;�Xb ���]@��d�}��p����lA�<�R=xAF=�a=��_=@�?=�g�<pV�;x���-�������q6���s��ȗ��ᲾN�Ⱦ�׾�ܾSQپ*�̾��ɞ��ނ�W4J�������   �   ���pF�;&E=l�J=��w=���=�z=��L= ��<PM�; �����m^���$��iT�]�����˜��ʡ�Ҩ��������i�W,>�����ɽ�m�|%��`+�;�C= �J=��w=���=@z=L�L=��<���;��ԍ���V�=�$�fdT��V����-Ȝ�Vǡ�^��������񇾰�i��'>�O����Ƚ��m��   �   0���4F�<�S=AF=da=`�_=��?=�]�<p"�;`��X3������-v6���s��˗�]岾��Ⱦ�"׾�ܾ:Uپ��̾�����������d8J�
��R$��04�`ź�P��<��E= �=�)�=�D�=���=Jh]=r+=�<PJ��\�j���2��J+&��A��jT��W]���[�x�O��u;� ^ ���:����}�2j��   �    ?�;(��<�'=^�8=�*C=@�1=T��<��"<�஼������ V6���}�
�����ɾ���e���������S��W��P�v Ͼ����)���B�� ��3���Z����<�08=�:�=�4�=q�=c��=��=p_t=��%=P
�<P������ƛ�� s�ҡ ������	�H�H���ɽn ���pc��0�X�C��   �   tt�<���<~u=V�$=${ =tY =@�v<�7��H��pʽ�p%� �q������оO����K��#"�dt,��80��-�?A#����(, �=Ծ�Ԧ��Yv���&�`RĽX#����;��#=0х=�Q�=�,�=_��=,�=�b�=xR�=6�K=�&�<��<�"C��m ��XD�,�w��ڋ� u����������V�T�#���ռ��=�@�.;�   �   ��<���<�=�j=���<�<�r�ҍ �,����nqR�xi���ƾv6���-�N.�]@��.L�`hP�i�L�dA�G	/�������i�Ǿ3┾�rM�I��,tm�@pƻ�=Pۂ=R�=8�="��=Nf�=V��=���=��=��y=�8=lw�<��`< U�9 �-�,�������ż���<Ĕ��EE��画�,y;@�L<�   �   �6�<0*�<�K�<�M�<�B�<�< qj�8OI�+�Ƚ��&�}Pz�pƮ�.q�y���"-���F��[��?h��l��~h�b�[��3G��l-�nx��M���4p����՘��a�����<�*}=SO�=��=���=l��=���=0�=���=ni�=�k�=Ls=,�@==���<<n�< ]G<�	<p��;�'�; ?�;x2*<`�f<���<�   �   ��<�4�< ��<�þ<hO|< �8`μB'�����n?�[ጾ��¾�D���h��p>�{.Z�f(p��M~�z����j~�Mp�o9Z�};>�/�����.o��s���%�*�s]��_ϼD¾<��t=N��=j�=���=�`�=Bp�=���=���=0Z�=�p�=�1�=ӎ=D�t=
NO=�a.=fb=H��<T��<�<�<���<|ˣ<襧<x�<�   �   �r�<���<4��<\��<��3<�I��:k�W������N�C�����ϾH��r�(���I���f���}��3��@��5��p�}��cf���H���'����WPʾm��7�gKƽh���,n�<\mn=��=���=h��=�6�=p��=�I�=���=���=|��=��=�=f�=|�=�bh=x�I= t.=*=e=P?�<�G�<x��<Xf�<�   �   �NZ=$�U=ģB=��=��<��$���Z�����J��ܜ�Ut����nWE�?Ts�GՏ��u���겿ZԼ��?���м�ײ�@��0p���r�ޠC����[1۾~���\5��6�������<� �=j_�=2��=`�=���=p�=���=t��=��=���=�:�=�I�=zpu=^=��L=�{A=h�;=XQ;=��>=��E=�N=#V=�   �   B]V=*bT=$dC=��=�G�<����O���^�E��Y����ܾ[���A��n�TK�������گ������㢹�:ӯ��z��������m��@�����־]����0� :��T����=읊= ��=Z��=�=Q�=���=^!�=a�=�"�=0	�=Ƈ�=�y=��[=X+D=�3=��)=k&=��(=8//=�9=b�D=��O=�   �   ��I=�?O=l	E=D�#=��<�5�v}0���ͽ��6��*��|PϾ-L���6�4"b�Nꅿ+d��e���XO��.����b��_���i���Ʌ�oza���5�?��Eʾ!��M�#��ߛ�p�G�:h=�+�=��=�C�=���=�{�=���=by�=���=I[�=$��=v�U=�S-=�=Ȕ�<8��<���<��<(��<؇�<)=�'=��:=�   �   ��2=��D=$�E=.�.=��<ֵ;M�������G�`�~�UL��[���;7&�"N�ݼt�����������7Ȥ��᡿F��w����u��N��%��r�����n�s�N������@)��(\ =��=*U�=�M�=��=>��=|�=�>�=�Q�=��O=�=(^�<�"%<��`:`O��@q��`C�`�a� m(;��(< 2�<X7�<Z	=�   �   �P=�1=0nB="B:=��=`��<`�������ҍ��_V�����{nݾ9���4�4SW� v�q=�����#摿�W��s����w�*3X��T5�3@���ܾ�㝾QO��K콆�>�PV�;��3=Ȏ=*�=�V�=�=��=���=��^=h�==�<�1��𖶼<���\G�vxa���f���X�N�8���
��\�������<�y�<�   �   �I�<*	=�8=�B=No,=�#�<��C:�n�E���M)�%��������� 6�d�P�Gf���s���x�
{t��2g�:R�7��X� i��ez��,-����&�⳽�輘r�<(�F=ؙ�=0�=���=0$�=8�=�&4=le�<�����	�ko�(q���Uҽ������������ҽ�����ـ��$�d����^;�   �   �g;I�<T�#=��D=��C=ʲ=���< .h��t�f��jE�����p��`!��"I���)���;���G���K��GH�m:=��+�]o������ľ𒾩}K����0�t�0�'��9�<J�U=@�=˞�=���=$Ve=��=h�'<�߬���e�� ��G���V%�w@���R��N[��X��"L��6��=����m���=Y�����   �   l#���z<x=�==%U="F=J�= �"<�ּs�������P��=��M��������y��y0������dA�h>�`�辏s��I喾N�]�p��:���l� ��;ز=61^=P�=@�}=^�S=��=`;X����V��d ��*�,���]��1����������}���N ���W���Gp�tlB�x����ȽH1g��   �   v�J���!��q�<�,=�/^=�;h=�[J=��=`_�;�����`	�� H�Ԅ����������9پ���Z��©�Jݾ��ǾHW��R���|Z�'����ǽ��J�H�!��w�<*�,=/^=�9h=�WJ=һ=��;���3&���d	�H�kׄ���������>پ̙�9���vNݾ��Ǿ�Z���T��f�Z���\�ǽ�   �   M?��xr�Pe�;:�=J1^=#�=��}=j�S=��=�;�����N�������,�@�]�8.���������	��|��������T���Ap�vgB�p��}�Ƚ(g����X�<�=r�==�#U=LF=��=��"<P�ּ�旽����P��@�� ����<����+3�������C��@�X���v���疾��]����   �   q����t�H(��5�<��U=A�=��=���= \e=��=X�'<xƬ�^�e�������P%��p@�c�R��G[���X��L�n�6��8�҆�`g���3Y� ����lg;<O�<��#=r�D=��C=��=ȴ�<HJh�j#t����@nE�x���s��Q%��kK�Y�)�|�;�{�G���K�eJH�==�R�+�vq�������ľP��K��   �   ��&�`峽L��n�<~�F=1��=1�=4��=�&�=��=�.4=�y�<@]��B���Zo��g���Kҽ}ｲ����������O�ѽK����Ӏ��$��v�� i^;Q�<:=�8=Z�B=Hm,= �<�PB:�u�����)�CÁ��������6���P�f�j�s�s�x��}t�O5g�r<R��7��Z��k���|���.���   �   <SO��N�h�>��D�;��3=KȎ=�*�=�W�=��=�=җ�=��^=��=�R�< Ά�P{��p���MG�ia���f��vX���8���
�$J���ּ�x�<���<,S=f�1=TnB=&A:=r�=��<�����������bV�����qݾ�����4�TUW�k"v��>��"��r瑿Y�������w�5X�gV5��A���ܾ�坾�   �   @�s��������7��j[ =��=�U�=�N�=Q�=��=�~�=vA�=�T�=�P=�=�q�<�L%< xc:0������`��`a���(;�)<X<�<?�<=��2=��D=�E=�.=8��<`��;\U���ī��I��~�N�������8&��#N���t������������Pɤ�	㡿G��]���$u�BN�&�%�At��]����   �   �!���#������G��g=�+�=u��=@D�=���=�|�=��=;{�=8��=�]�=���=��U=PZ-=��=d��<\��<��<�*�<���<̏�<N,=B'=^�:=d�I=�?O=	E=Z�#=ط�< >5���0�2�ͽ~�6��+���QϾ M���6�e#b��ꅿ�d��-���$P�������c����Ij��ʅ�Z{a�k�5�Ӎ��Eʾ�   �   Y]��ԡ0�q:�������= ��=>��=���=��=�Q�=N��=J"�=0b�=$�=�
�=H��=H�y=�[=�.D=�3=x�)=�m&=��(=1/=	9=f�D=6�O=�]V=(bT=�cC=�=�E�<`���O�f��O�E��Z����ܾ�����A���n��K��렠�aۯ�����m��G����ӯ�K{�����:�m�@�W��8�־�   �   S���5�Q6��������<�=�_�=T��=z�=���=|�=���=���=��=���=�:�=�I�=fpu=�^=��L=V{A=8�;= Q;=��>=d�E=�N=�"V=|NZ=��U=��B=��=��<�$�`�Z��
�J��ܜ��t�����WE�aTs�WՏ��u���겿`Լ��?���м�ײ�@��#p���r���C�x��'1۾�   �   �\����0��8����H�=���=���=���=��=�Q�=d��=Z"�=<b�=($�=�
�=V��=h�y=.�[=�.D=V�3=��)="n&=X�(=�1/=�	9=L�D=:�O=�^V=bcT=8eC=��=LI�<8�� �O�n����E��Y��i�ܾ����A���n�K��3����گ������ ��y����ү��z��c���&�m�7@�����־�   �    ��˦#�xݛ���G�k=-�=:��=�D�=���=
}�=,��=X{�=L��=�]�=��=ؙU=�Z-=�=L��<���<���<�,�<��<���<�-='=J�:=��I=>BO=�E=J�#=���< �4�{0�o�ͽ��6��)���OϾ�K���6�F!b��酿�c���󦿚N��j���/b������h���ȅ�Iya���5�q���Cʾ�   �   ΄s�N~�z�����_ =��=�V�=MO�=��=S��=�~�=�A�=U�=�P=�=r�<�M%< �c:P���0�������`� );x)<�@�<�C�<�=��2=�D=��E=<�.=��<P�;�E������8F�R�~��J������6&�� N�G�t��~���������$Ǥ��ࡿ�D������u�cN���%�np��h����   �   �MO�?G�R�>�0��;0�3=(ʎ=,�=�X�=j�=e�=��=Զ^=
�=TS�<�̆��z��$��&MG�jha��f�juX��8���
��E��P���(�<��<�V=B�1=�rB= F:=`�=|��<�惼������]V�	���Plݾ���>�4�FQW��v�@<������䑿�V��6���Mw�1X��R5��>�E�ܾ�᝾�   �   1�&��ܳ���(�<|�F=A��=x2�=��=*'�=T�=D/4=�z�<p[��
��LZo��g���Kҽ@�W���q�����v�ѽA���|Ҁ��$��p����^;�X�<~=\!8=ԑB=�s,=H-�< �D:�g� �|)�L����ﶾ�������5��P��f���s���x�>xt�0g��7R��|7��V��e���w��+���   �   �����t� �'�0G�<
�U=)C�=���=}��=6]e=t�=0�'<�Ŭ�(�e��������P%��p@�F�R��G[�\�X��L��6�18�����e��l0Y���`�g;�W�<��#= �D=��C=�=<ʓ< h��t����JfE�c���m������F�d�)��;�ՆG���K��DH��7=�d�+�m����p�ľ[풾XyK��   �   J4��$b� ��;��=<7^=/�=D�}=.�S=��=��;����N�������,�7�]�3.���������	��b���e���`T��uAp��fB�ƹ���Ƚ�$g����<D$=��==Z*U=jF=0�=�"<�}ּ�ڗ�H��u�P��:�����y�⾌������-�%��E��>��;����o�� ▾$�]�L��   �   b�J���!�̇�<�-= 5^=�?h=6^J=T�=g�;������_	�� H�Ԅ����������9پ��O����Iݾr�ǾW���Q��|Z�~��V�ǽD�J�@�!�\��<" -=5^=&Ah=~aJ=h�=ࠟ;L������[	�`�G�ф�9���j���n5پ2��t����XEݾF�ǾbS���N���vZ�t�0�ǽ�   �   d ��x�<'=��==�)U=XF=n�=��"<l�ּ0�������P��=��K��������z��v0������XA�W>�7��]s��喾��]���b9��:i� ��;B�=�6^=��=��}=��S=$ = X�;�����G����;�,��]��*��������~��T��������P��@;p��aB�x��:�Ƚhg��   �   �h;D_�<x�#=l�D=��C=��=4<�)h�"t�0���iE�����p��]!��!I���)���;���G���K��GH�f:=��+�Mo������ľ�$}K�q��t�t���'�TA�<��U=eC�=���=J��=�be=��=�(<(�����e������� K%�zj@���R�.A[���X�bL�Z6�63�}�
_���%Y��Ẽ�   �   \a�<*=�"8=��B=�r,= (�< �C:�m����:)���������� 6�e�P�If���s���x�{t��2g�:R��~7��X��h��:z���,���&��೽Է輤x�<��F=>��=*3�=x��=?)�=,�=�64=���<`���8��bJo��^��Bҽ�w��Q���c���ѽ�����ˀ�j�$��_���_;�   �   �Y=�1=8sB=�E:=�=��<TR�������_V�����xnݾ8���4�4SW� v�r=�����$摿�W��s����w�#3X��T5�&@���ܾ�㝾�PO�$K콖�>��h�;x�3=�Ɏ=n,�=�Y�=��=�	�=�=&�^=��=dh�<�k���_������=G��Xa���f�gX��8�j�
�2��Ё����<,��<�   �   ��2=�D=̰E=��.=���<pߵ;�K�������G�W�~�RL��Z���;7&�"N�ݼt�����������9Ȥ��᡿F��v����u��N�	�%�~r�����2�s����������>^ =>�=�V�=�O�=��=��=��=BD�=;X�=�P=�=@��<�v%<�Ef:P������P�滀_`� �);�9)<�K�<�L�<�=�   �   ��I=�BO=�E=��#=D��<�5�}0���ͽ�6��*��zPϾ,L���6�5"b�Mꅿ,d��f���YO��0����b��a���i���Ʌ�lza���5�9���Dʾ!���#�Lߛ��G��i=�,�=@��=E�=���=~�=���=}�=Z��=M`�=І�=��U=&a-=�=��<�<h��<�8�<p��<d��<t1=�'=T�:=�   �   l_V=�cT=ReC=t�=�H�<0����O����Y�E��Y����ܾZ���A��n�TK�������گ������䢹�9ӯ��z��������m��@�����־]��q�0��9��<��<�=U��=���=��=�=LR�=��=*#�=9c�=N%�=��=Ҋ�=��y=��[=82D=��3=�)=q&=�(=�3/=�9=��D=L�O=�   �   _b�=�H�=��n=-=}<�Zռ�����.�����~zܾ���7Q�?����/������3�ؿ�k�/������*���M�Nؿ�����a��M�����N��D���վ*���4����� �9�%;=+\�=�=�=D{�=p�=+��=r��=*�=�=�4t= R=8�7=�}&= �=\S =�**=|�:=P�O=�g=xc}=h}�=�   �   ���=. �=PQm=v/=4�<سļV����P*��K��_�׾��WM�e,���\���L����Կ�{�?��i������o��Կػ�è��_?��;K��e�=�Ѿc������R}�� �:�V==Nћ=w
�=P|�=J`�=�P�=,s�=Ԙ�=}9�=�t�=zhV=�!2=Tu=��=���<"=�w=1!=j�9=X�T=�n=��=�   �   Tx=ֳ|=�h=�<3=��<8���B��|��ڳ���ʾ�D�6B��x��%���۲��rʿ;ݿV�|@�,�[3ݿ�zʿ���W���.w��Q@���r2žU�{�*�@�^�@c�;�2C=���=ت�=��=���=C޻=֧=]��=~�e=�m.=�X�<=�<�3A<��;`�;�<P~U<�Х<�[�<>:=��B=0�b=�   �   ��O=�7d=�_=*�7=d��<�b�Xw����2�k��������~0�>�b�"H���������8;˿.\ֿ�Jڿՙֿa�˿�P���B���<���Ab�$q/�S ��౾1|`��?�Z0� |A<��J=��=�i�=��=G�=�=��w=n3=7�<���;@��p��Z��M�������#ȼ`%U� ��9�pr<�.�<4)=�   �   �=t">=h�M=�-:=�o�< 4�:ʖ/�wlڽv�E�����U⾑,��@G���u��4������x���Β��*¿�꾿9��і��U���cov�:|G�������Ee��u�=��Ľ������<l�Q=��=�f�=d�=���=��L=��<Ps�; D��Zo2�Q��������=Ž5\ѽ�PϽ��Q������d+�����:85�<�   �   `sy<;=�j1=��6=R�=`�Z<�����ƞ��4��o}��<���� ��(�#vP��ww��������'�������I죿de��R⍿�'y���Q��)�B���v����{�r��̐��	\����<U=��=ը�=�j=8&=$@�<�L���9�Lţ�y%���� 4-�OQ>���E�e�B�YJ6��>!�Z��O�̽�v��Ri�@!��   �   G� Kr<Ԗ=��*=�%!= ��<�l�h}B��n޽^�@�MĒ���;�����)��sJ�P�g����	���ʉ�\{��nM��V�i��L�1�+�V	�_�оh֔��
C�/j޽ �7�@I�:n�=^�Q=�jg=�N=*�=p,<,Ҽٷ��>��:�"�+�R�k�}�������G��|���m6��Ʉ���a�:�4�!�{����w>��   �   ��?�� U�<4�=4�)=��=px<�3���������>W������Ͼ���"Z�j]6��wI���U���Z�*�V�j*K���8��� ��'���Ծ`���"_�p������է�@��<��=||E=��:=(��<н�;�����F�����ҬF��-��DX��O��d�ؾ���e����>Tܾ��ƾ}��^ԋ��W����x����   �   U���T�� g�:�K�<��(=V/=>=0�<$��	j��R���6Y�G㕾���[뾱��@���!�^w%���"�e��v�OC��Ǿf���z?f��9�Ś��������:HP�<��(= /=�=�<p��p�����f<Y��敾���`�~��G��4�!��z%��"�[��(!�H��Ǿ�����Df�{=��   �   5s�����ৼ���<�=�}E=\�:=,��<p�;�}��+?������F�/*��T��MJ��;�ؾt��������5Oܾ��ƾx
���Ћ�PW��������>�?����l\�<��=t�)=Џ=��w<�C��F�����WW������Ͼ���\��`6�.{I�K�U�C�Z���V��-K���8�W� ��)�'�Ծ>�Z&_��   �   C��n޽��7�@��:d�=Z�Q=�mg=вN=l�=�S<d�Ѽ����A��D�"�F�R���}����,����B��)���Z2��hń�D�a���4���l����l>���F��^r<��=��*=�$!=D��< kl��B��t޽~�@�ǒ�U�;ڋ�B�)��vJ���g�#�����̉�+}��$O��v�i�ȢL���+��W	�g�о�ؔ��   �   �{����ϐ�8\�<��<�U=��=Ϊ�=��j=*&=�T�<�WL���9�����������--��J>���E���B�D6�69!�R����̽�o��^^�8 �Ȋy<�>=�l1=��6=��= �Z<`ȿ��ʞ��7��s}��?��� ��
(��xP��zw�U��M�������ǵ��g���㍿^*y�$�Q��)���x���   �   �f����=�԰Ľ0����<~�Q=M �=h�=���=���=��L=���<�ҿ;�'��:_2�b���񞫽�3ŽRѽ�FϽ����XI��ʳ�*X+�٤���:�A�<=%>=��M=�-:=�k�<���:t�/��pڽ\�E����^X�9.��BG��u�6��������x����+¿�쾿���3�������}qv��}G��������   �   �᱾�}`��A��\0�hwA<��J=M�=k�=k�=0I�=��=��w=�3=K�<�	�; ���U��X���>�0y����@ȼ��T� X�9�r<:�<~)=��O=d9d= _=~�7=���<p�
]w������k�d��ǌ�9�0���b�'I����������<˿�]ֿ_Lڿ.�ֿ��˿�Q���C��}=��Cb�@r/�,��   �   B3žt�{�����^�p]�;�2C=���=���=*��=:��= �=bا=!��=� f=u.=�h�<N�<WA< b�;�]�;��<0�U<ޥ<�f�<�>=>�B=��b=�Ux=̴|=�h=�;3=ر�<����C�����Ҵ��=�ʾ�E�KB��x��&���ܲ��sʿ;ݿ\�A�-�A4ݿe{ʿȮ���/w��R@�s��   �   ��Ѿ�������}����:�V==�ћ=�
�=�|�=a�=�Q�=Wt�=0��=;�=�v�=dlV=�%2=�y=8�=��<=,{=,4!=�9=t�T=��n=/�=㩇=L �=6Qm=�/=��<L�ļ�����Q*�EL��1�׾R��WM��,��J]��pM��O�Կ|�����i��P��&p�v�ԿVػ�	����?���K�.f��   �   ��վ������R��� X9n&;=\\�=>�=.�=f{�=��=<��=���=9�=)�=�4t=*R=8�7=�}&=�=0S =^**=<�:=(�O=�g=Dc}=D}�=Bb�=�H�=h�n=Z�-=�}< \ռH��2�.�ٚ���zܾ��8Q�T���0������C�ؿ�k쿈/������*���M�Nؿ�����a��9�����N�yD��   �   v�Ѿʯ������ }��A�:.X==қ=4�=}�=*a�=�Q�=^t�=8��=;�=�v�=llV=�%2=�y=V�=p��<8=r{=�4!=��9=��T=T�n=��=H��=� �=ZRm=P/=��<@�ļװ���P*�mK���׾���VM�,,���\���L��f�Կ{�����h��H��-o迒�Կ�׻�X���?���K�qe��   �   )1žl�{�����^� ~�;x5C=���=&��=���=t��=D�=zا=0��=� f=*u.=�h�<LN�<�WA<�c�; `�;H�<P�U<tߥ<�h�<�?=b�B=4�b=dWx=��|=0�h=�>3=���<�����@�����8����ʾYD�kB��~x�`%��=۲��qʿWݿa�}?�+�e2ݿ�yʿC��������,w��P@���   �   ߱��y`��;�~T0��A<��J=��=�k�=��=�I�=�=�w="3=0K�<P
�;����U��"���>��x����
ȼ��T� ��9��r<L=�<T)=��O=�;d=._=P�7=���<�T��Sw�u��D�k�Z����}0���b�CG����������9˿�Zֿ�Iڿv�ֿ�˿}O���A���;���?b��o/�:� ��   �   Mc����=���ĽT�켬�< �Q=�!�=i�=?��=���= �L=(��<0Կ;�'��4_2�_���잫��3Ž�QѽiFϽE����H������V+��դ�@\�:�E�<�=(>=2�M=2:=�w�<@��:\�/��hڽ�E�B���S�'+��>G�a�u��3��1�򄴿3���j(¿G龿���W�������
mv�<zG��������   �   ��{�H��ǐ���[� ��<�U=��=㫆=$�j=�&=�U�<pVL���9�껣�������--�J>���E���B��C6��8!������̽o��@\������y<B=�p1=��6=2�=`�Z<$�����2�l}�q:��B� ��(��sP�1uw�-��㬚�d���'���}ꣿ�c�������$y�J�Q��)�����s���   �   �C��c޽�7� C�:�=~�Q=Lqg=�N=��=8W<|�Ѽ����5��B�"�C�R���}����*����B�����F2��Iń���a�X�4�2�]���~j>���F�Hlr<��=ĺ*=P+!=h��< �k�uB�Ei޽��@�������;���N�)��pJ�2�g�2�~����ȉ��y���K���i��L���+��S	�ޢо�Ӕ��   �   l�K����§�Ɓ<p�=�E=��:=d��<��;X|���>�������F�.*��T��NJ��;�ؾr�������"Oܾ�ƾU
���Ћ��W���������?�0��0d�<��= �)=��=hx<�"��A���8���W����'�Ͼ`~�{W�lZ6��tI�U�U�/�Z���V�'K�s�8��� �1%�l�Ծ����_��   �   O������#�:�_�<��(=�/=B=�<��輷i��:���6Y�E㕾���[뾳��B��	�!�^w%���"�_��l�0C��Ǿ8���?f� 9���������m�:`Y�<��(=@ /=�!=��<0�輊c����01Y��ߕ����IV����M���!�-t%���"�\����=>񾫊Ǿ�����9f��4��   �   }?����tm�<ؕ=0�)=��=�x<P0��#������+W������Ͼ���!Z�k]6��wI���U���Z�)�V�e*K���8��� ��'�[�Ծ2����!_��o�P����ϧ�\��<�=��E=z�:=���< K�;�f���7��c���F��&���O���E��0ؾ��u��]��Jܾ.�ƾ%��;͋�W�l�������   �   8�F���r<*�=>�*=�*!=���<@�k�|B�fn޽E�@�FĒ���;�����)��sJ�R�g����	���ʉ�]{��lM��Q�i���L�%�+� V	�<�о<֔�a
C�,i޽h�7� ��:��=��Q=Zsg= �N=�=�z<��Ѽ����x佘�"���R�8�}����Փ��">������ .��z���8�a���4�r
�Κ���^>��   �   `�y<�F=s1=��6=j�=@�Z<L���)ƞ��4��o}��<���� ��(�$vP��ww��������)�������I죿ee��P⍿�'y���Q��)�5��cv��h�{���ː���[�L��<,U=Q�=s��=(�j=&=�h�<@&L���9����`����&'-��C>���E���B�t=6�3!�����̽�g��pP�H���   �   �#=V+>=�M=�2:=v�<@t�:��/�lڽ^�E�����U⾐,��@G���u��4������x���ϒ��*¿�꾿9��Ж��S���_ov�4|G����s��&e��(�=�R�Ľ��켄��<Z�Q=2"�=(j�=��=�=>�L=��<�.�;����O2�����t����)Ž�Gѽm<Ͻ¢��%@��
��bI+����� x�:�S�<�   �   8�O=2>d=V_=t�7=���<]�,Ww�����k��������~0�?�b�#H���������:;˿/\ֿ�Jڿՙֿ`�˿�P���B���<���Ab�q/�K ��౾�{`�%?�X0�`�A<��J=��=�l�=B�=zK�=��=�x=*#3=`^�< b�;��� ;��6s��0��j���� �Ǽ��T� ��9�r<�I�<,#)=�   �   �Yx=�|=�h=�>3=ط�<|����A��h��ճ���ʾ�D�6B��x��%���۲��rʿ=ݿW�}@�,�[3ݿ�zʿ���V���.w��Q@���d2ž6�{���H�^��m�;�4C=���=���=W��=���=��=�ڧ=���=f=,|.=<x�<_�<�zA<0��;��;�<��U<|�<�t�<�D=n�B=F�b=�   �   䪇=5!�=�Rm=~/=��<�ļ6����P*��K��_�׾��WM�e,���\���L����Կ�{�@��i������o��Կ ػ�è��^?��9K��e�6�ѾZ�������}���:vW==�ћ=T�=m}�=�a�=�R�=bu�=s��=�<�=8x�=.pV=*2=�}=��=��<l=L=8!=r�9=��T=^�n=\�=�   �   �I�=�{�=P^s=,,=�f,;<DS�;E��su�@�ž�+�C�M��H��4^���ѿP��L�	������Ш!�h��*k�h�	�|�9�Ͽ� ��H͆���J�u	��o���lg���뽆�����<B�q=�ܧ=�ٿ=�^�=��=*g�=�(�=�4�=tV=��)=��=4S�<((�<$��<4��<t��<r�=TP>=kc=�ւ=�ɏ=�   �   � �=S!�=�Zp=��=��x;��I��l�׫o������H�<�I��ۅ�@g��ܓͿ~?�2���������������"l�Փ�ӕ̿-��#~����F��O�����bb�ּ�����2�<��p=���=���=�H�=�ط=V4�=�Ɏ=�Ti= �4=��=���<�_�<0+J<PH<h@|<D�<Pi�<�!"=��K=��r=�p�=�   �   �=���=|�f=$U=��;$�.�,����^��������w�>��}�ɠ��_ÿ_w�h� ����.U�
�.m������ �o5�:�¿,퟿F�{��c<�Zc��6��ӶR�.ѽHV߼C�<��m=J?�=Pޮ=���=�6�=w�=�R=VW=\*�<@
�; ���|y�t���L<���h�Ѐ���ϲ;�d�<�o=�?8=N�c=�   �   n1G=(�^=­T=�=��@<�[��Zʽ��D�梾G���hc-�n�g�lJ���h���ҿA��h��l�L�
������o���[ҿ�Y��$풿�Vf���+����ɉ����:�D�������<�e=�[�={��=��=��i=�O#=�K�<���̌üjX1���q��֎���������6�Z�f��4��@Ƚ:Xa�<�=�   �   �]�<��'=�7=�:=)�<t������$�$��^�Ծ�g�~yK����O�������#ӿ�t濵��ۃ��p���K�bԿKt�� }��6���0K����~Ҿ�"���t����XP�l��<��W=�{=:�p=��>=��<@�:ༀ~m��>��ɯ�5/�D)��t!�n�����������ͽ������3�h䃼��<�   �    ؍9'�<L�=��=d��<��껔O`�����`a�x����E��Ĵ+�:]��ԇ�h��k����jƿu_ѿU]տ��ѿlǿ����g1������r*^�,F,��j�����]��D��ȣE�@�:�D=��?=RPD=��=�X�<x_��2M�j�����	�u�4���[�"{�����$���߀��^e���@�����ٽ����t,��   �   \����<��̝<��< n�<��;̏ �帳�j *��e����ɾ��
��4���^�����W���ä�[��ٍ��G����ѥ�����d��y>a�f�5����˾�*����)���(��b1<��=�=<t�<(r<Tھ�.��V���{2���o�������.�ƾ5վ�ھL�־�/ʾݵ��ٛ���|�W\@�*�
梽�   �   � ���k� 6��и�<��<���<Ѐ�\W��>�2�H�l<��}վ�"��/�=�P�o��u���8��}���ȋ��{���q���S��1��z�B�ؾ�I��=M�L
�\�PG����<D��<�2�<�n�;��Ѽ�N������M�Ǖ��N����$��K����`����2J��M����_t��&͔�ȕY��Z��   �   B^�B:���˼�b�;0��<�h�<@�!<H姼D8�����MmU����¶ξ,����ތ5���H�*U�D�Y�KV��J�=8�t �����5Ծ��`.^��Z�:5��|t˼P|�;���< d�< �!<H���}>��8��sU�K��T�ξ�����i�5�p�H�&U�M�Y�@V���J��8�w ���3:ԾW��q3^��   �   &AM����\�W����<L��<p;�<��;X�Ѽ�G��� �d�M�瑎�vI��R��������r	��F��J�d���o���ɔ��Y�<V�����c� ���p��<P��<H��<0���W��E�
�H��?���	վJ%��/���P��o��w���:������ʋ��}����q��S���1��|���ؾ�L���   �   -���*����(��@[1<��=\�=��<�<$¾�3��,�｢u2�H�o�F�������ƾ�վ?�ھ��־�*ʾTص��՛�n�|�~V@���ߢ�B~� <��ԝ<��<�k�<��;�� ����.$*�9h��.�ɾ/�
�y4���^�����Y���Ť�� ��%��������ӥ�����f��qAa���5�����˾�   �   ����]��H��X�E� ��:�D=��?=�TD=� =�k�<pE_��"M�����ʂ	���4� �[��{�9뇾N��۝���ڀ�:We�Z�@����{ٽ�󆽨� Ǒ9�1�<"�=Z�=��<�뻖V`�*���7a����GI����+��]�sև�<��o���mƿ�aѿ�_տ��ѿ(nǿ����3��m����,^�H,�xm���   �   �Ҿ@$��fv�?���XX�8��<8�W=n�{=��p=��>=�2�<@��:��߼�lm��4�����)��"�n!����������ܲͽw�
�3��΃�`<�i�<X�'=�7=�:=<%�<���y��� $��%����ԾCi��{K�,���	��C����%ӿ�v�������w��M�Կ�u��m~��7���2K�K���   �   2 �ኞ��:������������<.�e=�\�=eØ=��=��i=6X#=�`�<�-��pü�H1�ʺq��͎�����G啽e����Z���������:�p�<�=�5G=��^=֮T=2=�@<t_��]ʽ��D�袾s����d-�8�g��K���i���ҿ�B�i��m�.�
���j�����]ҿ�Z���Wf��+��   �   �c��7����R�N	ѽPX߼�B�<��m=@�=�߮=���=�8�=E!�=t
R=@_=T<�<�Y�;�2�pPy����l&����g��4��@�;s�<�u=�D8=��c=��=���=��f=�T=��;6�.���콚�^�߶�������>�\�}��ɠ��`ÿpx� � �V���U��
��m�X��)� �L6���¿�퟿8�{�Kd<��   �   �O������b�'�����2�<p�p=��=h��=�I�=�ٷ=�5�=vˎ=�Xi=~�4=��= ��<�j�<�@J<`H< T|<(�<8q�<�$"=��K=��r=�q�=+�=�!�=[p="�=@vx;��I�ym��o�����vI���I��ۅ��g��g�Ϳ@𿈖�&��(�H������`l�>��)�̿G-��W~����F��   �   P	�|o���lg�5�뽨�����<��q=ݧ=�ٿ=�^�=�=Fg�=�(�=�4�=�V=̱)=��=<S�<((�< ��<���<(��<<�=P>=�jc=�ւ=�ɏ=�I�=z{�=�]s=�+=�\,;ES��E�,tu��ž,�q�M�I��N^���ѿP��V�	������Ҩ!�d��&k�^�	�|�#�Ͽ� ��1͆���J��   �   !O�����Fb�;��t��h6�<��p=z��=���=�I�=�ٷ=�5�=}ˎ=�Xi=��4=��= ��<�j�<�@J<�H<pT|<��<�q�<8%"=��K=�r=r�=z�="�=
\p=��=`�x;�I�ml�p�o������H���I�\ۅ��f����Ϳ?������|����N�v���k�A��P�̿�,���}����F��   �   �b��5��
�R��ѽPN߼|I�<��m=�@�=�=���=#9�=X!�=�
R=D_=P<�< Y�;@3�`Py�􄝼0&����g��2����;t�<\v=XE8=��c=З={=�f=`W=@#�;��.���콻�^�ڴ��)����>��}�jȠ�/_ÿ~v��� �"���T�f	��l�*��� �i4�S�¿e쟿��{��b<��   �   ��4���Q�:�ڕ���盼���<<�e=�]�=Ę=��=�i=dX#=a�<`-��pü�H1�ںq��͎�����4啽>�����Z�h����� �:�r�<�=*7G=��^=��T=�=x�@<�W�dXʽ��D�L墾����Ib-���g��I���g��>ҿ�?�h�l�l�
�.��̯����jZҿ{X��쒿�Tf���+��   �   �{Ҿ!���q�����6�d��<��W=ȋ{=��p=��>=�3�<@��:D�߼�lm��4�����$)��"�n!������}�����ͽ���3�0̃��<�m�<��'=T�7=�?=,2�<P���~��l$��"��S�Ծ>f��wK����������"ӿ�r濴��ˁ��d~��I翍
Կ�r���{���4���.K�X���   �   J��]��>���E� ե:K=��?=xWD=0=�m�<�C_��"M�����̂	���4��[��{�<뇾N��֝���ڀ�We�+�@�Ƌ�4{ٽ��� ��97�<��=|=L��<@��@H`����a�5����B��в+��]�bӇ���������hƿF]ѿ[տl�ѿ�iǿ�����/��e����'^��C,�g���   �   A(����)���ȴ���1<��=z�=��<(�<T�������～u2�L�o�I������ƾ�վA�ھ��־}*ʾGص�՛�4�|�6V@�4�,ޢ�|���;�`ܝ<��<<z�<�@�;�� �׳��*�Rc����ɾ��
�D4���^�1���U������"����������ϥ�	����b��B;a���5������˾�   �   8M��� \�h"����<h�<HC�<��;l�Ѽ/G��� �Z�M�摎�xI��Y� �������q	��F��J�P���o��lɔ�ʏY��U�����n`� μ�lǢ<P��<��<a�bW�08�ɺH�~9���վZ ��/���P�Q	o��s��^6��I���Ƌ�|y����q�
�S�ټ1�x��ؾ�F���   �   V�=.���^˼P��;��<�s�<��!<�ৼ�7�����5mU����¶ξ.������5���H�.U�F�Y�KV��J�98�t ����5Ծ���	.^�&Z�4���m˼���;���<\v�<��!<xҧ�,2�����hU�4���ξ�����z�5��H�?U�B�Y�QV��J��8��p �Ǹ�\1ԾG���(^��   �   �򧽲V� ���΢<���<D��<@t�zW�7>��H�c<��zվ�"��/�A�P�o��u���8��~���ȋ��{���q���S��1��z�$�ؾ�I���<M�I	��\�`7���<\�<�I�<���;ȕѼ�@��m���{M�C���E��-�4���}���p����C��G����Ak���Ŕ���Y�%Q��   �   �p�@k;�X�<��<Dz�<�,�;8� �$���6 *��e����ɾ��
��4���^�����W���ä�]��ڍ��H����ѥ�����d��r>a�]�5� ����˾�*��,�)�������u1<��=��=̎�<��<���������ｲo2��o����?����ƾվ��ھ)�־)%ʾ^ӵ�$ћ���|�P@�F��֢��   �    P�9PC�<��==T��< �껖M`�F���@a�q����E��Ĵ+�:]��ԇ�j��m����jƿu_ѿW]տ��ѿlǿ����e1������k*^�"F,�tj���󮾲�]��C���E��j�:JJ=b�?=[D=0=�<_��M�@���0}	�%�4���[��{��懾��������ր��Oe�l�@�����qٽ7놽<���   �   �z�<z�'=��7=�@=�0�<���]���^$�$��Y�Ծ�g�yK����Q�������#ӿ�t濷��ۃ��s���K�aԿJt��}��6���0K����}Ҿ�"��Et�����D���<��W=`�{=d�p=8?=�E�<��:8�߼&\m�%+�����&#����g!����l��Iu����ͽn锽��3������:<�   �   �;G=�^=��T=��=��@<�Y�eZʽ^�D�v梾D���hc-�n�g�mJ���h���ҿA��h��l�L�
������n���[ҿ�Y��#풿�Vf���+���񾳉��b�:�����8D��<j�e=�^�=�Ř=T�=Z�i=|`#=�t�<@p�LUür91�,�q��Ď�����cܕ��熽�Z�l��`���\�:$��<\=�   �   ��=�Á=@�f=�W=��;�.�ޤ���^��������v�>��}�ɠ��_ÿ_w�i� ����.U�
�.m������ �n5�:�¿,퟿C�{��c<�Tc��6����R��ѽ�S߼�F�<��m=@A�=��=j��= ;�=�#�=�R=�f=�M�<���;���p$y�|n�����8�g�0㼻�]�;���<�|=�J8=�c=�   �   N�=�"�=�\p=��=��x;l�I��l�˫o������H�<�I��ۅ�@g��ۓͿ~?�2���������������"l�Փ�ӕ̿-��"~����F��O�����Nb����B��|4�<J�p=���=��=cJ�=�ڷ=�6�=�̎=:\i=��4=X�=��<(u�<�VJ</H<8i|<L�<hz�<)"=,�K=Ƞr=!s�=�   �   ��=к�=&�^=�0�<D���c���8�� ���w��/';��I���©�:/տ�� �hl�D*��:�"�E���I�ƚE�x�:���)�4�������^ӿ觿�F�7�>a���T���\-�cf���bt���'=���=Rӧ=&��=~�=Q �=��z=�C=lZ=�I�<�ZE< ��; �;�&8;���;h<v<��<�I=�jH=
u=�&�=�   �   �c�=V�=��Z=ȁ�< q�嘤��<4�a����[����7���}��Ԧ�z�ѿ�G��d���P'��P7�4B���E�.B��C7��'�h�J�����Ͽ�!��x�z���4��������)��~���24��'=��=S��=Ub�==��=�b]=Z� =D�<(]7< �9����)��P��v��`Ɋ;�<���<�l+=Ɓ]=���=�   �   R�m=:�q=�L=���<��7��Ք�u�&��a��>���b-��pp�{P���4ǿ��(�������-���7�vV;�@�7���-�����g���ƿ����m�{�*����2i�����~�~� �ܷ��#=_��=b�=���=u�=8!J=�M=�2Y<p_���������N<7��aG��A�dP%����@�h�`�0;��<Rj=��K=�   �   ��&=�@B="�3=�!�<�4˻��y�Ge�����
{Ծ�k�yY[�������&�ݿR����Tn��X(���+��(�J��nV�����zݿ�}��B���Y�`��2�о�u��+�	�hoT� �x;�0=��c=�t=�kZ=��=L��<�wƻ��qk�����qʽL����c���HԽ벽3���8f-��ď�p8�;���<�   �   h�v<��<җ=d�< �A��?�d��5a��]���1	�@�@����f8��Vſ�G�X�����^���^�Z��b[�p��`N�m�ſ:e��צ�Ͼ?��������6[��佐!�p�; )=��6=�(=|G�<��>;xo����Hz˽x�
��,�?�F�$|X�nz_��"[���K��a3�P���Uཧ���j � ���   �   앣����;Φ< ܦ<`��;�%�:S��H�4��Ė�����@"�XeY�̞��� ���@ƿ��߿
g��Z� �XR��F����ٕ�߳ǿ~9���M��Z��Q"�.4��p���1��ݯ��ּ�W.<
�<T��<�ր<J!�ޔ;�<b��TW�� E�~�y�����������d︾ɕ���h���잁�ݘO��S��ν�f��   �   uL��X�μ� �:J<���;U��D���Zk�r|j��뵾M���1�جc��ǋ�V�������˿K ׿�Lۿ�׿�AͿ�6���?��m(��̺e�Wr2�|�������Mj�����v��$c�h�;<���<��<0���"i��+߽��/�*mw�E`���;ƾ�[�,� �ԛ	����.t
�y��e��hJ˾�������f�9�҃��   �   �/��QԄ��]¼ �9�T�;Ů�HW�J����)�����u�Ⱦn�	���2�כ]��R��Q~���ۣ�`2��)����譿�"��������`��l5�y��p?˾HV���,�_������`ox�P8<�;H��q�"��Nf@��-���1��mz��>��'� z9�3"E��I��#F�dY;��*��������¾/���L�H��   �   0�C�����R_��@�P;`�v; bk��oS�^}޽�M>�x����*˾���G�'��WH��oe�l�|��ƅ�2���Pa����~�Gh��eK���*�r��M�ϾrD����C�c��K_��惼 �P; �v;pzk��yS��޽�R>������/˾�����'��[H�te��|��ȅ������c��L�~�1Kh��iK�(�*���q�Ͼ�G���   �   �X��+,�񰹽�����x��><��;T	��P	q�>��^`@��)���,���t�;�?�'� v9�E�T{I��F�rU;�8*���2��~¾������H� (���΄�`P¼ ��9PS�;`ᮻ|^�����)�����j�Ⱦ��	�� 3���]��T������ ޣ�5��Ҭ���뭿%����������`��o5�Ŝ��B˾�   �   b���kQj�x���v��-c���;<dǔ<8�<d����i��!߽Z�/�tew��[��46ƾ�U��� �d�	�=���p
�>��}��1E˾$���F����9�{�F��pμ@��:�%J<��;�]��>���n��j��l��j1�(�c��ɋ�����x�����˿#׿DOۿ��׿IDͿ�8���A��:*��ʽe��t2�T���   �   �6��r��P1��௽ּXX.<��<���<��<H!���;��X��VQ�\E�(�y�U���u���,���鸾|����c��[��⚁���O��M�νP�f�����,�;�զ<(ަ< ��;`*�cW���4��Ɩ���C"�hY�p����"���Bƿ ࿦i���� ��S��G�����"���ǿ:;��1O��b	Z��S"��   �   ��>���&9[�n�	!� �;�*=��6=V�(=�X�<��?;hR����o˽M�
��
,���F�OtX�zr_�[�J�K��Z3�\���K�=����� b���v<d�<h�=��< wB���?�q��8a�`��:3	�D�@����9��ſ�I�z���������_�����\�~��2P���ſ�f����p�?��   �   W����о�v��B�	��qT���x; 2=��c=\�t=rZ=��=���<0ƻ&��`k�����&gʽ|��)�����>Խ�Ჽ򷇽X-�D������;t�<ޝ&=�CB=��3=�!�<�E˻�y�g� ����|Ծ�l�4[[�����	�����ݿ�R����ho��Y(���+���(�H��PW�X���{ݿ�~���B��^�Y��   �    �*�����i��8����~� @޷��#=P��=� �=���=�w�=�'J=�U= YY<����ݴ�����.7�8TG�dA��C%�t���rh�@�1;�&�<Fp=f�K=��m=&�q=��L=���<p�7�xה���&��b������c-��qp�KQ���5ǿ/��Җ����T�-���7�RW;��7���-�X��jh���=ƿ�����m��   �   �4�C�����&)�	���/4�B'=o�="��=ec�=H��=G�=�f]=� =��<Xt7< 6�9����w)��6��F�� ��;�< ��<p+=|�]=���=�d�=wV�=ޑZ=���<�q�����=4�����\����7���}�?զ��ѿMH����� Q'�HQ7��B�$�E��B��C7�'�Dh������Ͽ�!��֠z��   �   �7��`���T��F\-��e�� Wt���'=�=�ӧ=M��=��=m �=.�z=D�C=�Z=,J�<8[E<p��; �; &8;���;�;v<���<�I=NjH=�u=Y&�=��=���=��^=�/�<ܿ�����`�8�� ��x��^';��I��é�[/տ�� �vl�.D*��:�(�E���I�E�n�:���)�&�������^ӿ�秿���   �   �4����:���)�u}��@4��'=��=j��=�c�=b��=V�=�f]=� =��<0t7< 1�9���w)� 7�pF�����;�<L��<:p+=Ȅ]=���=�d�=�V�=��Z=���<�q�f���\<4�$���D[����7�p�}��Ԧ�'�ѿ8G�� ��bP'�rP7��B�6�E��
B�C7�X'��g�����6�Ͽ7!����z��   �   ��*�7�h�������~� ���`�#=&��=`!�=��=�w�=(J=�U=�XY<`	��0޴�����.7�DTG�fA��C%�(��rh� �1;�'�<�p=0�K=��m=��q=��L=���<��7�FԔ���&�a��H��Ab-��op��O��54ǿ"�𿞕�X����-��7��U;�j�7��-� ��Bg���ƿ;����m��   �   ��F�оSt��"�	�*iT���x;�5=��c=Ȼt=�rZ=L�=T��<�ƻ8��`k�����<gʽ���5�����>Խ�Ჽ˷���W-����P��;��<^�&=�EB=��3=�)�<`˻�y��c������yԾ�j�X[�
�����׋ݿKQ����Tm��W(�n�+�̝(�<��zU����+yݿP|��A��a�Y��   �   %�P����3[���� �`B�; /=z�6=�(=�Z�< �?;R����o˽[�
��
,���F�^tX��r_�[�F�K��Z3�F��|K�⋖���]��v<$�<؝=�!�<��@� �?�����2a�\��r0	���@�h��7���ſF�J�������N]���,Z�T��`L翭�ſ�c��a��ؼ?��   �   �0供n��`1��د�	ּpu.<��<���<p�<@!�,�;�rX��TQ�bE�3�y�^���|���4��긾����c��T��֚��ڑO��M��~ν��f�T~���A�;ݦ<��<@ҁ;���N��`�4�~���?"��bY�S���%���>ƿi�߿�d��� ��P�JE�~���p�ῴ�ǿ�7��L��aZ��O"��   �   {����Hj�|���v�Xc� <<є< �<Е���i��!߽P�/�tew��[��:6ƾ�U��� �h�	�@���p
�>��v��%E˾���.��i�9�lz�-E���jμ �:�;J<���;F������Xh�Rxj��赾m��I1�֩c��ŋ�C���������˿�׿�Iۿ[�׿?Ϳ04���=��}&����e��o2�`���   �   >S��,���������w�X[<@0�;����q�Л�B`@��)���,���t�;�D�'�v9�E�Z{I��F�sU;�6*���!���}¾������H�>'���̈́� I¼ 8�9 ��;����N�a����)�芈���Ⱦ�	���2�a�]��P��|��'٣��/������H歿���p����d�`��i5���s;˾�   �   $�C���B>_�҃���Q;�cw;HQk�
mS��|޽rM>�o����*˾���K�'��WH��oe�r�|��ƅ�5���Qa����~�Gh��eK���*�h��6�ϾRD��>�C�M���G_�݃� cQ;�xw;x>k�~dS�v޽�H>�?����&˾[��#�'�TH��ke��|�,ą�Ő���^���~��Bh��aK���*������Ͼ�@���   �   ����Ǆ�L9¼ \�9��;�����S�7��n�)�����l�Ⱦn�	���2�ڛ]��R��S~���ۣ�c2��+����譿�"��������`��l5�n��R?˾ V��*,���������x��\<0M�;P�����p�ғ��Z@�&��\(��Qo�8���'�r9��E�wI��F�oQ;�~*�C��j��By¾����H��   �   (>��Wμ��:�HJ<���;�K��Ġ���j�7|j��뵾K���1�ڬc��ǋ�X�������˿O ׿�Lۿ�׿�AͿ�6���?��k(��źe�Nr2�r������KMj�t��n�v�c�@<<֔<� <�����i��߽��/�0^w�=W��1ƾ�O羲� ��	����Um
��}�h�뾿?˾o���W��F�9��p��   �   Lh��`�;��<<�<�ρ;�!�R����4�lĖ�����@"�XeY�̞��� ���@ƿ��߿g��Z� �XR��F����ו�ݳǿ|9���M��Z��Q"�4��p��l1�\ܯ�xּ�p.<�<p��<���<�� �6w;�gO���K��E�*�y�ϓ���������举*����^���z��������O��G�uν �f��   �   @�v<�(�<\�=�$�<��@� �?����F5a��]���1	�@�@����h8��Wſ�G�Z�����^���^�Z��b[�p��^N�j�ſ9e��Ӧ�ʾ?���r����6[���`!��5�;�/=l�6=8�(=Pj�< 8@;�6���ze˽i�
��,�{�F��lX��j_�4[���K��S3����@�������@0��   �   N�&=JB=�3=�+�<�˻��y��d�����{Ծ�k�zY[�������'�ݿR����Vn��X(���+��(�J��nV�����zݿ�}��B��	�Y�Z���о�u����	�mT���x;�5=��c=f�t=RxZ=��=���<��Ż���&Pk�B���]ʽډ�C��ے�i4Խز�9����H-���� ��;��<�   �   ��m=Z�q=z�L=��<��7�Ք�H�&��a��:���b-��pp�zP���4ǿ��*�������-���7�vV;�B�7���-�����g���ƿ����m�y�*����!i��J���~�  ˷ �#=���=u"�=���=Az�=.J=l]=�|Y<0����ƴ�<���!7��FG��A��6%�u��Fh�`*2;�7�<hw=Z�K=�   �   �e�=�W�=��Z=܄�<Hq������<4�Z����[����7���}��Ԧ�{�ѿ�G��d���P'��P7�4B���E�.B��C7��'�h�J�����Ͽ�!��y�z���4��������)��~��`!4�0'=��=���=Md�=v��=��=Rj]=F� =�$�<p�7< 7�9�b��])���`���$�;�4<���<2t+=�]=*��=�   �   ���=��}=�<=�+s<$E��cｔ�n���ʾ���lc������ʿK����j��4�[M�j�b���q���v���q���b�t�L��93��_�{���K�ȿ|���y�_�	��žԅe��޽�����<\�_=�r�=�K�=�͐=2�x=L�@=��=ෆ< �.;��	�ā�LP���x���?�`�P-<`�<R4!=��V=
�~=�   �   �=��r=Ry7= �r<��m齐Ri�"�ƾ����D_������ǿ��������0���I�d~^���l���q�$�l��k^��0I��40�l��c�����ſ���T�[��&�-���vb`�)ؽ����k�<��Y=��=F%�=�م=��\=0x=�۲<�@�;�#�����I���d	���(�ϼ(`p���P�8�t<�/�<0%;=�h=�   �   0GN=�YR=
p&=0&m<���"�ֽT�Y��f��F4��2S���������j��X��'�d�>�~�Q�H_�J�c�HH_��-R�H�>��'�V�������1����yP���� ��r�Q��@ǽ`Ǽ�(�<�<G=�	t=�vp=�H=$N=HW<�C�\G����H��у�����c"��)V���ϊ�b�\����}}��4�;�:�<Σ&=�   �   V�<fu=��=2Y<ؼ�.����A���������X@�����r��?Yڿ*������g.�[?� �J�dO�r3K���?���.�>@�J����ٿ�/�����:f>�R��e��2�:�*���,z��h��<�%=9=NE=ɩ<��J��d ���{� �����F[�����c"�\��r"�S�����ǽ;���z ���5��dO<�   �   ��L��k�<$\�<0O'<������b�#�r�����]l(���i�E*���¿���n������))���2�\l6��V3���)�.��>�	�T���V¿�����i�dO'�~⾬t��Z5����P�o��W�<��<H\�<���;�����g�[�ǽ$E���;�y�b�W��=a��fQ�������:����h��B����׽�!��p<��   �   ��-��)A�0�; ��;X�{��l�Ĉ�^�k��ν��x��.F��������})ʿ�.�P=��d�jl�zk�����L��A����|˿�b��5탿�@F�� �����lh�X���
�[���0� m<�'<@��������l3�b�A������ڟ�㻾�LҾ���1��vZ�h�ԾJW��<ޣ��턾�,J�x\��Ү��   �   Mƽ4J�<���`û���N�8�)���½<�5�i��.�5� �3�W�ޞ����g�Ŀ9v޿Ϳ�� �t}�j� �9����࿅�ƿ����Ċ�s7Y���!����𕾪�4��뾽@��H � !� 'c��3�����Z��v�g�L���0^˾h���'�3����(��,��)��^ �@�f���l)о�)��>,p��.#��   �   ��(��ƽ�*F��\����X�X�WJ��p��M�_��O��+����R)��Z����,���B��]�ÿ5�ο��ҿ.�Ͽ��ſ���%�k���,�\�D1+��%���ாx^a���x�����ؼ��9�����(�7�����]#�\s{�����q�O��_D2�<�L�g�a��Jo��`t�xcp�l�c�*AO��5�f��W��D��+���   �    }����������$��ّ�����؛��,��j]��ox��S��R�����$���L�w6s������"��z砿�*������d���;��V�v� �O�m�'��� �Rn����|����냮���$��ב�L������2���a��ux��W�������$���L�;s�����q%��L꠿�-��͜��ng��->����v���O���'� � �r���   �   �㮾�ba����������ؼ��9�x���N�7�O��ZX#�Rl{�B��5l���u@2�ަL���a�Fo��[t��^p�Şc��<O�5��b��R�@���'����(�i�Ž�"F�hU��0�X�\⼁N�����R�_�]S��ݥ���U)��Z�������E��PĿH�ο��ҿ;�Ͽn�ſ�"����v�����\��3+��)���   �   ���U򕾚�4�eﾽ
�� ����躠c���3��������g������X˾��$�P����(���,��)�&[ ��<�.��� $оF%��`%p��)#�nEƽ�J�̧��p���H�N��)���½��5�!���1㾶 !�b�W�Π�������Ŀy޿��� ��� �;���J����ƿ1���PƊ�H:Y���!��   �   *"�����ooh�����6�[�ؔ0� y<H�'<�ų����؂���-�J�A�k����՟�~ݻ�wFҾL�����&T�q�Ծ�Q��k٣��鄾
&J�W��ʮ���-��	A��?�;���;��{�Z�l�2��-�k��ѽ��z�1F����r����+ʿI1��>�f�n�&m�l��TN�PC�W��~˿|d���CF��   �   �P'���v���6������o��[�<���<�j�<@$�;�|���g�ջǽ�>�P�;�G�b�����\���L��~���6����h��B�����׽��� $뼀�J��w�<tb�<Q'<D��ɮ����#�F��F��.n(�4�i��+���!¿��꿤��
��V+)�|�2� n6�JX3��)�r��V�	�'��X¿�����i��   �   _g>�$��z����:�~���8{����<<�%=6!9=�L=ܩ<�%J�V ���{����o�(U����^]"����k�D�����ǽХ������5� �O<Lb�<Zy=��=�1Y<�ؼk1��ЉA�%�����hZ@���������Zڿ��� ��h.�d\?�v�J��O��4K�
�?���.�&A�
����ٿ�0��ϻ���   �   kzP�z�����J�Q��Aǽ�`Ǽ�*�<�>G=0t=L{p=(�H=�U=�@W<@��-����H�1ʃ�����T��@N��Ȋ��x\�����S}��z�;�H�<$�&=KN=\R= q&=@$m<���7�ֽ �Y��g��*5��3S���������k�Y���'�T�>���Q�l_�p�c�\I_��.R��>���'�����	쿍�������   �   ��[�"'�l����b`�C)ؽ��`m�<�Y=���=|&�=#ۅ=��\=�|=��<0r�;�l#�X����:��D]	�f�� �ϼPFp���O���t<�7�<l(;=��h=V=|�r=�y7=��r<����齨Si��ƾ=���E_������ǿ�������0�H�I�^�d�l�t�q���l�xl^��0I� 50��������8�ſ����   �   D�_���Êžr�e�޽����<޻_=�r�=�K�=�͐=t�x=��@=�=@��<��.;`�	��Á�@P��y���?�@�@O-<�_�<4!=\�V=��~=���=��}=��<=�(s<F�*d���n���ʾ��mc�8����ʿo����j��4�[M�x�b���q���v���q���b�d�L��93�z_�Y���+�ȿ\����   �   ��[�d&�a���Ra`�e'ؽ@�⼀p�<�Y=>�=�&�=:ۅ=��\=�|=��<�q�;�l#������:��V]	�v���ϼFp� �O���t<88�<�(;=��h=�=J�r=�z7=`�r<����4Ri�܃ƾw��}D_�����@�ǿ����j��8�0�R�I��}^�*�l�2�q���l�bk^�0I�>40�������g�ſ���   �   xP��������Q�3>ǽ\WǼ|0�<�@G=Vt=�{p=��H=V=AW<��$.��֠H�Iʃ�ح��c��LN��#Ȋ��x\�����R}� }�;�I�<Ʃ&=LN=p]R=,s&=81m<ֿ���ֽ:�Y��e���3��1S�I������i�jX�b�'���>���Q�4_�&�c�*G_��,R�^�>�R�'���������t����   �   �d>�0�����Ұ:�����Hn��X��<�&=�"9=^M=ݩ<�"J��U ���{������7U����i]"���o�A�����ǽ��������5���O<e�<f{=��=�CY<@	ؼD,����A�R������W@�����n���Wڿb������f.��Y?���J��O� 2K�p�?���.�8?�l��!�ٿ�.������   �   �M'����r���2�Ǌ��`to��e�<��<Dn�<�,�;�{���g�ջǽ�>�`�;�\�b�����\���L��
~���6����h���B�����׽~���!� `J�D|�<�i�<�f'< �������.�#����}~��j(���i�)��2¿���T��b��^()�L�2��j6�U3��)�ҋ��	�G��?U¿V����i��   �   ������ehh�I���p�[� s0���<��'<p�����������-�L�A�p����՟��ݻ��FҾV��ɀ�/T�t�Ծ�Q��d٣��鄾�%J��V��ɮ� �-���@�_�;Ɋ;P�{�~l�B����k�j̽��v�e,F����ϔ��r'ʿV,��;�c��j��i�*��DK��@�k��Uz˿�`���냿t>F��   �   ���F핾��4��徽���� ����b� �3�u�������g������X˾��$�V����(���,��)�([ ��<�(���$о7%��0%p�:)#��DƽBJ�䟗����P�N���)���½��5�����*��� �Y�W�����刺��Ŀ�s޿Ҽ�b ��{�͂ �$|�������ƿ҈����K4Y�N�!��   �   Oݮ�#Ya����K�����ؼ�9�𕑼�7�_ ��X#�8l{�?��8l���{@2��L���a�Fo��[t��^p�Ǟc��<O�5��b��R�@���'��t�(�0�Ž�F��I���uX���E�������_��L������O)��Z�������/@����ÿ3�ο��ҿ�Ͽ��ſ���<���z�\�B.+� !���   �   3�|����|��Ԓ$�@Ñ��}����U+��]�Xox��S��R�����$���L�~6s�����"��~砿�*������d���;��U�v���O�g�'��� �6n��J�|�l��>���j�$�@ȑ��z�����W&��&Y��ix��O��b�����$��L�+2s����� ���䠿�'��1���b��29���v��O�'�� �j���   �   N�(���Ž|F��?��(pX�\	�OH�������_��O��$����R)��Z����0���B��a�ÿ8�ο��ҿ1�Ͽ��ſ���#�i���&�\�<1+��%���ா^a�0��:����ؼ��9�������7�����fS#��e{�	���f쾸���<2���L��a�0Ao��Vt��Yp��c��8O�&5�\_��L�<��0$���   �   .<ƽzJ�ؐ���`����N�ė)�;�½��5�K���-�3� �5�W�ߞ����i�Ŀ=v޿Ͽ�� �v}�j� �:����࿂�ƿ����Ċ�m7Y���!������4�$꾽x�������纰�b�p�3��x��K��8�g�i���tS˾���� ������(���,���)�@W ��8������о� ���p��##��   �   ��-���@� ��;pފ;��{���l����k��ν��x��.F���������)ʿ�.�R=��d�jl�|k�����L��A����|˿�b��2탿�@F�� �c���lh����v�[� y0�h�<(�'<�s�����_z��R(���A�[����П�ػ��@Ҿ��\z��M�a�Ծ8L��hԣ�Z儾�J�9Q�#����   �    �G���<r�<�m'<`���c����#�R�����]l(���i�E*���¿���p������))���2�\l6��V3���)�.��>�	�R���V¿�����i�^O'�g⾃t���4�\��� |o�Tg�<���<hz�<�t�;0c���g�ܱǽ�8�Q�;�a�b�����W���G��_y��2��N�h���B�< �7�׽���h��   �   8s�<V�=��=`HY<�
ؼ�-��a�A�s������X@�����u��BYڿ*������g.�[?��J�dO�p3K���?���.�>@�J����ٿ�/�����4f>�L��J��Բ:������r�����<�&=�&9=�S=h�<�nI�H ���{�a�����6O�P���V"����L������ǽ䜌�X����5�`�O<�   �   �PN=�`R=0u&=p4m<<��h�ֽ"�Y��f��E4��2S���������j��X��'�d�>�~�Q�J_�H�c�HH_��-R�F�>��'�V�������0����yP������5�Q�(@ǽ8[Ǽ�/�<�AG=�t=�p=��H=]=�cW<p�
�����H�������]��YF������pj\� ���&}�pȳ;<Y�<�&=�   �   D=�r=�{7=��r<����{Ri��ƾ����D_������ǿ��������0���I�f~^���l���q�$�l��k^��0I��40�j��a����ſ���U�[��&�%���Zb`��(ؽ0��|o�<`�Y=��=�'�=}܅=��\=�=��<�;�R#�T봼�+���U	�چ�X�ϼ�*p� �M�0�t<�A�<�,;=��h=�   �   �Ot=�K`=r�=@g�:$n���H����=x8��p��r����鿢�fW1�0�Q��r�����������@����ن�"nq���P��0�����Y翁���B���{�5�+r쾢7��q� V� ��;
-=�iv=X*�=�qw=.�I=�X=X�<  �6��y����fL�S�6�8x� ;���ρ��sK<�6�<�s4=l�a=�   �   )b=�/T=Ȏ=�ŗ:�g�xq��ꍾ�:�:5�a��X����`���9.���M��m�>��f������mk���	��̵l��3M�--�B��C����Tq��rS2�^��*<��L�>P� ?�;�&=�!j= x=��^=FN*=p��< ��;@�R����B0��:T��fb��FY� �9� ���j����:, <��=�I=�   �   ��*=��.=ذ�< �1:V���
�~U޾��*�ov�r���ڿ*���S%���B�M_���w�Ev��]���t����9x��^_��}B�
�$�n����ؿ�����s��(��wھ�����4�.@����;d=4aD=�>@=��=��<�،�P_�f?W������κ���ѽ}�ڽ��Խ����㞽��h���X���\Q<�j�<�   �   tT�<��<��< d���<������Qn���ȾRO���`�]����ȿ2K������2�t�J�-`�&�n�)t�.>o�f�`��K�vU2�:������� ȿ���z_�����ž��h�Y���#)�@4�;Xb�<x=�ؾ< h�;�޺��j`�::�����ER�H�4�� E�@K��F���7�wl �Z����(�v���� s���   �   (���`�O;�D<`%��ԭ!���нUL�)��������E��-���j��+�߿J������2��wD��nP�"�T�Q��qE�
�3�b���{�C�߿�:��2�����D��b�����z�G� �Ƚ��� Ԝ�0Q<�p<Г>�TK0��1��_q�4 8��i��9��v��ɼ��:�����Z➾����J�o��/>���q.uF��   �   �ރ�l��w5���<�X�8ݨ��_&����̣���&�1�g�jԘ������������l���'� R1���4���1�`�(�������P�n]���3��-�g���&�����N��
y#�Ӧ���w��8�����<μ��s�^�ܽ��+�>�p�8��t����ྒྷ���q�����A��������yDľ����w���1�z'��   �   ���x������#��ā��k(��� ��a��������S=�{�{�����u¿�������V���P��1�$��ơ�N%�����ÿV꠿TW}��>��/�]崾��`��F��L^~��T뼠c���0�ᑌ����ooE��n��4���-��`����(���:�,lF�d�J��AG�IW<�I�*�"��=���lþ֑��0K��   �   G%R�f��R���)$��'���F�zt��x�'��&��<�Ͼ���Q�F�v�~�N���綿<�οW��f1�a���%�g����п�߸��k��r�����H���saѾ�ۉ��(��`�C��=��Hd�n捽�+����M������վ�|�hi/��:Q��Jo�䊃��D�� ��oԋ������q���S�H�1�&����پ;m���   �   ���[�E����PҀ�ؽ�f����}����B�������۾���A�/yo�����堿_#�����Y���oǺ��v�����{C���r�EyD�x��:x޾މ���E�8��cπ���������}�ӥ��B�����{�۾3��� B��}o������蠿o&��"�������ʺ��y��勢��E��*�r��|D�N���|޾�   �   �dѾ7މ�(�V򺽴�C��9���]�����g#����M�������վKy��e/�j6Q��Eo�6���)B��8���ы�p�����q�6�S���1����پ�i���R��������%$��'�$�F�3y��X�'��)��DоL����F���~�ž���鶿W�ο����4����r)￯����п]⸿.n��c����H�d��   �   �1��紾
�`��J���a~��R�HZ���'���������hE�nj���}����򾳋�d�(�/�:��gF���J�"=G��R<�@�*�����6���gþ!ґ��*K�(������|��@�����#+���� �P�a�����7��tV=��{�ͺ��¿��⿑ ����R�l3� ������&�R�<�ÿV젿�Z}�(>��   �   ��&��ᾃP��{#�����x�����[���ͼ��s�@�ܽ%�+��p�R��������ྡ��˜����h=���������>ľ\���P�w�l�1���׃���b5��<�Z�F਽rb&�4��������&��g�5֘�����=��\���n�t�'�T1���4���1�*�(����
��S�[_��C5����g��   �   W�D��c�B���[�G���Ƚ��� ���@"Q<��<xf>�<<0�(��]k��8���i�<5��X��l������Ȱ��Nݞ�𩍾zo��(>�M�M嶽8gF�𫈼�6P;�S<P ��d�!���н
L�@�������E�/��;l��2�߿~����6�2�pyD��pP�0�T�Q�rsE���3�����|���߿<��I����   �   �_���E�ž3�h��콦$)� @�;Pi�<�}=��<���;pú��Y`�@0�������K�B�4�wE��8K���F���7�f �|T�p���8�v�p�@:��lb�<@��<���< d�J�<����=Tn���Ⱦ�P���`���� �ȿ�L������	2���J��.`��n�+t��?o��`�<�K��V2���)���ȿ����   �   λs���(��xھ ���25��@����;�=�dD=D@=�= �<����$F��0W�����	ƺ�f�ѽG�ڽr�Խ`����۞���h���o�X|Q<�v�<�*=��.=4��<�s1:zV�����V޾��*�zpv�R���ڿԕ�lT%���B�HN_�(�w�w�����'���;x��__�V~B���$������ؿD����   �   �q���S2����Q<��h��=P��E�;l�&=�#j=�x=*�^=�R*=���<�Խ;@R����0�42T�^b�>Y��9�����]���:�ˠ<��=�I=+b=�0T=�=���:��g�Dr�[덾�;��5�������%��Ĩ�::.���M��m����f�������k��
��N�l�D4M�j--�x�����J���   �   #���I�5��q�j7���p�V�p��;�-= jv=�*�=$rw=v�I=�X=��< ��68�y�t��NL�S�6��x�;���с��rK<H6�<Js4=�a=rOt=rK`=��=�P�:$n������(�qx8�q�������鿶�|W1�H�Q��r�����������;����ن�nq�z�P�t0�����Y�_����   �   �p���R2�u�羄;��W�;P�`S�;��&=l$j=x=b�^=�R*=��<�ӽ;hR�4���0�V2T�&^b�">Y�,�9�����]�� ƛ:�ˠ<��=�I=�+b=�1T=F�=@�:Ļg�*q��ꍾM:��5�4����)��&��r9.���M�Rm�����e��*���k��Z	�� �l�R3M��,-�����㿌���   �   ��s��(�ovھx���,3�T@����;�=BfD=�D@=D�=��<@���LF�1W�����&ƺ���ѽ`�ڽ��Խt����۞���h�����n��}Q<x�<�*=*�.=���< V2:�V��i󄾖T޾N�*�4nv����:�ڿ����R%��B�L_���w��u�����������8x��]_��|B�F�$������ؿل���   �   �_�����ž��h�L��h)�0e�;(o�<x=��<;�º��Y`�L0�������K�W�4��E��8K�ͯF���7�$f �xT�\����v� o�� ��e�<d��<��< �b���<������On���ȾWN�v�`�x����ȿ�I�����2��J�j+`�X�n�8't�T<o���`�j�K�<T2�6�������ǿ����   �   ��D�a�����N�G�M�Ƚ��� �0Q<��<�a>��;0�(��^k�8���i�K5��g��y������Ұ��Wݞ�����!zo��(>�8�嶽DfF�Ȩ��@]P;�b<0�\�!���н�L�j���G���E��,��"i��k�߿8�8���2��uD��lP��T�	Q��oE�f�3�����z�K�߿
9��㽇��   �   ��&�R��yL���u#�p��� e�����`=�x�ͼ^�s���ܽ�+��p�W��������ྰ��Ӝ����m=���������>ľV���<�w�@�1����փ�з��Q5�`�<����ب��\&��������&���g��Ҙ����\�迄��bk�Һ'�2P1���4���1���(�b��6��/N�K[���1��[�g��   �   �-�%ⴾ��`��?���R~��?��M��&$��]����hE�jj���}����򾹋�n�(�9�:��gF���J�)=G��R<�C�*�����6���gþґ�~*K����1���L��`��4p���#���� ��a�����$��Q=�<�{�����¿���������$O��/�F������#����I�ÿ(蠿�S}��>��   �   W]Ѿ�؉�R�'��纽�|C�h'��X�ߍ�a"��|�M�腙���վNy��e/�r6Q��Eo�;���-B��;���ы�s�����q�5�S���1����پhi���R������f$����F��n����'�$����Ͼ.��0�F���~����x䶿B�ο���-����}"�}㿹�п�ܸ�bi��Y���}�H�I��   �   .���zzE�����Ȁ�����~�}���潠�B�㝗���۾ ���A�5yo�����堿d#�����\���sǺ��v�����zC���r�AyD�p��"x޾����rE�o�齚̀�������Z�}�֗�2�B�����Q�۾J����A��to������⠿g �����$���Bĺ��s��A����@��]{r�wuD�^��as޾�   �   �R����W��`$�f�x�F�9r��Ό'��&��)�Ͼ���S�F�{�~�Q���!綿?�ο\��j1�e���%�g����п�߸��k��p�����H���QaѾ�ۉ�(�e캽ҀC��&���S�eڍ�����M�6�����վAv��a/�'2Q��@o�����j?��g���΋�������q���S���1�Ͳ�hzپce���   �   ���s������x��0o��a%��� ���a�v������S=��{�����x¿�������X���P��1�&��ơ�N%�����ÿW꠿PW}��>��/�0崾�`��D��X~�|A뼨G����샌������bE�xf���x�����/��l�(���:��bF���J�~8G�pN<� �*�ݳ��0��qbþ�͑��#K��   �   qσ����75� �<����ڨ��^&�֠�������&�3�g�lԘ������������l���'� R1���4���1�`�(�������P�m]���3��*�g���&�k�ᾖN��Ax#�W����h��H��@��ͼ��s���ܽ��+�e�p�����J���t���x��5��J���9�����:��-9ľi����w���1�u��   �   ,�����P;Pv<�����!���н�L����{����E��-���j��/�߿L������2��wD��nP�"�T�Q��qE�
�3�b���{�B�߿�:��0�����D��b������G�C�Ƚ.�� ����>Q< �<�8>��-0�����e�"8���i��0��`��&���e��s���3؞�9����qo�J!>�-y�D۶�$WF��   �   $u�<���<蓲<��b���<�W���xQn���ȾPO���`�_����ȿ6K������2�v�J�
-`�(�n�)t�.>o�f�`��K�vU2�<������� ȿ���x_����žG�h�	���)��e�;�s�< �=���<��;t���J`��&��s����E�r�4�AE�.1K�o�F���7��_ ��N�O����v��S缀Ȝ��   �   N�*=��.=���<��2:tV�����qU޾��*�ov�s���ڿ,���S%���B�M_���w�Fv��]���t����9x��^_��}B�
�$�n����ؿ�����s��(��wھd���L4��@����;= iD=&I@=b�=X$�<04���.�@#W�Ж��������ѽ1�ڽn�Խ���Ӟ��h�F���C�ؠQ<��<�   �   F.b=�3T=��= �:��g�Jq��ꍾ�:�:5�b��Y�����`���9.���M��m�>��f������mk���	��̵l��3M� --�@��C����Sq��rS2�X��<����<P��N�;ҕ&=�%j=x=6�^=bV*=L��<�;HeR�hv��0��)T�XUb�h5Y���9�β��O��@��:@֠<&�=~I=�   �   p�Z=:�D=(��<��/�����5�@��������O��5���ȿ���"�X�F���m��|��!����)��!F���#��~i���+��:�l�ΡE�x!��� ��ƿm����LM����_�����0�����0���=��R=�h=3T=�o"=,*�<P��;@9c�4���^E2� mU�ƹb���X�ܿ8�&k�tS���2�:�0�<�=�F=�   �   �G=N�7=��<`�1�e���p�1�䂣�4.�L�K�[����8ſ�������7C�0i�.}��=���U��~\���[������F���Bh�,*B� ��tq��$oÿ�)����I��^�t���2�,��p�������<h}E=��T=dL9=d =�Q<����<��v]=���x�ܱ�������z���f�֧F�\����0��&<��< �+=�   �   

=��=@�<`�:�����N&���������T�@�_���i���
�����8�.�[��"~� ���~���>��/���zG��H5~��U[��D8�$9���H���∿��>�����h���v�!��V��8�@��<�[=��=8��< =�;˛�<�:�X(��ZHý��(N�[��P�jc�tȽ�N��RsH�ݷ� <;h��<�   �   � <�[�<�AA<x�W��=�����P��V径�/�%�|�{����߿���TL)���G�~e��<�u���!ˋ�QĈ�4��Jf��H�TA)�\q���޿�'����z��.�@���'���@���t�0�#��5u<h�<hp7<��!�*�!�5����#������:�b�U��g�U,n���h�}DX�h�=�h���������0�8�[��   �   !��0��`�J�����(�d�  �קn��Ǿ����^�q��K�ƿ�����T��C0���H��]��l��sq�̹l�4�^���I�N1�n��c���ƿe��t�]����1Už_k�����$Y��sl� $�P���@8޼�}��PڽF"��@Z�f����Y�� ������G�ƾϭ¾}���&J���ي���^���&���⽢1���   �   Ƃ����7�|�ȼ0�ͼ�LL��ԽE�=���#�!�<�� ��bҪ��yֿX��
I��<+���;���F�� K���G�p�<��d,�ZF��<�HG׿�)��,*��8;<�4� �������B�-�Ͻz�B�����:��2G+��u�����zL�ZČ�!`���ݾ
V �>������;�Tx�b����߾�2��?g��.Q� ���   �   ���X���V\�<c�>�?�"���h]�����~}Ͼ�&��zU��F���v���@ؿ?}��t�d��.2$�Nn'���$�X}�j��M���5�ٿ����%V�mb��kϾY���3�6ѧ��9������R�~�������i��*��
�۾�z
�I&�K?���R�2z_��d�U5`�OT���@��(��?���޾�ק�hnm��   �   �au�&��\����h���D�7���s��`�F�Lٞ�����'��9`��Ҏ� ��c�˿�^�dG��(w������$���@�C�Ϳ����o����a�(�(�/�h��V3G��:�Ȇ�x�@��Vc��b�������q��l���������LF��k��b��Qr��x囿����f���Z���kn��H�Hw!�����ո���   �   B�����g�2S�_o���s^�~�]����v���e�_!��������)���Z�e���ᒞ�Eǳ�=|Ŀ�NϿ�Gӿ��Ͽ
�ſ�E������܇�-�\�ؒ+��8������ڞg�P�l��Lr^���]��#��.��e�Q%�����&�)���Z�߈������fʳ��Ŀ�RϿAKӿiп[�ſ�H�����Y߇� ]���+�a=���   �   ��|k���6G��>�nɆ�r�@�Pc��\��&��U�q��h��2������nHF��k��_��]o��e⛿�����c���W��@����n� ~H��s!�=��������[u�|�F����h�r�D�� ����齧�F�~ܞ�!���'��=`�+Վ�5#��{̿Pb�K��y�����������YC�7�Ϳ���������a�կ(��   �   d��nϾ�Z���5�ӧ��9�����R�����Z��Mi�)&��/�۾w
��D&��?���R�u_�nd�70`�rT�4�@��(�y<���޾bӧ��gm���ZR���N\��_�j�?����P`������Ͼ$)�~U��H��y���Cؿ~����u�f��P4$�zp'���$�P�,��a�����ٿE��������'V��   �   ==<��� �������B�C�Ͻ��B� ����+���;+�Pm������rL�ӿ���Z��Vݾ{R �a{�ۯ����7��t���l�߾�-���b��4'Q���:{��h}7���ȼ�}ͼ�NL��ԽE��¥�����<�5"��[Ԫ�#|ֿ��J��>+���;�&�F�>#K� �G���<��f,��G��=�gI׿�+���+���   �   G�]�����Vž ak�����%Y�jl� ��L��d޼&}��Eڽ�"��8Z������T��o������8�ƾާ¾�}��E��Պ��^�*�&�|���)���
��H�� hJ�0�����d�� �Ԫn�!Ǿ�����^��r��!�ƿ����0V�ZE0���H�*�]�ll��uq�,�l�T�^���I��1����M��l�ƿ����   �   �z��.�����(��zA�`�t�{#�Eu<���<��7<�w!�"�!��񘽼潒��r�:���U���g�$n���h��<X�\�=�*}�u��Ȳ����0�8�[��> <�e�<�KA<��W�R?��(	� R��_���/��|����M�߿|���M)�P�G��e��>�����K̋�lň�*���f�H�VB)�&r��޿�(���   �   Q㈿��>����������!�;W����H��<�_=>�=`��<���;س��f�:�] ��v?ýN��I�>��K��Y��kȽ�F��fH�Ƿ� �;�ı<�
=��=�B�<H�:����P&�Η��)���t�@����j���N��t�8�\�[��#~�� ������?��
���:H���6~��V[��E8��9�g������   �   -*����I��^�����R�,��p�� ����<�E=��T=6P9=, =�0Q<����̞��T=�^�x��������.v��^���F������0�x;<H��<B�+=G=��7=���<H�1�^���P�1������.���K�О���9ſÈ��(��8C��i��}�����`V���\��-\��c���dF��Ch��*B�<���q��goÿ�   �   L���eLM����!���n�0�+���0�滢�=.�R=d�h=f3T=,p"=�*�<@��;�8c�����8E2�mU���b���X� �8�Pk��S�� )�:$0�<(=��F=�Z=��D=���<��/�e��~�5��������ƹO�6��,�ȿ4��6�"�r�F���m��|��,����)��!F���#��ui��y+���l���E��w!�~� ���ƿ�   �   �)���I�^�����#�,�No�����P�<d�E=F�T=nP9=> =�0Q< �����
U=�v�x�������=v��^���F������0��;<���<��+=�G=N�7=D��<��1�˦���1�����.�	�K�)����8ſ����v��&7C��i��|�����jU��\��8[�������E���Ah��)B�����p���nÿ�   �   ∿��>����A�����!�YT�� �ܬ�<ba=�=0��< ��;������:�q ���?ýt��.I�Q��K�	Z�lȽ�F��fH��Ʒ���;Ʊ<�
=n�=xG�<�:�����M&����������@����i��
� ����8�0�[�F!~�N���}���=��L����F���3~��T[��C8�n8�l~�] ���   �   ��z�&.�)��x&��a>�^�t��f#��Qu<���<�7<Pu!��!����潤����:���U�Ϟg�"$n���h��<X�h�=�2}�r�����"�0�(}[�@D <�i�<�YA<X�W�7;�����O����m�/���|���w�߿���LK)���G�`|e��:�Y����ɋ�/È� ���f�ZH�*@)�lp�A�޿k&���   �   7�]�����Rž�[k�C���Y��Ql� �� :���޼�}��Eڽ�"��8Z�ʟ���T��������J�ƾ�¾�}��E�� Պ��^��&�>��y)�����Xx� (J��t���d�� ��n��Ǿ���ك^��o����ƿ�����S�:B0���H�η]��l�
qq�b�l���^���I��1���5���ƿ����   �   �8<�l� � �����B�G�ϽD�B������#��$9+��l��Ԓ��rL�ؿ���Z��eݾ�R �l{������7��t���p�߾�-���b��'Q����hz���z7��ȼ�oͼXDL��Խ��D�������<�D���Ъ��wֿ���G��:+�p�;���F�~K�d�G�H�<�c,��D�6;��D׿�'���(���   �   `�hϾlV���/� ˧�p9��}���R�������(i�%&��3�۾w
�E&��?���R�u_�yd�@0`�{T�9�@��(�w<���޾Sӧ�xgm�>�Q��BJ\�Y���?�槪� Z�j���jzϾ�$�xU� E��{t��P>ؿ3z��Xr�r��0$�$l'���$�V{�������d�ٿ�����썿�!V��   �   ���_e��].G�H3�����l�@��Ic��Z������q�ph��0������tHF��k��_��co��k⛿�����c���W��C����n��}H��s!�0�������T[u�k{�3���h�<�D��������F�X֞����;�'�Q6`��Ў����x�˿�[��C��@u������n����<�*�Ϳ˥�� ���H�a�*�(��   �   ����Řg��K��d���e^�l�]�������e�B!��������)���Z�i���撞�Kǳ�D|ĿOϿ�Gӿ��Ͽ�ſ�E������܇�+�\�Ғ+�x8������P�g�1O�)i��i^���]�X��{�$�e����������)���Z����1���Dĳ��xĿ�KϿ.Dӿo�Ͽ��ſyB�����ڇ���\�j�+�-3���   �   �Tu��v�)��h�h�R�D�G�����齪�F�ٞ�����'��9`��Ҏ�� ��h�˿�^�iG��*w������&���	@�D�Ϳ����m����a�!�(��h���2G�U8�Ć� �@��Dc��U��z���q�Sd��̆��$��`DF�`�k�=]��l��_ߛ������`���T�������n��yH�@p!�a��� ����   �   ���I���@\�T��?�ک��f\�Z���\}Ͼ�&��zU��F���v���@ؿB}��t�f��.2$�Pn'���$�Z}�j��O���7�ٿ����%V�bb�qkϾ�X���2��ͧ�r9��z���R�%���.��x�h��!����۾�s
�A&�X?��R��o_�Cd�+`��T���@��(��8��޾�Χ�=`m��   �   r��o7�d�ȼ�hͼ�DL��ԽFE������<�� ��eҪ��yֿZ��
I��<+���;���F�� K���G�p�<��d,�ZF��<�HG׿�)��+*��1;<�%� �}�����B���Ͻ@�B���������.+�e������kL�����U��B	ݾ
O ��w������3��p�T���߾(��X^���Q����   �   ����xU���I� p����d� �F�n��Ǿ����^�q��N�ƿ�����T��C0���H��]� l��sq�ιl�4�^���I�P1�n��c���ƿe��p�]����Užm^k�����Y�PNl� ������t޼,�|��;ڽH"�L1Z�H���tO��������;�ƾ��¾4x���?��pЊ���^�l�&�p��!���   �   �g <dv�<�hA<��W��;�����P��?征�/�&�|�|����߿���TL)���G�
~e��<�u���"ˋ�RĈ�4��Lf��H�TA)�\q���޿�'����z��.�$���'���?��t�`f#�0\u<��<@�7<�J!��!�1阽2�r����:��U���g��n���h�5X�/�=��v�Q��b���
�0��M[��   �   �
=|�=�L�<��:�;��XN&���������S�@�_���i���
�����8�.�[��"~� ���~���>��/���zG��H5~��U[��D8�$9���I���∿��>�����H����!��U�� ����<dd=��=���<�г;䝛�L�:�����6ý ��1D�6��F�`P�cȽ�>��&XH�P����f; ձ<�   �   �G=��7=4��<Д1�����<�1�؂��2.�L�K�[����8ſ�������7C�0i�.}��<���U��\���[������F���Bh�**B� ��uq��$oÿ�)����I��^�h�����,�9p�������<��E=b�T=�S9=P =PEQ<����p���L=���x�h���5�nq���T��F�p�����0��R<��<b�+=�   �   �G=Tq0=C�<P���L��d�J�O��$����`�����wz׿J}��=/�f�W��
����s���Ը�W���ϸ�,ȫ��A�����D�V��F.���
�ֿ爞���^�y����>uG������4�<�8=��O=�:=�_=P�u<�d����żL?*�8�b�{ƃ�Hw��ׄ���f�D�/�D�Ҽ�һ�kW<�"�<�82=�   �   f�2=8K"=x�<|A��ڤ���dF�V������\��圿c�ӿ�-	��3,�z�S�8�~������>������������t��|~�ԲR�Y+�"f�U�ҿ�ڛ�D�Z����g��XQC������@���!�<�R*=�:=`~=lx�<ł;���*� �̶o�i���a����������6���ku�@�'��}���z;D��<և=�   �   ���<(~�<p!p<$^���j���>:������	�n�P��唿(|ɿ��Ɓ#��G�ZYo�}z������	}��y������cۜ�����o��}G���"����Suȿ�
���hO�f������~n7�䢤��<���:�<�d�<P��<`z�< �}��H����n�
������$��N������W����FS��Pw�R��7»�v<�   �    �c98*< ��;����ƚ�S�'�vb�������Y>��\��5.��-?�=�6�6��X�4�z��(���U��G	�����|s��&F{�"Y��6�2�n��}��� Ç��P=��-�����_%�؂��PE���L�;0cI<��;����&�T�AV����jd-���Q�ĉn������������p���S��/��V��%��.�]�i���   �   l�&�$厼p)<��6ڼ�	��as����g�پ��&�O�p�IY��S�տ�����!�D�>�(.Z���q��(���,��i��"�r���Z�l$?�x4"������տ8��&p��O&�Ęؾ[������j�� ̼�U����E�� ���s����7�|�s� e���ܱ�W�ƾАԾNvپ�վZ�Ǿ)���ژ���v��^:�^Z�Cٟ��   �   ��ƽ6{e���
w��|���󽏑[� ��>��ctL�����w����濂[�#�
9��qK�`�W�t�\�xX��DL��9���#����!S�P�������BL�=^�5]��/Z����Xv�dn	��P���]��v½p��e����Ǿ�;�_/��P�%���(��x%�6�����&���~ɾ!����h�����   �   �Y/��>۽�>�G�4o�Ʒǽ/�����|㾈�&��Vg�𛘿�T�����@��<e���'��1��4��1��`(��:�6���� �����f�g��&��"_���E.�7�Ž��j��&C�������׽2-�Vׁ��.��;��2/�� 5�n�O��yd�3�q���v���r��ie��P��G6�eg�E�p���F���   �   J���0�/��8ڽ���$�t�.ܢ����r^��������\6�W�r��V���Ż�T�ۿ����'�u������|���J���ݿ�⼿+��.t��7��O��V��hD^����
��|ir�o㋽��׽�].�����zHþA��^�-�`\W�zS�R��85��G%���X��Ă��Kܟ�T"��遀���X�T'/���)�ľ�   �   ô���e���!���Ž����=����Ľ�8 �Qy�����	���8��Om������.�������ӿ.߿�$�G�߿rԿ�¿�E���x��F�n��:���	�����*c���� �w�Ž�~���?��N�Ľ�< �R�J����!	�A�8�XTm�C����1��	�����ӿ�߿�(���߿�uԿD�¿�H��{��x�n� :�B�	��   �   �Q��Y��:H^������fgr��ߋ�[�׽}X.� ����Cþ$����-��WW�4N�O��2���!��MU�����1ٟ�y��\��+�X��#/�+����ľ�����/��3ڽj���
�t��ޢ�^��^�,�����`6�c s�rY���Ȼ���ۿ����)�6w������p��GN���ݿ\弿g-���t��7��   �   O�&�2�.a��0H.�6�Ž8�j�,!C�[�����׽t-�uӁ��)�����j+�7�4���O��td���q���v�x{r��de�D�P�MC6��c�I��{B��LT/��7۽������G�po���ǽ /�u���.#��&�>Zg����9W�������:g�֦'� 1�x�4�l�1��b(�|<�ܜ����X"��r��_�g��   �   �DL��_�A_���!Z�7���Xv��j	�"I�v�]� n½m� e��훾?�Ǿ�4�+��L��%��(�/t%� ���I ��yɾ{���Ih������ƽXpe����u�,!|�`��֔[����!���vL�n������!��
]��#�,9�@tK��W�(�\��zX�VGL�$�9�T�#�`��gU��Q��#����   �   p�%Q&���ؾ�������j��@̼�>�p�~�T8����rh��o|7��s�`��Fױ�8�ƾd�Ծ�oپ�վN�Ǿ}#���՘�\�v��W:��T��П�p�&�,Վ�8<�h5ڼu��4u�{����پ��&���p��Z��F�տ����!��>�\0Z�Z�q�A*��D.��rj����r���Z�&?��5"����?�տ����   �   �Ç�R=�N/�������`%�T���B��Pm�;�}I<�;�ߥ��T�OL��.���]-��Q�`�n�P���5��������o�&�S�n�/��P��� �]��Q�� (l9�#*<�ː;���\Ț��'��c������B[>��]���/���@��>���6���X�F�z��)��W���
��E����t��H{��#Y� �6��ġￇ����   �   ���iO�������o7�'���D:��$@�<|m�<���<|��<@"}�0���n�}z������8I�O�����R�S��K�� �v�������� v<��<���<0'p<,_���k��J@:�Ⱥ����	���P��政-}ɿZ����#��G��Zo�Q{������~��}�������?ܜ������ o��~G�^�"�,��vȿ�   �   �ڛ���Z�L��h��zQC������>���$�<�T*=T�:=v�=���<��;������ ���o�{���\�������z���1��"cu���'��p�� �;엱<&�=��2=�L"=�x�<�B��⥳��eF��V��o����\�-朿 �ӿ6.	�\4,��S��~������͛��W��}���������~�8�R�XY+�Tf���ҿ�   �   È��J�^��x�����tG�w��������<��8=�O=:=4`=��u<pb�� �ż?*��b�jƃ�Gw��!ׄ���f�x�/���Ҽ�һ�jW<"�<�82=��G=�p0=�A�<�Q��M��ˠJ����S��ƨ`�˥���z׿b}��=/���W��
�� ������Ը�W���ϸ� ȫ��A�����&�V��F.���
�Uֿ�   �   ڛ���Z����g��6PC������:���'�<�U*=Ĩ:=��=���<0��;����� �ʭo�����\��ɻ��{��2��>cu���'��p�� �;$��<d�=0�2=`M"=|{�<�>��7���TdF��U�������\�|圿�ӿ�-	��3,��S���~�?���������C��o���������� ~�:�R��X+��e���ҿ�   �   �	���gO���������l7����h2���D�<tp�<L��<h��< }��/��
�n��z��4��
�MI�c�����R�j��K��,�v�x�`����"v<̜�<���<@1p<0W���h���=:�踨���	���P�d唿t{ɿ@�(�#�2�G�:Xo��y��ƺ��|��u�������sڜ�5���Jo��|G���"���Xtȿ�   �   ����pO=��+�� �h]%�
��,7��P��;��I< 0;dޥ�܂T�PL��9���]-��Q�}�n�]���D��������o�6�S�z�/��P�����]��P�� tm9�,*<P�;����Ú���'�Ma�������X>��[��)-���=��<��6���X�P�z�m'��oT���������Kr��D{�d Y���6�,�͞�/����   �   �p��M&�)�ؾ{���}��e��(̼�.���~��6�J��Sh��r|7��s�*`��Vױ�L�ƾx�Ծ�oپ�վ`�Ǿ�#��֘�`�v��W:��T��П��&�Ў��<�(ڼD��.q�l��X�پ^�&�T�p��W����տ���<�!���>�,Z�^�q��'��l+���g����r���Z��"?�3"������տ����   �   @L�R\�lZ��"Z�����Mv��c	��D���]�Lm½?��e��훾I�Ǿ5�+��L��%�(�(�9t%�)���R ��yɾx���0h�ò��ƽ�me�0���m��|����A�[�������/rL�K������N�� Z�n#�9�|oK���W�Ɣ\�ruX��BL���9���#�z���P�N������   �   ��&�=�X\���A.���Ž�j�C�+���b�׽-�`Ӂ��)�����o+�@�4���O��td���q���v��{r��de�L�P�SC6��c�G��^B���S/�Y6۽c���p�G�o�9�ǽ�/�����-�E�&��Sg�
���QR��Խ远��Vc���'�r1���4���1��^(��8�t����r��p��	�g��   �   @M�6S��?^���Q���\r�n܋�L�׽�W.�؀���Cþ#����-��WW�=N�O��2��"��RU�����5ٟ�|��^��-�X��#/�&����ľ⠇�"�/�d1ڽ����@�t�y֢�#���^������
Z6���r��T��+û�5�ۿq���%�s�r����~��	G��< ݿ�߼��(��$t��7��   �   �����_���� �׌ŽMx���8����Ľ8 ��x�����	���8��Om������.�������ӿ4߿�$�N�߿#rԿ�¿�E���x��F�n��:���	�а���b���� �^�Žz��8���Ľ�4 ��s����3	�<�8��Km�!���,��{�����ӿ ߿$!㿋�߿�nԿ��¿�B���u����n��:���	��   �   T���$�/��*ڽp���B�t� آ�P���^��������\6�X�r��V���Ż�W�ۿ����'� u������~���J���ݿ�⼿+��+t��7��O��V���C^�������v\r��ً���׽~S.��}��-?þ=����-�nSW�)I�AL��/�����R��>|��֟�����|����X��/�����ľ�   �   *N/�T.۽G���4�G�po�N�ǽ�/�����X㾁�&��Vg�񛘿�T�����D��<e���'��1��4��1��`(��:�6���� �����c�g��&����^���D.���Ž&�j�lC�ᮃ�K�׽�-��ρ� %������'��4��|O�|od�L�q�n�v�vr�a_e�f�P��>6��_���|>���   �   #�ƽ,ae�j��8j�R|��󽼐[����2��btL�����{����濄[�#�9��qK�b�W�x�\�xX��DL� �9���#����"S�!P�������BL�/^��\��VZ�+���Ov�|a	�v>��]�9e½����d�雾��Ǿj.��'��H�u%���(��o%� ��D�y��-sɾ����bh�����   �   ��&�������;�D#ڼ���Zr����?�پ��&�Q�p�LY��U�տ�����!�F�>�*.Z���q��(���,��i��"�r���Z�n$?�z4"������տ8��%p��O&���ؾ����~�9g��t
̼H���~� +����]���u7���s�O[���ѱ�G�ƾ�Ծ^iپ)վ>�Ǿ����И���v��P:�O��ǟ��   �    �v9�F*<��;���xĚ���'�Ab��p����Y>��\��8.��/?�=�8�6��X�4�z��(���U��G	�����}s��&F{�"Y��6�2�p�����Ç��P=��-��f�_%�����(7����;X�I<@�;�ǥ��sT��B������V-���Q�Cyn��������F�����o�x�S���/��J�����]�`7���   �   ���<l��<�;p<U��i��w>:������	�m�P��唿*|ɿ��Ɓ#��G�\Yo�}z������	}��y������cۜ�����o��}G���"����Uuȿ�
���hO�`������n7�a���l3���G�<�v�<���<ș�<��|������n�_r�������C���P���M���潄B��P�v������ Cv<�   �   T�2=�O"=�~�<�<�� ���zdF�V������\��圿c�ӿ�-	��3,�|�S�6�~������>������������t��|~�ֲR�Y+�"f�V�ҿ�ڛ�B�Z����g�� QC�����@<��8(�<�V*=�:=��=X��<�!�;t{��H� ��o�����W�������u��-��Zu�L�'�b���5	;`��<z�=�   �   >>=�%=���<4/Ƽv�ŽP�U�斿�V&�ݰi�0���mi߿*���"6�na��q��q���u1��a���G`��)����%��I|���E����`�j�5��I�$�޿�G�� i�\���Ⱦ��}T��ý����D��<h-)=�HA=��*==�<�)<X�!�I���D� 
~�Ҩ��?9����H��x8F������-���<���<��'=�   �   �2(=H@=�K�<05Ǽ;����gQ�ʻ��7���e�a颿Ȼۿ�B���2��\�]����������Y��
����[��o	����hh���f\���2�^���1ۿR|����d�÷�����)P��п�`տ��'�<J�=�v+=lf=�j�<�V��T[���:�������1��������,���尿�.��V�=�VƼ�c캼�<x$
=�   �   �j�<ē�<H�6<8�̼b��*�D��԰�Ļ�YY����R
ѿ�]���)�B�P�|�z�D���=6��꫱�G��۷���C��b�����z�FQP�\�)�� ��п X����X��K��"����C�zp��<�ż8�C<��<p��<��J<Xn��?�~(��:,����������O�n
"� ��4U��8��~�½͇�d�� 	%��)=<�   �   �v�`N�;�:� ݼxU��b�1���"���XF��̍��H��fT����N>���b�=���8����f��/J���|��K���C����b� J>����2�����#���@�E�6�
_����0�ᙦ���ּ�ɬ:���;��@���ּ
�q�%�Ƚ���9�Q�^�,R|���������ꇾ��|��U_�v�9���ʽ`mu�,�ݼ�   �   ��<�薴�lW���l�+���������{8.�j�z��٪��4޿��
�\t(�`�F��_d���}�g���vي��ˇ�
5~�µd�PG���(���
��&޿㻪�laz���-�v�Ă��������������x��^���F9�6������6�C�&)��tȟ��3��N�о��޾���1/߾XѾ�����[��������D�e�	��c���   �   *�ս��}�6f"�,%�����h���g�����&�8U�zb���f��+�￢��4�)��A�T�
�a��f��b���T�blA�J*�~#�������d���"U���=���>g�t������f�"�X���z�)Խ@H'��s�������Ѿ"@�����ׂ"�V�,��0��,�P�"�6:������Ҿ�O���Pt��O(��   �   N�9�MB뽯����_��K��R~׽w�9�EH������$.��Eq�O�ȿ���U����J�.�؆8��<�v�8���.�	 ����a��pȿ���uq�}4.����,���z9�]�ֽ�t��� ^�J���4��A�8�=n��"俾h����j�6Z=�N�X�-kn��D|����!z|�I�n�/HY��=�c��{���2���z����   �   f���΂:����C=����������;���j�򷾱�1�>� �}�Oՠ��~ÿS��� �"������� ;����V8�)!�Y�ÿ�*����}���>��@������j�p,��@����D��������9��/���k;�J���5��a��;��}��L̥���$���������З�1����a�Dy6�n���ξ�   �   �ʾ7@���7+�o�ս�b���H���:ս,�*�r�����ʾZ���aA���w�����YS��e�ɿWܿ���������bܿ�"ʿ6Ĳ�A ��fcx���A�#�(�ʾ}=��t4+���սb��zJ���?սH�*�������ʾO��ieA�*�w�o���zV��ܴɿ	ܿ���������vfܿ�%ʿ6ǲ��"���gx�L�A����   �   2C����� k��.�PB����~��������9��+���f;�G���5�a��8��z��ɥ�[﮿!��I�����Η�������a�|u6�j��%ξ���9~:���}:�����������>���j�����-�}�>�1�}��נ�Ӂÿ����� �6�������,=����.:�l$�+�ÿ�,����}���>��   �   �6.���3.��}9�x�ֽet��6�]�퍒����N�8�2j���޿������f��U=�>�X��en�?|�<���zt|���n�>CY���=����H���J��������9��:�?���P�_�YL����׽��9��J��q��x'.�Iq��񞿎 ȿ��W������.�X�8��<��8��.� �p��L��rȿ�!��xq��   �   +%U����a����@g����������"�>��,�z��ԽB'��s�t���t�Ѿ9������~"�Պ,�0���,��"�S6�����Ҿ�J��It��I(���սX�}��_"��)%�⊽:���g�F����:U�7d���h�����8���)��A�Z�T���a���f�Tb�r�T��nA�*��$��𿷁��'f���   �   tcz��-�x�������/���p����x�`K���89��v�����ƺC��$��>ß��-����о&�޾��㾐(߾�QѾڰ���V��R�����D���	� [��6�<�\���dN���k��,������􊾘��R:.��z�*۪��6޿�
��u(�N�F�8bd���}�汇��ڊ�Q͇��7~���d�G��(�� ��(޿=����   �   򎍿o�E��6�`����0�]���\�ּ P�:`�;�'@���ּh�q�ةȽ��l�8�L�^�vI|�F�����懾c�|��M_���9�
�W�ʽ�]u�,�ݼ`�u�`{�;��:` ݼ
W���1�0���C��&ZF�	΍��I�� V����tO>�N�b�Z�������h���K���}������E�����b�RK>�����������   �   �X��N�X�/L�W#��I�C��p���ż`�C<�%�<��<ذJ<�C�3�� ��Y#������p��HJ��"�����O�=/���½�Ň�:��X�$��G=<Xu�<h��<�6<8�̼wc����D��հ����XZY�P���_ѿX^���)�\�P���z�(���?7������X��ั��D��(�����z�&RP���)�!�֞п�   �   �|��<�d�������)P��п�lӿ�+�<��=
z+=�j=u�<����\L��n�:�����ܶ��Y����'���ꦽ�)��V�=�dHƼ��뺼��<�'
=<5(=�A=@L�<�6ǼJ����hQ��ʻ�8�m�e��颿h�ۿ�B�d�2���\�ʋ������T��1Z������\���	��k���h���f\���2����2ۿ�   �   �G����h�+���Ⱦ�4}T�]�ýH������<�-)=FIA=�*=�=�<X�)<�!��H��DD��	~�����=9����n���8F������-�`�<,��<B�'=�>=��%=Ж�<�0Ƽ
�Ž��U�-����&��i�U����i߿B���"6��a��q�������1��i���G`��#����%��;|���E��b�`�N�5��I���޿�   �   �{��0�d�3������(P��ο�4Ͽ��-�<��=�z+=�j=Du�< ���xL����:�,�����ﶺ�m����'��립*��d�=�lHƼ@�����<,(
=�5(=xB=�N�<�2Ǽ����,gQ��ɻ��7�]�e�+颿{�ۿRB���2�t�\��������J��Y��z���[���������g���e\�2�2����1ۿ�   �   2W��N�X��J�m!��ȺC��m��Жż��C<�(�<��<вJ<(C��2�� ��n#��������aJ��"����P�^/���½�Ň�*��x�$��I=<Hw�<���<ȩ6<�̼=`���D��Ӱ�6��RXY������	ѿ4]�0�)�`�P�J�z�~���Q5��媱�7��˶���B�������z�0PP���)����п�   �   �����E��4�`]����0�蕦��ּ@��:�+�;�@�P�ּ�q�ҩȽ��~�8�b�^��I|�U���+��(懾��|��M_���9�
�P�ʽ�]u���ݼ�uu�Ќ�;��:ݼ�R����1���H��YWF�$̍�G�� S�����L>���b�:������Ke���H��<{�����(���J�b��H>������t���   �   �^z���-�js�Ӏ�����᭖��
����x�TF���79��v�����ĺC��$��Iß��-���о<�޾ �㾧(߾�QѾ鰻��V��Z�����D���	��Z����<�D����E���d�?'�����g�����6.�]�z�5ت�3޿��
��r(���F��]d�0�}����׊�\ʇ�P2~�l�d�fG�,�(�h�
��$޿L����   �   = U���\����9g�3������0�"����z�z�Խ�A'��s�t���{�Ѿ9������~"���,�0���,��"�\6�*��� �Ҿ�J��It��I(��ս��}�["��"%�X܊��|�A�g�8���{��5U��`���d�����.��n�)�~
A�F�T�H�a�6�f��b�`�T�"jA�d*��!���}���b���   �   �1.����,)��=v9���ֽ�n����]����������8�j���޿������f��U=�J�X��en�?|�C����t|���n�GCY���=����I���A���������9��9�񳓽��_��F���x׽��9��E��1��x".�nBq�Wힿ}ȿ��T����
�.�f�8�n<���8���.� ���B��|mȿb���qq��   �   x>�%���j�D(��9������
���Ր�0�9��+���f;�G���5�a��8��z��ɥ�c﮿!��Q�����Η�������a�|u6�f��ξᜎ��}:��}��6��|��/���&8��j��p�3�>�0�}��Ҡ�	|ÿ��<� �����b���8����n6���_�ÿ(����}���>��   �   ��ʾ!:��l/+��ս/[���C���7ս:�*�.���y�ʾT���aA���w�����]S��l�ɿ_ܿ���������bܿ�"ʿ;Ĳ�C ��hcx���A���ʾ:=��|3+���ս]���B���3ս��*�s�����ʾ���!^A�0�w����_P���ɿ�ܿ�����(��_ܿ(ʿ�������^x��A�)���   �   3���lx:�w�H3��{��ǌ��d:��j��񷾥�,�>��}�Qՠ��~ÿX��� �&�������;����X8�,!�\�ÿ�*����}���>��@������j�+�n<��b���@��� �齜�9�](��b;�D�.�5�}a�<6��&w���ť�쮿������a	���ʗ�Ռ��ȡa�|q6�+���;�   �   ��9�I1뽥���z�_�5F���z׽^�9��G��v���$.��Eq�P�ȿ���U����L�.�܆8��<�z�8���.�	 ����e��"pȿ���uq�t4.����+��jy9�ǽֽ6o��$�]�=���-�齆�8�bf���ٿ�����,c�SQ=�[�X�h`n�x9|�b����n|���n�6>Y�$�=����������������   �   ��ս��}�S"��%��܊��}���g�_����8U�|b���f��.�￤��6�)��A�ğT��a��f��b���T�dlA�L*��#�������d���"U��� ���@=g�	������"�0��<�z��Խ
<'��s�������Ѿ>2�����Xz"�f�,��	0��,�Ͼ"�a2�����Ҿ�E���@t��C(��   �   ��<� n��$:��pb��'����������r8.�i�z��٪��4޿��
�^t(�b�F��_d���}�h���xي��ˇ�5~�Ƶd�RG���(���
��&޿绪�laz���-��u�t������Z���,	���x��5��.+9�
n��	����C�g ��>���(����о��޾>���!߾sKѾ���cQ��޶��f�D���	��Q���   �    �t�P��;��:�ݼS����1������XF��̍��H��gT����N>���b�>���9����f��/J���|��K���C����b�"J>����5�����#���=�E�6��^��<�0�v����ּ �:0X�;`�?���ּ��q��Ƚ����8��|^�A|�θ������ᇾ��|��E_�p�9����ʽ�Lu�Ծݼ�   �   ԃ�<���<x�6<ؚ̼�`����D�f԰����YY�����U
ѿ�]���)�B�P�~�z�D���<6��쫱�G��ܷ���C��c�����z�FQP�\�)�� ��п X����X��K��"��2�C��n��ԗżP�C<\/�<d�<h�J<���&�������h���C���D�'�!����J�r%��+�½���@��h�$��j=<�   �   �8(=�D=R�<�0Ǽ~���RgQ��ɻ��7���e�b颿Ȼۿ�B���2��\�]����������Y��
����[��o	����gh���f\���2�^���1ۿU|����d����q���)P��Ͽ��п�|.�<ޓ=�|+=Nn=H~�<�Յ��>����:��������������y"���妽O%����=��9Ƽ ��`�<X,
=�   �   �5?=`�&=<��<��ļǇŽ��U��ʿ��X���i���g�߿@��~w6�,�a�����E�����ɡ���L��$���v��gX��Z����a���6�H����A��pvj�����G���V���ƽh�Ǽ.�<B�%=�1>=��'=���<�+<�S0�З����G�S���;���Z���ߒ��G���F� ?���y+��� < ��<��(=�   �   NV)=�W=�0�<��żC���6�Q�� ���l���e�$��-ܿN{��P3��Y]���i�������B��D���A��Z������_����]���3�����hܿ�m��Ef�e���x��7R���½@�ȼ�͊<�F=�H(=�!
=�<�
��(ȼ��>�0������R���Cýc��5���Ro��ʨ=��wż�6Ժ�<l>=�   �   �l�<���<��9<��˼fZ���E���������Y�?���4jѿd��@L*�D+Q���{��i�������������R��Jg����{�LQ�u*�Z��)�ѿk2��#Z�7>��|����E�0@��\[μ $5<tE�<��<��;<Hu'�ʡ�������ý�f��,�4Z���"�p4�B��W����½������H�!���@<�   �   @	j��(�; r6:�xܼCi��w2�;������F����W����������d?���c��P��?R��:������*�� <���=����c�l?�����$������G���
G��	�������2�3���߼ ��9���;�4� �߼�v���˽�����:��@`���}����������f��\�}���_��(:�V"���ʽ��t���ܼ�   �   PR<��ֳ��Ɓ��b�Rb�����E������.��]{�i]���޿�y��+)���G���e�*B�sc��~z��xP��@��\e���G�)�,r���޿�o���{��.����4���Zz�J��������Do����=�X9��vi
���E�>��`����l��-&Ҿ������߾�Ѿ���Q���`���N�D���	��E���   �   �ֽ�~� �"�$�%��C�����C�h�p���=����U��풿)�����P��V�*�B��U�|�b�آg���b�ƃU���A�`l*��t����i���钿lV���ƿ���h��*�yɋ���&���#��q�c�ֽ�)�Bu�쥾�Ӿ����l���^#�@Y-�=�0��>-��.#����4f����Ҿ�y����t��l(��   �   ��9�E��o����`�9䄽Voؽ��:��陾���.�Wr�x���Aɿ�U���� ��/��[9��<�`;9��L/��L ��������ȿ����1r�+�.���t����:��ؽ9E��X�a�Ȯ��v콴y:�p����N������s���>�LZ�U�o�^}�����7}��Yo�2�Y�"&>���*������.���   �   �펾��:��W�8��7]��ͱ��f�d(l�J㸾�����?���~�����-�Ŀ���V���=�.���E����`�j�9q忛<Ŀ�s��l�~�S_?�s���Ƹ�l����Բ�g���,Y��}��b;�#7����ξ>4��7�glb�M���O����������ò�D���k��>���Å�s�a��6�h��fξ�   �   �|˾���z�+�Z�ֽ7���=���<�ֽ^,��ׇ�s�˾�����B��8y�᝘�4T��q�ʿ�ݿ��������ܿFsʿ����V����x�)0B�~R��x˾T�����+���ֽW�������ֽy,��ڇ���˾���P�B�Z=y�����XW����ʿݿ���մ���近�ܿ�vʿ���GY��8�x��3B�3U��   �   ����ɸ�l���ֲ�]���hU������\;�l3����ξ�0��7��gb������L��`���&�������䐯��g��J��?�����a�F�6�d��maξ�ꎾY�:��Q�m���]��o���?� -l��渾R���?��~�����.�Ŀ��B���?�d�� H�Ơ�j��k�}t�m?Ŀv��C�~�Pb?��   �   ~�.�I������:� �ؽ�D��Ϊa�o����m콺s:�a����I��_����o��}>�6Z�ؘo�VX}����2}�$To�@�Y��!>����#������P*��,�9������>�`��䄽�rؽ2�:��왾���-�.��Zr������ɿ�X���� �n�/��^9���<��=9�2O/��N �\�����!�ȿ����4r��   �   �V����)ȿ�O�h�-,��ɋ��&���#��d��ֽ��(��9u��楾�yӾv���k��cZ#��T-���0�D:-�`*#���R_���Ҿ�t���{t�g(�o�սl�}���"���%��D�������h����/����U��,+��c����>�*�LB���U�Rc���g�Z�b�H�U���A�*n*��u����T��]뒿�   �   )�{���.����h����{����������[����=�0��wc
�)�E��9��"񠾱f���Ҿ
�P��R�߾��Ѿ���B���܁�6�D�1�	�=���E<�Ƴ������a��c����%G�����β.�g`{�_��!�޿4{�`-)���G�R�e��D��d��	|���Q�����^e���G�t)�Ds�v�޿�p���   �   RH��G�Y
�������2��3��\߼ ��9���;��~�؍߼ �v�V}˽ʤ�ȩ:��8`���}�|��X���>b����}��_��!:�h��}ʽ��t��ܼ�i��U�;�)7:�xܼ�j��22�{<������F�������]���Ȍ��?�~�c��Q���S��z;�� ��G,��9=���>��L�c��?�~��&�������   �   �2���Z��>�;}��,�E�~@�� Yμ /5<hN�<T(�<�<<�J'�����{���ý�\�����T�F�"��.��������u�½g�������!�XA<8w�<p��<��9<��˼�[��TE�������Y����=kѿ��M*�`,Q�b�{��j����� ����������A��h����{��LQ��u*�����ѿ�   �   -n��hEf�����x��>7R���½l�ȼ4ъ<I=(L(=�%
=���< >��ȼB�>�c����觽'M���>ý��8{���j����=��iż�Ӻ�<�A=�X)=DY=d1�<h�żM���(�Q����%m���e��$���ܿ�{�DQ3�zZ]�z����@��C�������A�����d�������]��3����9iܿ�   �   �A��3vj�O��hG����V��ƽ��ǼX/�<��%=h2>="�'=l��<x-<�R0� ���d�G�>���1���Z���ߒ��G��H�F��?���z+�h� <P��<d�(=�5?=��&= ��<��ļY�Ž�U�%˿��X� j�#󥿒�߿X���w6�J�a�����E�����ϡ���L�����j��WX��I����a���6�.����   �   wm��WDf�վ��w���5R���½�ȼ�ӊ<�I=�L(=,&
=艖< =��4ȼV�>�t����觽@M���>ý/��R{���j��ؠ=�jż@}ӺL�< B=*Y)=Z=4�<(�ż����֊Q�� ��el���e��#���
ܿ{�xP3�fY]�������5��B������w@�����z��������]�<�3�$��Lhܿ�   �   �1���Z�P=�L{����E�;=���Pμ895<�Q�<0*�<0<<�I'�����{��"�ý�\�����T�^�"��.���˨����½x�������!�`A<y�<���<��9<��˼�X���E�/�����Y�����{iѿ���K*�d*Q���{�i�����菲��������O��gf��N�{��JQ�0t*���� �ѿ�   �   mF��B	G�_������2�$/��߼ ��9 ��; �~�d�߼Ҥv�N}˽Ѥ�٩:��8`���}�|��h���Pb���}�%�_�":�r��}ʽ��t�|~ܼ@ki� g�; 8:�mܼbf���2��9��
����F�*��C���?���ʊ�2?��c��O��Q���8��G���)���:��|<����c�?�~���"��k����   �   ��{�/�.���>���iw�o��4��$
���V��2�=��/��bc
�%�E��9��.��f���Ҿ
�g��i�߾��Ѿ��N���܁�7�D�!�	��<��jD<�����@���>[�{^��r��C��ۅ�v�.��[{�\��g�޿�x�r*)��G�e��?��a���x���N����`Ze��G��)��p���޿�m���   �   � V���ÿ���h��'��Ë�ȅ&��#�.b�P�ֽJ�(��9u��楾�yӾ����t��oZ#��T-���0�Q:-�l*#���`_��&�Ҿ�t���{t��f(���ս��}� �"��{%�4?����ӈh���������U�X쒿'��b��ܚ���*��B���U���b���g���b�.�U�v�A�xj*��r����@�� 蒿�   �   |�.��󙾴�:�'�ؽ?��`�a�!���Ul�Ys:�H���|I��_����o��}>�AZ��o�cX}����+2}�2To�L�Y��!>����#������;*����9���뽮����`�߄��iؽ^�:��百=��*�.��Sr�}����ɿ�R���� �ԁ/��Y9���<��89��J/��J ��������ȿۄ��.r��   �   ��(ø��l�r��Ͳ�А���Q�����6\;�B3����ξ�0��7��gb������L��e���-�������쐯��g��O��D�����a�I�6�a��]aξpꎾ��:��O������W��諲��
��#l��߸������?��~�����^�ĿY��~���;����C�j��L�.h��m忟9Ŀ5q��>�~�\?��   �   t˾������+�»ֽ����=����ֽi,�:ׇ�P�˾�����B��8y�❘�9T��x�ʿ�ݿ���� ����ܿMsʿ����V����x�+0B�yR�~x˾���	�+���ֽW���^���`�ֽ�,�~ԇ�Z�˾�� B�U4y�H���7Q���ʿݿA�����9��4�ܿ�oʿ�����S��=�x�`,B��O��   �   �掾��:�I�2����V��x�����'l�㸾�����?���~�����0�Ŀ���X���=�2���E����d�j�=q忟<Ŀ�s��o�~�O_?�g���Ƹ�Rl�J�7в�����O����뽜W;��/���ξ�-��7�cb������I��/���ͨ��5��������d��E������%�a�G�6�%��Z\ξ�   �   ��9�7��X��b�`��ބ��kؽ�:��陾���|�.�Wr�y���Bɿ�U���� ��/�\9��<�d;9��L/��L ��������ȿ����1r�%�.����%����:�l�ؽ�?����a������d��m:������D��'����k��y>�L�Y���o��R}�����u,}��No�8�Y�9>���M��V���2&���   �   x�ս��}��{"��w%�`?��J��f�h�5���0����U��풿)�����R��V�*�B��U���b�ڢg���b�ȃU���A�bl*��t����k���钿iV�ٞ��ſ���h��)�ŋ���&�l�#��V���ֽ��(�92u�"⥾�sӾ�������.V#�IP-�"�0��5-�&#��{�EX��	�Ҿ�o���st��`(��   �   �6<�ԭ�������X��^����0E��և��.��]{�i]��!�޿�y��+)���G���e�,B�tc���z��yP��B��\e���G�)�.r���޿�o���{��.����䃋�Hy����T��0��@F����=�'���]
�
�E�@5��젾a���Ҿvྞ�侺�߾��Ѿ/
������ׁ���D�&�	�k3���   �   ��h����; 9:hjܼ�f���2��:������F����Y����������f?���c��P��@R��:������*�� <���=����c�n?�����$�������G���
G�	�t���Δ2��0��� ߼ ��9��;��}��t߼<�v��s˽���:��0`�f�}��w��Ŷ���]��$�}��_��:�G��sʽ �t��dܼ�   �   ���<d��<�9<8�˼�X��tE���������Y�@���5jѿf��@L*�F+Q���{��i�����퐲��������S��Lg����{�LQ�u*�\��+�ѿj2��#Z�/>�u|���E��>���Qμ?5<DX�<�4�<�%<< #'�����t����ýS�����O���"�M)����ڞ����½�������h~!�X8A<�   �   d\)=v\=D7�<P�ż������Q�� ���l���e�$��,ܿP{��P3��Y]���h�������B��D���A��[������`����]���3�����hܿ�m��Ef�c���x���6R���½��ȼ�Ԋ<4K= O(=�)
=ܒ�<����l�ǼB�>������㧽 H��;9ý���/v��f��B�=�[ż��Һ���<JF=�   �   H�K=�B4=|��<�c���̶���J�ិ��_� �a��R���bؿP �l=0�@HY�:c��<o��lG��[x��f
���|���_���������"&Z��1����ħٿ�Q��>"c�
��mS����M�-㺽������< �.=pPF=N�0=���<>L<��fۼ��4���l�l����������li���0��]Ѽ�û@�b<�
=6=�   �   ��6=�%=8�<D���@8��4�F�=���x����]������ԿH�	�0C-�>AU�!������0V���;��<����6���^��N0��D�����U��.���
�ֿ�u_���g���ZHI��4��������<�V =X�0=��=|��<�©:X���F�,�^4{��u����� n����zŚ�d�v��Q'�LD��@+2;�)�<�<=�   �   �Z�<��< d{<䀢��2����:�	p��-f
���Q�ط���ʿ�N�x�$�
�I��.r��l��D����u/��G�������d��ar�d<J��9%�����˿5{��ES��X�g檾=��笽�6��8d<l��<L��<P�j<��޻Z��4�|�Y������W�	�NT���p�����3轷����4v�|#� (��u�<�   �   �}_:�=4<�١;�z���ߚ��v(�24���q����?�O������'�����8��[�І~�&^��:����9��'w��9��N~�:�[��8����ղ�@���։��@������g���j*�6*��9����i;�a<�c&�l���Rc�(���b~	�1B2�N�V��Ns��Ȃ�?υ�$o��r�"�T��S0���C���z\�е���   �   "\%������{7��aټV���Q�^���j�۾[(���r�gܥ�ؿ�<��#�\FA�F�]�~�u�=��Y���_����u���\�H�@���#�2&��'ؿ7��is�
�(���ܾ兾����T��@����L�������+��#���x��=�}	z�qΚ�$d��d]ʾ��׾�(ܾ�>׾�}ɾ4?��Q���yw��:�4O��^���   �   �ǽ��e�z��6�V&~�	��Z�]��ݷ�k �ܥN�e0��B�����ZN�jz%���;��N�
	[�nB_��Z�\�M�;���$�����#�5���&����N��b�t���^�QM���K��r��v ��xk�y�ʽq-!��Ik�Բ����˾	��T��v���`'�n�*�'��-�����Q��%CʾD,��_�h����   �   ("0��mܽ����EJ�fZr�_eʽ.D1��u��J���(��kj�Ÿ��ÿ�H���	�����$*��v3�ؒ6��3�Xx)��	�PH	�u3�Ra¿�G����i�ʤ(���ᨓ�n�1�X�˽�u�HN���Y߽�	2�\��/E�������&��Q8��S��g��'u�͇y�S�t��g�!�Q��(7�r�6��|����΃��   �   4���	`1���ܽҿ����y� ��
:���a�௱����t-9�C�v�Μ��о��:߿�����	�RA�$�������?���& ޿Kʽ�=
���u�Ň8�^��rU���oa��N�����Ȗ{�����v޽Q�2����;KǾ#c�Q#1�CJ[��ၿ��������pE��&���奔l�쒿�����Y���/�zu���ž�   �    CþC���
#��ɽW닽T ����ɽѲ#��6���,ľՌ�i(<�:pq�z���
����ĿD�ֿ����w�:S��տ�ÿ�
��s"���	p�� ;���
�)?þ�����#��ɽwꋽ"��Q�ɽɶ#��9���0ľ���,<��tq�(������Ŀ�ֿV���{��Vῦ�տb�ÿ����$��p�$;���
��   �   ���rX���sa��P�'���{�:��3p޽F�2�Y|��\FǾ�_�f1��E[�߁� ���y���B���"��d쩿O렿꒿��k�Y�G�/��r�|�ž󀈾�[1��ܽ���D�y�����<�2�a�Q���H���09�X�v��М��Ӿ�7>߿���� 	�tC�N���� ��ԃ��S޿ͽ������u���8��   �   �(��������1�o�˽4�u�� N��ꉽ�Q߽�2�k��@��5���*#��M8���R���g�"u�,�y�Ҩt��g�V�Q�G$7���1�������ʃ��0�wfܽ����BJ�|[r��hʽBG1�x��澣�(�"oj�纚�� ÿ�K쿖�	����"'*�y3�H�6��3��z)����I	�K6뿱c¿�I����i��   �   !�N�Qd�7v����^��O���K�������lk�t�ʽZ'!��Ak�䭟��˾���q��C��J\'���*��'�)����J��x=ʾ�'����h�����ǽ�e�&�X4�z(~������]�0෾L"�r�N�2��D������O�B|%���;���N��[�,E_���Z���M� ;���$���&���((���   �   ks�z�(���ܾC慾���U��T�㼀�L�����p�+�����r��=�� z�Yɚ�l^��0Wʾz�׾-"ܾd8׾|wɾ�9��k����pw�%�:��I�8V��P%�l�i7��_ټ�����R�� ���۾�\(��r��ݥ� ؿ>���#�2HA���]��u����������8u���\���@�L�#�B'�F)ؿ����   �   �׉�?�@������h���k*��*���5���%j; |< $��꿼�Bc����^x	�5;2�x�V�lFs�MĂ��ʅ��j����q���T�(M0��y�÷��P�[�������a:�S4< �;|z��ᚽ9x(��5��"t����?�P������(���V�8�ȿ[��~�^_�������:��sx��`��>~���[�>�8����3��O���   �   �{�� S�Y�窾�=��笽�4��H)d<8��<���<��j<�y޻���.�|�����/���	��N�]�� ����p*�g���t&v����ܫ����<e�<��<Pj{<ȁ��=4���:�(q��g
���Q������ʿhO�F�$��I��/r�am��:��	��}0��C�������e��.br�>=J�v:%������˿�   �   %����_�1�������HI��4��D󩼸��<Y =��0=ԓ=���<���:����ܒ,�+{��p��d����h�����������v��I'��6����2;�2�<
@=D�6=\�%= �<����:9���F��������H�]�����I�Կ��	��C-��AU�����N	���V��<��ɵ��x7��"_���0������<�U�&.�̐
�jֿ�   �   Q��"c�܂�'S��9�M��⺽<����<��.=�PF=��0=x��<H?L<0��0fۼ��4���l�T����������li�&�0�(^Ѽ�ûP�b<�
=�6=��K=xB4=T�<,e��bͶ��J�%����_�:�a��R��cؿh ��=0�^HY�Kc��Ko��wG��bx��h
���|���_����������&Z��1������ٿ�   �   s����_�u������2GI��2��塚x�<�Y =�0=�=��< ��:�����,�$+{��p��{����h��	��������v�J'�7��`�2;�2�<L@=��6=$�%=��<�����7����F�����F��B�]�圝�f�Կ�	��B-��@U�ڰ��t���U��;������d6�� ^���/������0�U�`.�6�
��
ֿ�   �   jz��S��W�'媾1=��䬽�,��x3d<T��<���<P�j<�w޻���4�|�����H��,�	��N�x��������*轇����&v���0۫����<�f�<t�< t{<�y��1����:�Jo���e
���Q�Q���b�ʿRN�޶$�6�I�n-r��k��d����n.��A������d���_r�X;J�9%�|��݊˿�   �   �Չ���@�����f��Ah*�T&���*�� ^j;��<��#�l鿼6Bc����`x	�C;2���V��Fs�\Ă��ʅ��j����q���T�>M0��y�÷���[�`��� �a:0\4<�;�o���ܚ��t(�3��Rp��ʛ?�:N�������%����8���[��~� ]����@8���u�����4~���[���8����'������   �   �fs�6�(��ܾ.ㅾ����O�� ����L��{����+�n���r��=�� z�dɚ�z^��BWʾ��׾C"ܾ{8׾�wɾ�9��z����pw�+�:��I��U���N%�xꋼ�Y7��Rټ�����N�����W~۾�Y(���r�ۥ�gؿ�;���#��DA�4�]��u��������ނ�&u�^�\�r�@�z�#��$��%ؿ����   �   L�N��`�Kq�� �^��F��!F����� �Zik���ʽ '!�~Ak�⭟��˾���y��M��W\'�
�*��'��)�*���J���=ʾ�'���h�����ǽJ�e���<-�R~���� �]�J۷�����N��.��)@������L��x%���;���N�l[��?_�j�Z���M��;� �$���7!����$���   �   .�(������B�1���˽ƅu���M�=艽.P߽s2�P��@��3���-#��M8� S���g�*"u�<�y��t��g�b�Q�R$7���8�������ʃ��0�,eܽ�����:J�2Pr��_ʽ�@1��s�������(��hj�ڶ���ÿ
F�$�	�����"*�Xt3�l�6�B3�v)����F	�l0��^¿�E��x�i��   �   ���Q���ja��J�Ө����{����n޽��2�,|��DFǾ�_�f1��E[�߁����}���%B���"��k쩿W렿꒿��r�Y�L�/��r�n�ž̀���Z1���ܽ������y�a���6��a���������*9���v��˜��;��7߿F���	�<?���������|����ݿeǽ�����u���8��   �   �:þS����#�>ɽ�㋽i����ɽܱ#��6���,ľ̌�g(<�;pq�{���
����ĿK�ֿ���x�CS�"�տ%�ÿ�
��x"���	p�� ;���
�?þX����#��ɽ�勽�����ɽ|�#�4���(ľ,���$<��kq�� �����]�Ŀ��ֿ���1t�{Oῃ�տ��ÿ������Mp�;��
��   �   3}���U1�ezܽ���l�y�����8�Ψa��������m-9�A�v�Μ��о��:߿�����	�VA�*������G���, ޿Pʽ�@
���u�Ç8�R��?U��oa�tM�_�����{���~h޽*�2��x���AǾ]��1�)A[�܁�"���\����>��i��驿+蠿 璿c����Y�h�/�go���ž�   �   �0�]ܽY����5J��Or��aʽC1��u��!���(��kj�Ÿ��ÿ�H���	�����$*��v3�ܒ6��3�Zx)��	�TH	�x3�Va¿�G����i�Ĥ(��澔���^�1���˽�u��M��㉽I߽/�1����<;��'�����LI8�3�R���g��u��|y�T�t�rg�u�Q��7����󾟦���ƃ��   �   �ǽe����)��~�C���]�_ݷ�\ �ץN�e0��B�� ��ZN�lz%���;� �N�	[�rB_��Z�`�M�;���$�����#�8���&����N��b��s��E�^��J��FG��d����^^k�v�ʽ�!!�:k�1���Q�˾�������,���W'���*�j'�]%�M��D���7ʾ�"���h�����   �   LA%��׋��B7��Mټ	���P����@�۾[(���r�gܥ�ؿ�<��#�^FA�H�]���u�?��Z���`����u���\�J�@���#�4&��'ؿ;��is��(�q�ܾ�䅾���EQ��,��`�L��k����+���8m���<�`�y�wĚ��X��*Qʾ�׾�ܾ2׾eqɾ
4��j~�� hw���:��C��L���   �    @d:�v4< ,�;`l��Dݚ��u(��3���q���?�O������'����8��[�І~�'^��:����9��(w��9��R~�:�[��8����ز�B���։��@������g���i*��'���*�� �j;�< �!�$ҿ�3c������r	��42��V�.>s�����Oƅ�^f��m�q���T�MF0��s�έ����[�����   �   �r�<�<�~{<�w��f1��E�:��o��&f
���Q�ٷ���ʿ�N�z�$�
�I��.r��l��C����v/��H�������d��
ar�f<J��9%� ���˿5{��DS��X�H檾�=�欽�-�� 9d<���<���<Hk<,޻̑���|�m������
�	��I������Ȃ�� �蚴��v�0� ������<�   �   ̍6=z�%=��<Ȕ��7����F�/���t����]������ԿH�	�0C-�@AU�!������1V���;��=����6���^��N0��E�����U��.���
�ֿ����t_����Y���$HI��3����,�<>[ =X�0=h�=६<�<�:h����,�R"{��k��c����c�����������v��A'�t(��`�2;,=�<ZD=�   �   $'c=��L=4��< ���Ě�]6�x駾S�	��aQ�vh���9ʿ�
��c$��yI�$�q�%W�����P,��i���1��3?��饍���r�2�J�P�%��$��̿Wᖿ�S���W���|Y:��졽��L�@��<N�A=�/X=�C=�L=4ə< �9�u�� ��Z�A��b���l�.�_�pC<�H�����U+;0�<`9=��N=�   �   ��N=nM?=�?�< :�}r��I!2������7��M�Eޒ���ƿ�� ���!���E��&m�dX��/���
J���e���C��D���I���P�m���F���"�J���ȿ�?��<�O�6���!�� R6��p���N�0`�<�:4=.�C=�$(=�[�<�<��K��L�O��ׄ���������l��[災z�G�,���P�!��2<���<B;3=�   �   =V�=�R�<@7)�h'����&�&����8��ɰB��w��^Y��D���>����;�N�_�Q��>���G>��+������ei���ځ� `��J<�"���4��U������T�D�N������*�:��� /X��<B�
=�=�.�<�P:`�Ƽ��Q�˞���νW[��t� �	�� �R��I-ʽTk��HF�$��@�a;�+�<�   �    �<�z�<��T<�J��倽����������t�1��� A��������lQ,��K��j��ʂ��݋�X���s����m���Cj�^�K��X,��&��s㿦��J�����2�@��)����6�������u��*≮�<���;Xx�&�9�8]�����
� ���B��j]��Yn�B�s�49m��S[���?�K_����&�����,��1G��   �   �H�7 �`������ڌe��P��q�^�ɾE���a� ؚ��:ʿ�f��`b��?4���M�|>c�n�q��v�vq�Ab�L�L��~3���&���^ʿ!2��ڻb�!���h˾�pt�����qo�8_��c���+��������v齄�*��d������Φ��`���ƾ��ʾ�ƾ�������勾��_�,�&��ℽ�   �   Pf�� �6�|�Ǽ8μr�N�/I׽q.H�ŋ��(T���?�N���8��Kۿ"x�����|/�HU@��fK��O���J�\I?�jX.� ����� 4ڿ<ޭ������-@�6��^{��kJ��)۽
�V�x�޼8�ټ�2A�����R���=V���������w�^1�L�8��ݵ��]�`��G��|n���$����Q�~���   �   )��پ�L�^�X��jD�ⳮ�@��P�����Ӿ�}��=Z�児�����ǔݿvl�(��6���'��j*��'�BD�����m �kܿ����zߏ���Y�s>�W�ӾT憾���.$��^J��	%�,�f���ý�X �$s��|��=�㾇��Z+��lD�$X�`d��]h��c���V���B�y�)�@T������:o��   �   x�K����8.o��	L�������9zL�������� ,�&f�ړ��g���jWѿ�1��� ��/�VM	���������Z꿬�Ͽ�;���r����d� +�!��у��HL�kM�0����\O�8�s���½p� �b>{�����|���Ü$�fIL��jr���������Y-��Ρ�Y������|܈��p��&J���"�N����s���   �   9��S�k�2p��Э��i�h�i�G������aYm�����!5��.��a�'R���碿�j��'ɿ�ӿW�ֿ^�ҿ��ǿ�����o�����1_�QZ-�	 ����T~k�m��ͭ��i���i�����X��_m������7�y�.��!a��T���ꢿ�m���ɿ��ӿ��ֿ��ҿ9�ǿ����or��%��+	_��]-�� ��   �   *�򾤆���!L��Q����
[O�n�s���½�� ��7{����������$�EL��er��􉿛���6*���ʡ�B�������و��p��"J�C�"�ѹ��co��x����y��)o�(	L�����
�~L����!���,��f�3���+����Zѿ5�ƕ ��1�XO	�z��5���^꿧�Ͽ�>���t��4�d��+��   �   �@�W�ӾM膾(��-&���J��%�h�f��ýrS ��s��w��>����V+�IhD�X��Zd�NXh�ťc�ҸV�g�B�z�)��P�F�ྔ���p�n�$�2Ӿ��^��T��kD�Ӷ��!��������Ӿ?���@Z�臐�k�����ݿn���8��'�&m*�� '�@F����,o �ܿᤵ�L᏿��Y��   �   �/@����Y}���J��+۽V�V�x�޼P�ټ 'A���������6V�]���_��tq侸-�+H��3���Ʊ�Z������*i��� ����Q�6���^����6�luǼ(μh�N�uL׽|1H�,����U�1�?�䙄�:���ۿ�y����x~/��W@�`iK�@O���J�~K?�HZ.������N6ڿ ୿틄��   �   ��b�|���j˾st���fro��Z���6��H�*��r� |���k齲�*�bd��덾mɦ��Z���ƾ��ʾ�ƾ��������l�����_���&���3ڄ��1�x � ������t�e�>R��q���ɾ���X�a�wٚ��<ʿ�h���c��A4���M��@c��q���v��q�@Cb�,�L��3�V��(���`ʿc3���   �   �����2��������7������u�)*<lŃ<`��;X�w���9��S������{� �,�B��b]�uQn���s��0m�L[�u�?��X����3���j�,�8G���<$��<(�T<ȝJ��怽|���������1���@B��J������R,���K���j��˂�ߋ�� �������n���Ej���K��Y,�V'�3u㿨���   �   �����D���/����*������*X�8�<\�
=�=>�< �:p�Ƽp�Q�����νQ��J���	�x����z$ʽ�c��� F��﮼�tb;d9�<"=v�=�U�<�8)��(����&�1����:���B��x��OZ��o�������;�~�_������2?��������/j��aہ�`�TK<����k5������   �   $@����O�b���!��$R6�mp���~N�<c�<:=4=>�C=�((=�e�<��<�vK����O� ӄ����&����g���⁽:�G�����w!� �2<`��<f>3=��N=�N?=�@�<�<�gs�� "2�P���m8���M��ޒ�8�ƿF� ��!�`�E��'m��X�������J��uf��7D������������m��F���"�|��0�ȿ�   �   4ᖿ��S�֙���� Y:�b졽`�L�x��<��A=X0X=v�C=M=�ə< 9du��ښ�*�A��b���l�(�_��C<�h������R+;�/�<9=B�N=�&c="�L=$��<��6Ś��6��駾�	��aQ��h���9ʿ�
��c$�
zI�B�q�2W����V,��i���1��*?��ܥ��v�r��J�:�%��$��̿�   �   {?����O����� ���P6��n��xvN��e�<>4=��C=)(=�e�<��<�vK����O�ӄ�$���=���h���⁽\�G����� w!�@�2<���<�>3=H�N=|O?=C�<�4��q��� 2�e����7�̞M�ޒ�b�ƿ�� �d�!�z�E�T&m�X��Ȕ���I��se��:C��Ɵ��ٌ����m�*�F�*�"����T�ȿ�   �   @���0�D�z�h
��6�*�~���HX�$�<�
=��=@?�< �:,�Ƽp�Q�����ν�Q��`��	������$ʽ�c�� F��﮼`xb;`:�<�"=֣=LZ�<�))��%����&�q����7���B�Nw���X��i������:�;�R�_����w���f=��>�������h���ف��`��I<�b��S3��_����   �   L���.�2��龟����4�𵆽(�u��6*<�Ƀ<��;0�w�`�9��S�������� �<�B�c]��Qn���s�1m�-L[���?�Y����6���>�,��G���< ��<H�T<�J��‽Q������h��\�1����@��{����fP,���K�h�j��ɂ��܋�&���F���yl��Bj�֢K�\W,��%�Rr�`���   �   ��b�i��Of˾Jmt�2��nho��M������*�Fq��{��zk齦�*�bd��덾xɦ��Z�� �ƾ��ʾ�ƾ�������{�����_���&����ل�P/�H � w��퉼��e�{N�L�q�l�ɾ���8�a��֚�=9ʿ�d��*a�h>4� �M�L<c���q���v��q��>b�P�L��|3�����#��]ʿ�0���   �   Q+@�d���x���J��#۽��V���޼d�ټ>$A�����]��h6V�V���`��|q便-�4H�4���Ա�Z������5i��� ����Q����]��$�6��lǼ�μ��N�ND׽J+H������R���?��Z6��#�ڿ�v�V���z/�&S@��dK�^O�*�J�(G?�vV.�R��H���1ڿ?ܭ�񈄿�   �    <���Ӿ�ㆾ�������J���$���f���ýS ��s��w��8����V+�PhD�(X��Zd�\Xh�ӥc��V�r�B���)��P�L�ྕ���L�n��#��Ѿ���^��M�aD�����������_�Ӿ�{��:Z����³���ݿ�j�^��4���'��h*��'�8B����k ��ܿ8���yݏ�w�Y��   �   ���g���>L��E������PO���s���½� �C7{�㙷������$�EL��er��􉿡���=*���ʡ�I�������و��p��"J�I�"�ҹ��Uo���
x�����w���"o��K�&�B���uL�}��{���+��
f�����Ӹ��mTѿ5.�
� �.�ZK	����Ζ��JW꿐�Ͽ=9��dp���|d�+��   �   ���3xk�gh�Bƭ�N�h���i�B�������Xm�ԏ��5���.��a�(R���碿�j��-ɿ$�ӿ`�ֿg�ҿ��ǿ�����o�����8_�TZ-� �����}k�$l��ʭ��i�n�i���������Sm�<����2���.��a��O��墿{g���ɿ��ӿ��ֿ��ҿ��ǿ���l��F��� _��V-�T ��   �   �x�Ί��q���o� �K�����I�nyL�H����� ,�%f�ړ��i���mWѿ�1�� ��/�\M	���������Z꿲�Ͽ�;���r����d�+��򾢃���L��J�4���zPO���s�`�½�� �)1{����������$��@L��`r�򉿭���#'���ǡ�*������׈��p�DJ���"�����j���   �   T�fʾ� �^��H�X`D����-�� ���S�Ӿ�}��=Z�慐�����Ȕݿxl�*��6���'��j*��'�FD�����m �pܿ����}ߏ���Y�m>�6�Ӿ憾���� �� J�T�$���f���ýN �� s�Rs���y�|���R+��cD�8�W��Ud�Sh���c��V�ԿB�`�)�JM�[z�����n��   �   �U��b�6� ^Ǽ��ͼ*�N�{F׽�-H�����T���?�M���8��Kۿ$x�����|/�JU@��fK��O���J�^I?�nX.������$4ڿ?ޭ������-@�,��){���J�'۽��V���޼|�ټ�A������s/V��
��3k�2*�SD��/������#V�F����ᾬc�����7�Q�`���   �   8�@���`��艼��e��O�y�q�2�ɾ<���a��ך��:ʿ�f��`b��?4���M�~>c�p�q��v�zq�Ab�N�L��~3���&���^ʿ%2��ڻb����h˾Lpt����*ko� L��`�����*��e��s��,a�'�*���c�.獾=Ħ�+U����ƾw�ʾ��ž>��������ۋ���_���&����rф��   �    �<h��<p�T< �J�L〽:������ؓ�n�1��� A��������nQ,��K��j��ʂ��݋�Y���t����m���Cj�`�K��X,��&��s㿨��J�����2�(������I6�_��� �u�0A*<ԃ<�<�;`�w��9��J�����.� ��B�F[]�QIn���s��(m�FD[�G�?��R����ۅ���,�p�F��   �   �(=��=8_�<�%)��%��:�&�����8��ŰB��w��^Y��D���>����;�P�_�R��>���F>��,������ei���ځ�`��J<�$���4��W������R�D�H�y����*�ɭ��XX���<�
=��=�L�<�:�Ƽ
�Q����̮ν�G��N����	�s���ʽ�[����E�Lخ��c;pI�<�   �   <�N=�Q?=�E�<�1��q��!2������7��M�Dޒ���ƿ�� ���!���E��&m�eX��/���
J���e���C��D���J���P�m���F���"�J���ȿ�?��<�O�3��!���Q6��o��XyN�`f�<:?4=��C=@,(=Hn�<��<�]K����X�O��΄�\���X���1c��<ށ���G����\!�P�2<$��<lB3=�   �   F��=
o=$$=`�y;^�g���b&��Ų�f�:��*��{��A�~b�Ш4�D�V�حx�X ��E��~����J��1?��|Hy���W�j�5����?k�I����އ���=���M������b�|���{��5=�j\=R�p=4^=$�/=���<X4.<p�Ȼ�㫼ZE�V�"�..+��2�D���X�����-�Ȳn<�=6B=�tp=�   �   ~�p=r�b=�k=�o;�a�Ƃ�������r`7��ۃ��|��>�����1�R�R�"�s��.��&���5w������9��%t�>�S���2��&�n�Ch���t��/�9��#�6����M��Wv�@�����
=bP=�n^=��D=(�=tm�< (`�h���
o��F�X3g�r�p�ڥb�x>�|o�T`���O;���<h "=�]W=�   �   ��7=r<=8�= �>;�Q�5o�rC���A�3|-�?Az�P���?޿��d�(�ȳG���e����7���ڋ�F����u���e��G��w)�0�� �߿BD����|���/�����T�����fd���̺,�<��)=Ԑ%=H��<8�3<H@�l���v��ئ���Ƚ�޽Bx��۽&Ľ|G����f�����h�~<6�
=�   �   �z�<X��<(&�< v:�r9�rG��)Rq�H�˾��5e�5���K�̿2b ��}���6��Q��Wg�r[v�x�{���u�6�f��xP��6� ��*� ���Ϳ?���K�f�߫�?�ξ�nv��� �зJ�@iP��<`��<�څ< �]�����n����ɽ��T&��u>���M�0RR��L�ʨ;�=�"���U뿽��p���ּ�ǧ:�   �   �s���;�$<��X��k ��>ӽNqO����/Y
��J�.J�������e忢�
���"�@�8��J���V�\�Z�4.V��I�L{7�t�!��Q
� �g׶������
K�6i��&���US�Z�ڽ�/���0p�;�ց:lp�S�t������*�D��Sw�r!���ã�ாM`���ﭾ����ɏ���q��$?��U��ⴽ�@��   �   �}��<���'� �5����K��n7*��"��d辽<+��n����ƿ���t2��d�~	-��6�~�9��5���+�1��&��x�P;ſд��5�m���+�b龘V����,��α��7�Huh��`���������J8���������ʾ��꾙�o
�2���j	��� ���羆�ƾ��$fy��o2�޾��   �   �������������ׇ�����i�
���B��JC����@���c�ȿP���>�B��|����2������jX���ƿv���;��I�B���
�ߢ����i��J��V��0_���ռ'�	ߜ��5�{OR��s���;ɾ�I�����:�/��bA�4�L��P���K���?���-�a�����qž�2��v�L��   �   �SU��Y��Ԗ�xJ+����D%S�k�Ľ2�.�0x����׾�M��,N�x냿b_��!h���տ�������՝��b��sC�v�ӿ�i��Y���Z����XL� �S־<��+.��#ŽV�����B2�����8��v�Y�%\��n�߾l��w�6�H�Y�x�I񇿻`������Ў�X톿��u���V��A4�"���Vܾ?����   �   ^����FJ�׃�i����&��(��������z�L�w����l	���I��x��䒿�����ҵ��V��[T¿���#|��5�K5����u��EG��&��V����mBJ�
~�f��b�&��(����b�����L��z���従���I���x�{璿�����յ��Y���W¿H���1����7��?�u�rIG��)�P[��   �   �V־�č�
/.��'Ž�V����<2������[�Y�X���߾��x�6���Y��x���]��4����͎��ꆿ��u���V�>4����Qܾs���LNU��U��ϖ��E+�F���)S�	�Ľ�.�{���׾�P�0N��탿�a��k��9�տk�迒���u�������F翆�ӿGl������T���\L��"��   �   ��
�������i��L�cX���^���ռ2'�؜�1��HR�Wo��6ɾC�������/�j^A�m�L��P�صK�r�?���-�²�����lž�.��G�L�.��֒���T|������ه�����i�+���r�rMC�����z����ȿR�꿤@��v~������f���>[�\�ƿ�����<���B��   �   j�+��d�aX����,��б� 8��hh�p`����}��b	��C8�T���{��ʾ�����
�h���f	�"� �@���ƾH��:^y��i2�D�罴v��x꼠�'�h�5�ą��N��*:*��$��3g��>+��n�{���!ƿ@���3��f�h-��6���9�
�5�z�+��2�R(�G{�R=ſo�����m��   �   WK�sj�^(���WS�b�ڽ�/�P�P��;�ۂ:@ם���S�tz�������D��Jw����c����ڮ��Z��ꭾ]����ď�S�q��?��O�Uٴ�x@���r���;��$<��X�n ��Aӽ�sO�����Z
��J��K�������g���
��"��8��J���V���Z�>0V�ʼI��|7�̹!��R
�� ��ض������   �   ��f�߬���ξzpv��� ���J��SP��<��<�< �\�����#f��J�ɽ�~�pM&�vn>��M��JR�$L���;��|"�
 ��´x�p��}ּ@	�:���<���<+�< v:u9�<J���Tq��˾���e�X�����̿c ��,�6�0Q��Yg�f]v�t�{�|�u��f�NzP�D�6���� ��Ϳ-����   �   {�|�?�/����xU�����tgd���̺��<��)=4�%=x��<0�3<p�?�nt��v�|Ц���ȽK�ݽ�n��y۽gĽ�?����f����PO���~<��
=b8=P<=��=`�>;�Q�Xp�aD��YC�3}-��Bz�+ª�@޿��0�(�ȴG���e�>�������ڋ����w�дe���G�Bx)������߿�D���   �   �t��q�9��#�c��� N��Wv� ����
=tP=Pq^=�D=��=@x�<��^�䃞��f�t�F�h*g�l�p��b�&>��g��R���oO;���<:"=�`W=��p=��b=Hl= o;��a�������p��a7�܃�K}���>�X���1���R�ؽs�/�������w��?���Z9���%t���S�F�2�'�qn뿅h���   �   oއ�h�=����������t�|���{�
6=2k\=��p=�^=��/=d��<�5.<@�Ȼ\㫼,E�0�"�.+��2�d���������-�бn<��=�B=�tp=��=�o=�$=��y;F�g� ��&�����:�+��:{��h�b��4�Z�V��x�a ���E������J��)?��fHy���W�T�5�l��k�%����   �   Jt����9��"󾉀���L��Tv��b��R�
=>P=�q^=h�D=��=�x�<��^�����g���F��*g���p�.�b�J>�h�S�� oO;���<V"=�`W=��p=d�b=vm=@2o;��a�t�����7��4`7�oۃ��|���=鿾�8�1���R���s�F.�������v��i����8��T$t���S�x�2�t&�qm뿻g���   �   *�|���/�W���S������ad� :̺��<�)=(�%=���<`�3<��?�\t��v��Ц��Ƚs�ݽ�n��y۽�Ľ�?����f����0O���~<�
=08=�<=ę=�?;�Q�Dn��B��Aᾊ{-�Y@z�����F>޿p���(���G���e����}���Gً�����Ht�z�e��G��v)������߿aC���   �   }�f����H�ξlv��� ���J� P���<,��<��< �\�����f��B�ɽ�~�{M&��n>�&�M��JR�@L�ԡ;��|"� ��´|�p�$}ּ �:���<���<(1�< Kw:�m9�zD��.Pq���˾���e�O���'�̿|a �}���6�>Q�NVg��Yv�~~{���u�l�f�NwP�̙6���H� �m�Ϳ��   �   �K��g�s$��DRS�[�ڽl/���`��; )�:,ԝ���S�/z�������D�Kw����o����ڮ��Z���ꭾo����ď�p�q��?��O�Aٴ��@�(�r�P+�;�$<�sX�,e ��:ӽ�nO�����W
��J�I������+d忎�
�F�"���8�F�J���V�>�Z� ,V��I��y7��!�`P
��忶ն�?����   �   D�+��^�-T���,�ɱ�.��Nh���_��*}����C8�B���{��ʾ�����
�s��	g	�.� �T���ƾR��D^y��i2����v���s��'���5�|�fG���4*�� ��Aa��:+�2n����ƿM��1�(c��-��6�l�9���5���+�R/�j%�Kv� 9ſ����J�m��   �   ��
�����!�i�@G��P���T�X}ռ�'��֜��0��HR�Fo��6ɾ C������/�r^A�x�L��P��K���?���-�˲�����lž�.��&�L����������o����"҇������h�2���P��GC�\���8�����ȿ}��Z=�~��z���J����>�pU�R�ƿ>���=9��^~B��   �   �N־"���'.��Ž>
V�6��F62����N����Y��W���߾��w�6���Y�x���]��<����͎��ꆿ��u���V�%>4����Qܾg���NU�pU�Ζ��?+�޴�(S�K�Ľ-�.�ru��@�׾IK�d)N�}郿]��de����տ���w���?������@�R�ӿ�f��ڨ��:���TUL�Y��   �   ^����<J��u��_����&��(���ړ���L��v����g	���I��x��䒿�����ҵ��V��cT¿���,|��<�S5����u��EG��&��V������AJ�f|��c����&�x(�
��&���p�L��s��h�~��I���x�MⒿ됦��ϵ�mS��Q¿ג��y��Tꤿ�2��Z�u��AG��#��Q��   �   �GU�#Q�qȖ�t9+����S��Ľn�.��w��߶׾�M��,N�x냿c_��"h��	�տ������ߝ��j��zC��ӿ�i��]���]����XL� �S־�+.��!Ž�V�"���12�[����}�x�Y�T���߾����6�A�Y�
x��뇿[��W����ʎ��熿��u��V�/:4���_LܾI����   �   ���͊��0��|f��^���Ӈ����i�ޚ��7��JC����?���d�ȿS���>�F��|���6������pX���ƿx���;��J�B���
�����m�i��I�wS���U�0wռ��&��М�),�bBR�5k���0ɾ�<��4���/��YA���L��P�%�K���?�Z�-�
��u��Pgž7*����L��   �   ln��^��'���5�B|�`I���6*��"���c辶<+��n����ƿ���t2��d��	-��6���9��5���+�
1��&��x�T;ſҴ��7�m��+��a�dV����,�5̱�0�`Gh���_���.v��B��V=8�L��w��kʾ�|꾇��
����Oc	��� ��}��ƾS���Uy��b2�����   �   �r��k�;�$<@QX��e ��<ӽ�pO�f��#Y
��J�-J�������e忤�
���"�B�8��J���V�`�Z�6.V��I�P{7�v�!��Q
��i׶������
K�0i��&��US���ڽ�/���p��;��:L�����S��p�������D��Bw����B���2ծ�9U��孾6��������q��?��I�[ϴ���?��   �   ���<��< 8�< �w:Tn9�F���Qq�+�˾��1e�5���K�̿2b ��}���6��Q��Wg�v[v�x�{���u�8�f��xP��6� ��+� ���ͿA���M�f�ݫ�)�ξvnv�� ���J��P�H$�<���<L��< $\������]��c�ɽ>y� G&�tg>���M�CR��L���;�Fv"�6��r׿�|�p�haּ@w�:�   �   n8=d<=�=�)?;Q��n�SC���A�.|-�>Az�P���?޿��d�(�ȳG���e����8���ڋ�G����u���e��G��w)�0���߿DD����|���/�����T�����:dd��G̺ �< �)=��%=��<(4<�?�$h�֎v��Ȧ�V�Ƚ;�ݽ�e佪p۽��ýi7���f�
��`���<��
=�   �   ��p=Z�b=�n= >o;��a����������q`7��ۃ��|��>�����1�R�R�$�s��.��$���4w������9��%t�<�S���2��&�n�Dh���t��1�9��#�(����M��Vv��w����
=`P=�s^=P�D=��=���<�]�|v���_�T�F��!g���p�f�b��>�(`��D��`�O;$Ķ<�"=ndW=�   �   �w�=�K�=~�U=�~�<�
����=�p�|�;	��2�g����;$ϿN���5�09��T�3k���z��M���{�dk��T��:��F����8bѿ�à�|4k� �"�W�Ҿ�!y�����<(���M<lw7=�%z=�/�=��{=t�R=4v=�*�<�E<=��h�q���������Ў���B�����\<L��<��6=n�o=��=�   �   5�=���=܄O=���<r���h3k���ɾ_��ɮc�X��T�˿x^����\6�h;P�|�f�`�u�K{���u�`�f�b�P��6�|��� ���Ϳ,���d�f�f��q>ξP�s�����&y"�P�L<��1=�3o=��{=�;e=�+6=���<@�Q<@Db�DǑ����H�0t�����CԼ�]^����:\��<D�=�^S=��=�   �    2g=Z�j=*�<=�՚<��B,ս�[�J����'�e�W�.^���¿�h�Q���,�R8E�D�Y�΅g��Wl��Mg�6oY��$E�5-�(��(�����ÿ�ו��Z�x�������cc�.E��O���F<�% =̍M=؏I=,� =`3�<`�H;������!��n�ǒ���Ʀ��櫽-m���$��<�[�.�� 3I�8h!<��<Ȟ>=�   �   j�=t^.=n�=�<�<�ż�����=D����c��H2E��-���ǲ�M�࿊��h&���4��zF�TR�
[V�n�Q���E�Z4����D��)ῌ��� ���G��k�ac����J���ƽ�T���0<T, =$�=Ԛ�< }*<��e�i/�T=�� ӽ�d�T\��h&�5D*���$����)���ǽ҈�����Ỹ��<�   �   �J;`��<Ŀ�<H`U<����C�����&�����J��De-��q�
��c�ȿ���P���} ��/��F9��<�X�8�֢.�.���<��
�>ȿ�0���q�u.��:�����+�ۂ���zļ@h�;X�<�m< h���⃍���{a�>�K��r��jD��2��,��z����m���D���Y�ԽVe}��ϼ�   �   �(%����`��;P��;8�r�Vnq��e��.s�;ľGd��:M�[���ˬ���ѿc���n
�F��N���^!�A�����[	�Q{��}п�������M�H��Wž�
v���	�0���Κ��%�: -�:p1v�8�>�����6q��"S�	i���S��ݫƾ�ܾ����#�v龼Yھ�Hþ�l���P���K��������   �   �mƽ8-H��咼@䳻H�X��A2���˽��=� N����쾕�'�g�`�._������Ϳ����2}���Z��;���X�-˿�S���,��I2_���&�h��;V���>��_Ͻ�;��l����9���]\�@ҽ5+�rz�.����ؾ���yx��&��/���2���.��u$��_�C0 �YUӾ�7����r�n2$��   �   ��+��ɽ��K� ��
y�����&�����
�˥k������5L1�S8d�_7��n��ߺ�:�˿:ֿǁٿ�SտS!ʿ��-��������a�c/����J_����i�Q
�q�����hN��|�Ƽ��X�zJҽ�11����Ak��+T��B��Wf;��YV��Rk�px���|�Qw�GGi��S��8����u��fR���U���   �   $ǁ��"�V��Rt2��ɮ�\α��7��g��X�%�����N����G�>w-���V���~�g֐�\��(ʦ�l��������X6��Id{��S���*�`:�ж��Dā��"��P���n2��Ʈ�tӱ��7��m��Ϋ%� �������J��z-��V�<�~�ِ��^��ͦ�
o��}������8���h{���S�	�*��<������   �   �b��R�i��S
�������K����Ƽ��X��Bҽ�,1�{����f��PN�����Fb;�LUV��Mk��jx���|�Lw��Bi���S��8���p��N��rR����+�\�ɽ&�K�|����y�<���+���B�
�֪k�@���X��JO1�<d��9�����ếF�˿C=ֿ��ٿ�VտH$ʿ��;0����x�a��e/����   �   ��뾞X��(�>��cϽV�;�l��H��p)���Q\�k7ҽX+�ojz�m����ؾ����t��	&���/�Z�2���.��q$��[�- ��OӾ3���r�-$��eƽB"H�ؒ�`̳���X�>F2�r�˽4�=��P������'���`�)a��Z��MͿ���6���~�������>���[忭˿V���.��;5_�"�&��   �   ���yYžv���	�U2��`Ϛ��~�:@��:Pv���>�״��Qk�<S��d���N���ƾ��ܾI��)ﾎo龚Sھ2Cþ�g���L���
K�������l%����`��;���;��r��sq�%h�z2s��=ľ2f�G=M��\���ͬ���ѿ�e��(p
������f`!��B����]	��}��п��N����M��   �   �v.��<�^��ҩ+�����P|ļ�v�;0�< +m<�ng�&�{��5���Z��}K���r�R����?��"-��T'��������l�b�D�{��Խ�T}�x�μ��J;���<���<�cU<����邚�!�&�y������g-�Gq����,�ȿ�����d ���/�:H9�6�<� �8�Z�.�����=���;@ȿ2��$�q��   �   �G��l��d���J��ƽ�V����0<j/ =J�=���<ȣ*< �e��Y/�A4����ҽ�^��U�Xb&�|=*�e�$����������ƽ|Ɉ�����w����<��=�b.=��=8=�<�ż�����?D�_������3E��.��4ɲ�С�p��z'��4��{F��UR��\V���Q���E��4������m*Ί���� ���   �   ��Z�������|dc�&F�RP���F<�' =.�M=��I=z� =<C�< LI;������!�	n�犔������ޫ�e��C���[�����I���!<H��<v�>=6g=��j=b�<=�՚<���3.ս��[������(���W��^���¿�i�hR�v�,�H9E�^�Y� �g��Xl�Og�<pY��%E��5-�������P�ÿ�ؕ��   �   ��f�����>ξ��s�����y"��L<��1=d5o=>�{=�>e=�/6=X��< �Q<��a� ���@��X�4l�.��05Լ�B^����:�ɚ<��=VbS=a��=& �=|��=6�O=���<��d��t4k�u�ɾ�����c������˿"_��X���6��;P��f��u��K{�.�u��f�ԐP�F�6��6� ��Ϳg����   �   F4k�ԯ"��Ҿ~!y�[���;(� �M<�w7=&z=�/�=�{=��R=zv=$+�<�F<P;����q�L�����������(B� ��\<���<��6=:�o=��=�w�=�K�=�U=�}�<h
���콣�p���;5��h�g�%���\$Ͽb���5� 09��T�3k��z��M���{� dk��T��:��F����bѿ�à��   �   ��f�Ԑ��=ξ!�s�����bv"���L<��1= 6o=��{=D?e=�/6=���<X�Q<@�a�$���h��r�Pl�H��d5Լ�B^����:�ɚ<��=vbS=}��=V �=ө�=@�O=� �<h�u�� 3k�b�ɾ'��x�c� ��
�˿^�����
6��:P���f���u�tJ{���u���f�ЏP�p�6����� �$�Ϳ�����   �   �Z���������ac�]B�HK� �F<* =��M=��I=� =,D�<�PI;$�����!�$	n����������ޫ�"e��d��B�[�̗�PI�p�!<���<ؤ>=�6g=$�j=T�<=�ۚ<dz�*ս��[�|���9'���W��]��L¿�g�0Q���,�|7E�F�Y���g�zVl��Lg�nY��#E�.4-�v��������ÿ2ו��   �   	G��j��a���J���ƽ�H���0<�2 =F�=(��<`�*<��e�tY/�)4����ҽ�^�V�ib&��=*�{�$���������ƽ�Ɉ����@vỴ��<��=zd.=d�=�E�<��ļ៺�<D��
�����1E�(-���Ʋ������x%���4�2yF��RR��YV���Q�$�E�4����Z���'�C������   �   8s.��7����$�+�e~���kļ@��;d�<�4m< Ug���z�����Z��}K���r�\����?��1-��d'�������l�z�D����Խ�T}���μ`�J;ܞ�<`��<(xU<�����|����&�������c-��q�����ȿ���2���| ��~/��D9��}<���8�H�.�ĕ�H;�q��<ȿ6/����q��   �   N��,Tž�v�t�	��+��8��� @�:@k�:v���>�M���$k�S��d���N���ƾ��ܾY��=ﾠo龮SھCCþ�g���L���
K����Ь��H%�(�����;`��;`�r�Bfq�2c�3+s��8ľ�b��8M��Y��7ʬ���ѿ�`��Jm
��������\!�\?�\��*Z	��x�{п�﫿?���M��   �   |��TS����>�YYϽ��;��Y�����l!��O\��6ҽ+�Hjz�_����ؾ����t��	&���/�e�2���.��q$�\�- ��OӾ 3���r��,$�heƽ, H��В�������X��82�s�˽��=��K��?��L�'�{�`�`]������&Ϳ�|�����{�H������7��V忌˿�Q���*��	/_�E�&��   �   �[��]�i��L
�#������9���Ƽ��X��Aҽ>,1�[���~f��DN�����Ib;�QUV�Nk�kx���|�Lw��Bi���S��8���)p��N��gR��~�+�e�ɽ��K�������x���������O�
��k�c����bI1��4d�D5����]ܺ�H�˿�6ֿ�~ٿ�PտVʿL�J+��s���4�a��_/�N���   �   �����"�fI���b2�����0����7� f��Ц%�����5����G�:w-���V���~�k֐�\��-ʦ�"l�������_6��Ud{��S���*�c:�ȶ��*ā���"�gO���i2�T���𻱼Z7�a���%�����Q���NE�t-��V��~��Ӑ�SY��OǦ�6i�����;���3���_{���S�v�*��7������   �   &�+���ɽ��K�t鲼��x�����ԗ��&�
�T�k������0L1�O8d�^7��p��ߺ�?�˿:ֿ΁ٿ�Sտ\!ʿ��-��������a�c/����7_��|�i�bP
�X������9���Ƽ��X�;ҽn'1����$b���H��d��b^;��PV�:Ik��ex�s�|�	Gw��=i��S�
�8�:�\j��aI���N���   �   �\ƽ�H�����}����X��;2���˽��=��M����쾍�'�d�`�-_������Ϳ��	��4}����^��;���X�0˿�S���,��L2_���&�]��V����>�^Ͻz�;��[�� ��l��LD\��.ҽ�	+�.cz�囩�dؾi��%q��&���/�%�2���.��m$�UX��) �QJӾn.��]xr�'$��   �   �%���P��;���;��r��iq�e�@.s��:ľ>d��:M�[���ˬ���ѿc���n
�F��P���^!�A�����[	�U{��}п�������M�E��Wžz
v��	�>.������ q�:��:��u���>�⫹��e�'S�X`���I��v�ƾ��ܾ��꾝�i�uMھ�=þ�b��GH���K���������   �   `QK;<��<H��<�U<䁚�}~��A�&�����3��<e-��q�
��b�ȿ���P���} ��/��F9��<�\�8�آ.�0���<��
�>ȿ�0���q�u.��:������+�)���pļ ��;�< Mm<��f�� ��r����㽦T�WvK�V�r�֡���:��T(���"��v���r�l���D��K�Խ>C}�0�μ�   �   4�=�i.=��=LH�<��ļQ���}=D����[��D2E��-���ǲ�N�࿊��h&���4��zF�TR�[V�n�Q���E�\4����F��)῎��� ���G��k�Mc��E�J�Q�ƽHM����0<�4 =r�=���<��*<�te�K/�|+���ҽJY��O��[&��6*��~$�q��d�����ƽ������������<�   �   �;g=��j=r�<=Xݚ<,{�v+ս��[�:����'�a�W�-^���¿�h�Q���,�T8E�F�Y�Ѕg��Wl��Mg�6oY��$E�5-�*��(�����ÿ�ו��Z�w������Tcc�qD�fM�`�F<+ =
�M=��I=�� =xR�< �I;������!��m�H�������q֫�]�������[�Њ���H���!<0��<�>=�   �   �!�=���=f�O=D�<N����K3k���ɾ]��Ȯc�X��T�˿z^�����\6�h;P�~�f�b�u�K{���u�`�f�b�P��6�~��� ���Ϳ,���e�f�e��m>ξ9�s�P����w"���L<:�1=(7o=��{=�Ae=N36=��<H�Q<@~a�ث�������~d�����&ԼX'^��Q�:�Ԛ<D�=VfS=	��=�   �   ă�=�~�=B�=,�=�&����r�8�������J�?�VЄ������}ۿ�������0�46B�N�M�:"R��M��XB�n
1�v9����}[ݿu������9C�������GC����`���`U�<�P[=��=ґ=�=��r=�ID=�=d��<��K<�l�;�Z��&��@k�:��<��<��<�?8=�p=I��=l�=�   �   �0�=���=c��=��=����s��24�+��� ��}<�����N�����׿T����X�-�P�>�t1J�F4N��(J���>���-�x��8s��ٿm���2��V�?�0��"u���~>��V��t^���r�<��V=3{�=7Պ=�"�=:XZ=�5&=�}�<`�V<���: S ��aX�H�j�8�4��h�p��;�:�<�\=f`R=��=	%�=�   �   �Ս=B�=�+v=��=����EӍ�>\'�V*����c2���w�{R��*�Ϳ�4�����%�d�4��r?�@C��I?��4�x%�:�����m�ο����%mz���4��q��nۛ��0����H�r�xB�<�4H=��n=��j=��G=.{=���< ��Q��&���8��9V��L]��$M�J'� �ܼ�v�p<ؽ�<t>=�ix=�   �   ��N=ڇi=H X=b�=�}Y��Oo��������ھ��"�H�b����Ƞ��4��Np�T���&��N/��i2�6/���%����6����=��ZӖ���d��d$���޾@j��z�N���'��=�<0�-=\"==N� =d`�<`1\;������?������-��D��N
��Ռ�F�ٽ@ಽ��fv���/�0�j<>%=�   �   h��<(2=x�)=��<@�Z;�9�P���v�g��Ͻ��\��H�#��Uڨ��BͿE𿸈����֩��=�JB�:$�^������̿ ����=����H��h�>K��ւm�_��>U��Z��(Y�<�=Ȏ�<��M<�wE�h2�H@��b����@d=��V�M�f��yk�`Rd�R�y6�����۽,{��H#�@�κ�   �   p�q�pm?<�R�<ȃ�<���;�@��L���<��@��*ﾭ�)��Ac�]���gﰿ�gϿ�.꿣��,��I�b��J����v���ͿO����9���b�Ui)�;���v���?��ǽ����:�d�<�9�<�R;�ü$?|���ܽPJ#���Z��+������0����=��D����̼��ۯ��0��z�����P�`���Ƚ�T��   �   [ف�g���|;��j<q�;@R��ඈ�l<�BOw�ގ����	�8:� Wo�bߒ�yϬ��ÿ�տ�$�a�㿾I߿��ӿ�������i��X+m�u�8����h۾��\w�zz��Q���峼 �S;��<`���<����$�UD�F���9ʮ�E�Ծ�i��^�X���&����m�����Ͼ����9{���:�6G��   �   #���Ʌ�x7ü �Ƹ���;�s�N,�o�Ƚ�6�[�����Ծ����D=�D�i��^�����������>����~G���o��.�����f�:�:�[��kAҾ�Ə��x4��#ǽa-�@��@�C; �g�������:��5�S�?����˾С �2���v1��TC���N�;�Q��xM�-hA�`�.�0������apƾq���4�K��   �   a�I�K��[l�<�� �y���I��K���]w��1��0�N�0Û��Lپ���2���S��q�����Ћ����.��+h����n���P�/�����ԾdO����I�=D��Rl�@2�� �x� J�W���gw�+9���O��ƛ��Qپ���%2��T���q�����ҋ�f���0���j����n���P�R/�S�%�Ծ�R���   �   �ɏ��|4��(ǽ�f-�(���D; �g�T�缄����� �S�;����˾֞ �����r1�`PC�D~N���Q��tM�dA���.���Y����kƾ������K�����Å��(ü ���`�;��$,��Ƚ,�6�^�����ԾE��H=��i��`��i������ز��������
J��r��E���B�f�<�:�� �EҾ�   �   K޾�aw�-}�6U���볼@�S;�< ��(����  ��ND�D���cŮ���Ծ�c���Z�Ø�#�:�������Ͼ���rw���:��=�ҁ� T��`a|;��j<�m�;�Y�������?��Sw�����	��::��Zo�cᒿ�Ѭ���ÿ!տ�'�=�㿈L߿M�ӿt������`k��z.m���8�����   �   ���x����?�b�ǽV�� u:Di�<D�<`%S;�ü�/|���ܽD#�,�Z�Z'������ᔲ�n8������LǼ��֯��+��L�����P�t��UȽ��T�x�q��?<l[�<��<���;�D��P���<�SC��m�׊)�`Dc�
���^�+jϿ;1�W!��v-�ZK�ƻ�����x���Ϳ$¯�1;����b�@k)��   �   Ij�M��O�m��	�(BU��`��\�<��=Ԛ�<�N<IE�`�1�7��M��v��]=�A�V�!�f�Xqk�LJd�[R�r6�����۽Zr��&��Nͺ���<�7=��)=���<@gZ;J�9�1���~�g�ҽ�J^��H�i���ۨ��DͿW!���B��0��?��C�t%�x��� ￊ�̿b����>��h�H��   �   �e$�6�޾Ak��J{�����*�x?�<��-=�&==�� =�p�<��\;h���t�?�0������g���8��������󽴬ٽ�ֲ�|v���g�x�/�8�j<-=D�N=��i=RX=��= �Y��So����皇���ھ�"���b����������0q�T��&��O/��j2�^/���%�
���7�<��^��BԖ��d��   �   ��4��r��ܛ��0�n�� �r��C�<L6H=v�n=��j=DH=�=(	�< Lظ8;����f�8��+V��>]��M�'�܎ܼ(K��3<���<�$>=�nx=O׍=4C�=�,v=ڏ=����ԍ��]'�_+����d2���w�IS��!�Ϳ�5��t���%�:�4��s?�*C��J?���4�$%�������4�ο:���nz��   �   ��?�`��`u���~>��V��t^���s�<��V=�{�=E֊=-$�=�[Z=�9&=ć�<�W<�[�:�8 � FX�Șj�(v4�@�g����;�D�<a=*dR=C�=0&�=�1�=>��=���=Z�=����u���24��+��� �D~<� ���Ʋ����׿�����Ʊ-���>��1J��4N�n)J�2�>��-����rs�F�ٿOm���2���   �   ~9C�Ώ�Q��qGC�r������\V�<hQ[=��=:ґ=��=�r=�ID=n�=���<ЏK<�m�; O��"�� m�:��<h�<��<j?8=ʾp=.��=Y�=���=�~�=�A�=��=@)�����Ǥ8�7���Ι�v�?�pЄ�ΐ���}ۿ �������0�@6B�T�M�:"R��M��XB�b
1�h9���_[ݿ�t��󙆿�   �   ��?����pt���}>�<U���Y���v�<ԸV=Y|�=�֊=^$�=�[Z=:&=��<�W<�\�:�8 �`FX��j��v4� �g� ��;�D�<a=:dR=J�=K&�=�1�=���=��=��=@���\s���14��*��T �a}<����������׿��B��-���>� 1J��3N�x(J�R�>�F�-����r�W�ٿ�l��F2���   �   ��4�p��Mڛ�u�0�!��0�r��I�<`8H=�n=��j= H=��=�	�< �׸�:����v�8��+V��>]��M�B'�,�ܼ�K��3<���<�$>=�nx=�׍=�C�=�.v=��=�ꞻ�э�B['��)�����b2���w��Q��n�Ϳ�3��@��n%���4� r?�\C��H?�*�4��%����� ��m�οĜ���kz��   �   �c$���޾�h���w�~��@��G�<��-=�(==�� = s�<��\;l����?��������i���8�����́�Ԭٽ�ֲ��v���g�P�/��j<�-=:�N=*�i=�X=L= {X��Jo�8������Z�ھ��"���b����������忈o�l���&��M/�\h2�
 /�j�%���6�Q�����?Җ�d��   �   gg��H��pm���67U�@%��Pf�<�=���<xN<(DE���1��6����h��]=�F�V�4�f�nqk�bJd�wR�0r6����۽`r����@Aͺ���<l9=~�)=���< �Z;̝9�d�����g�ν�y[�1H����ب�TAͿb𿤇�������f<��@��"�4������̿o����<����H��   �   ޚ�Lt��O}?���ǽb���}	:dt�<�K�< OS;T�üh.|��ܽ�C#��Z�U'������锲�w8������[Ǽ��֯��+��W�����P�{��?Ƚ�T�8�q���?<�a�<��<�0�;b9�sH���<��>��Q�Ȇ)�4?c��������eϿc,����*��H��������t近�ͿW����7��I�b� g)��   �   ؾ�Xw��v�bL��\ӳ��0T;h�<�B��"������zND�0���XŮ���Ծ�c���Z�˘� #�C������)�Ͼ���uw��ބ:��=�ҁ�pP�� �|;H�j<@��;�B�����F9��Jw�򋿾Ț	��5:�To��ݒ�Tͬ��ÿ'տ�!࿋���F߿��ӿ����B���g���'m���8�����   �   �Ï�:t4��ǽV-���� �D;�9g����E��M����S�;����˾Ҟ �����r1�gPC�L~N���Q��tM�(dA���.���d����kƾ����p�K�6�����"ü \���=�;(S��,�7�Ƚć6�������Ծ?���A=���i��\���������t�������"쳿�D��Wm�������f��:����P=Ҿ�   �   �I��;��El�H�� Po� �G��A��nZw��0����N�Û��Lپ���2���S�!�q�����Ћ����!.��1h����n���P�/�����Ծ]O��L�I�wC�DPl��)�� �q� rG��8��Rw��)���N�˿���HپY��]�1���S���q�Q����͋�a���+���e��8�n���P���.���(�Ծ�K���   �    ��S���Lü ���`J�;8Z�,��Ƚu�6�5���r�Ծ����D=�B�i��^��������%���E�����G���o��2�����f�@�:�[��eAҾ�Ə��x4��"ǽZ]-�h��`�D;`g� �缰��<��B�S�Y7���˾�� �l��(o1�RLC� zN�|�Q�_pM�`A���.����{����fƾˌ��T�K��   �   �ʁ�<;���};0k<���;|G������;��Nw�������	�8:�Wo�aߒ�{Ϭ��ÿ�տ�$�g���I߿��ӿ�������i��\+m�w�8����[۾��\w�z�lP���۳� "T;P�<`����;��$��HD�j�������9�Ծ�]��YW�A�����������	򾘵ϾF���{s��x~:��3��   �   �Rq���?<Tl�<��< 1�;2<�K��<��@��ﾦ�)��Ac�\���fﰿ�gϿ�.꿩��,��I�f��Q����v���ͿS����9���b�Ui)�4�ﾲv����?���ǽ ���	:�v�<�S�<��S;�qü& |��xܽ>#��Z�%#���񟾶����2���������vѯ�'��	���2�P�R��DȽn�T��   �   TӺ<�?=l�)=@��<��Z;��9�>����g��Ͻ��\��H�!��Uڨ��BͿG𿸈� ��ک��=�NB�<$�`������̿����=����H��h�1K����m����;U�5��4g�<̓=��<H=N<�E���1��-�����>��V=���V�&�f�6ik�HBd��R�k6�f��}۽/i����@�˺�   �   ��N=��i=�X=~= �X�LMo�c��s�����ھ��"�C�b����Ƞ��6��Pp�V���&��N/��i2�:/���%����6����=��[Ӗ���d��d$���޾+j���y�A������G�<f�-=.,==Z� =��< �];�u��X�?���U�����-�������v�2�ٽ�̲��m��PX��b/�P�j<�5=�   �   �ٍ=5E�=p0v=P�=�잻�ҍ�\'�B*�����c2���w�yR��+�Ϳ�4�����%�d�4��r?�BC��I?��4�x%�<�����n�ο����'mz���4��q��cۛ��0������r� I�<@9H=�n=:�j=�	H=��=P�< lŸ�%�����\�8��V��0]��M� �&��vܼ��Z<��<�+>=Htx=�   �   �2�=N��=���=d�=�����s���14�+��� ��}<�����M�����׿T����X�-�R�>�t1J�F4N��(J���>���-�v��:s��ٿm���2��V�?�/��u���~>�pV��X\���u�<
�V=�|�=E׊=t%�=�^Z=�=&=���<%W<��:0  �p,X�X~j�8\4�`Hg����;�O�<�e=.hR=��=�'�=�   �   xz�=Ş�=���=@�c=��<�0+�̡ ��Nw�M�ʾ�����T�
X������xdٿ�m����I�&�()��&�2_�:�G��]�ڿb���ڎ�`�W�^���Ѿ�2��4��L�i� �X���=�s=6Ґ=|�=�H�=���=��b=�%;=��=�#�< �<�[�<ܵ�<��<��<N�=��I=�h{=�A�= �=���=�   �   �0�=7O�=�H�=$�b=���<n�"������q�>�ƾ��J"Q�����O
��e�տ�Y��2�����"E#��@&��>#����֮������ֿL���S��>T�����̾Y^~���
���_� B|:h_=P@p=�;�=Xn�=���=�-s=�J=��=���<E�<@�K< x<PC<%G<h�<X��<`s'=h8]=�m�=�z�=Z��=�   �   V�=:�=EԘ=��_=�ѡ<>r�He�-�a�8Ժ����F���v��8�˿�~�����%�N.����&���(�����NI̿�S������kH�U-���q�l������	D��;�X=N�e=�$�={E�=�c=&�5=T}�<��<@�);��Ֆ�����hƼ4-����C� �/9��v<v� =6tD=�B�=��=�   �   �=�L�=���=f,X=t�<\�ϼfmŽ�eH��L��e���]�4���q���_�����ۿFu��t��X���/�4��3�����B�ۿ�����H����r�%V6����h����Q�]�ڽ����<�=B�Q=ZI]=*�D=��=D��<��������g+��|r�a���{��Hܧ�U��������L����� I��87t<��=p�\=�   �   0=�uc=t�n=��I=L�<`;t�9�����(��ϐ���޾,���~U�q���E ��]ĿV�ݿ��1k���K�B���W��9�ܿ)<ÿ�y��]]���U��c�\��3���x�/�M�����˼H]h<>2=�{2=��"=0��<���;t?��l�G��^�ݽV	�
I�N�)�N�,�;n&�T�������ƽ�C��HG
� ?n��W�<�   �   �8<��=(6=<�1=t��<�,��6.c�)#���l�"K��ݥ�95��=i�J��Kè�����п�rۿ��޿=�ڿ&fϿSҽ�%���IW����g��4����蹾�o�|	��{���;���<BC=f�=(�<�>����W�����f�!��M�ias�~���ّ��{��R7���k��1@j�!�A���2Oͽ�k�\e���   �   ,�É;`�<��=4�<��; �����vV6�t����#׾�p�;C?��il�PՋ��Ξ�����ȶ������"���g���i���n��C�i��V=����oվ쑾:Z6��Ľ`� ۱:���<� �<��<`<ػ�J)�v������L�x��TƤ��	��!Xվ ��y�澯��gҾ�`��D#�����v?��e�}����   �   _��PU���;���<d~�<�ql<�f�2hx������Z��~����(���:��I^�Mx}��ۊ�Mr���֔�iؑ�ŉ�ڴz�C[[�8�����)~����V��=����s� �l�8�J<`�<�6�<�D��Ώ#��'��^��2'g��q���
ɾ@J��[����$$$�l�&��0#�d.���	����þ�p����[�R��   �   ���J��hZ׼�M�;P��<�@�<`NE;L����T������Bl��R����߾�����(��iA� �T�r�`�rd��_��R��>�B�%�/�	�fpھ�v��p�c����`D��TK׼�o�;���<�=�<�E;h����Z������Hl�tV��S�߾�����(��mA���T���`�6vd�
�_�ɪR���>�m�%���	��tھz����c��   �   z�V�"D���s��l���J<��<�=�<�����#�{ ��p��� g��m���ɾ�D��X�-��� $���&�-#�+���	�-����¾m����[���t���K� M;D��<t�<0hl<x$f�rqx�����Z�����Y������:�0M^�`|}��݊��t���ؔ��ڑ�<ǉ�øz��^[�8�����
�4����   �   v�]6���Ľ�����:���<�%�<l�<��׻�>)�s��n}�s�L�������������RվC�⾋�������Ѿ�[�����j��Tp?��`�̎��8��;4j�<R�=�3�<�~�;H�����.Z6����>'׾>s�F?�ml�;׋��О�	���nʶ�$����$���i���k��op��e�i�Y=��sվ�   �   8빾[�o�^~	�� {�H�;���<�D=`�=,�< �=�����O��s��M�!�t
M�pYs�*����ԑ�Ew���2��hg��n8j�D�A�>��nEͽtvk�M����8<��=6=��1=ر�<`H���4c��%�T�l��M�����d;5�W@i��K��-Ũ���0�пuۿ�޿��ڿOhϿOԽ�됧��X���g���4�����   �   ��ྺ�����/�얮�4�˼Zh<>3=�~2=��"=8��<���;�&��J�G��塽ڌݽt���B���)���,��g&���4����ƽ;���8
���m�j�<�0=�zc=4�n=��I=��<hIt�`���r�(�xѐ��޾ֶ���U��������ĿA�ݿ-��Ym���L�_���T��	�ܿ�=ÿ*{���^��ʸU� e��   �   ގ�Bi����Q���ڽ����<��=8�Q=�L]=,�D=f�=�˗<@Q��@볼LY+�Hlr�#X��ir���ҧ���v��v�L�(���0��� at<n�=�\=q�=iN�=~��=�,X=��<��ϼ/pŽ�gH�]N��������4�L�q��򙿥���5�ۿ�v��T��D���0����3�L�����ۿʬ���I����r�RW6��   �   �-������l����lD���;PY=��e=�%�= G�=R�c=��5=��<`��<�f*;h��T���0����gƼ ��pzC� ":9Ȱv<R� =�zD=�E�=
�=��=>�=�Ԙ=��_=tϡ<�t��g�ړa�mպ�S���F�9�w��+�˿����&��.�^����B����p��J̿�T�������lH��   �   ���9�̾�^~��
�
�_��<|:�_=Ap=<�=4o�=Ɍ�=�0s=�J=�=��<dO�< �K< �<pZ<�;G<#�<8��<�w'=2<]=xo�=�{�=_��=x1�=�O�=�H�=��b=��<@�"�=����q���ƾ|��"Q�'��
����տpZ����� ���E#�A&�F?#����������ֿ[L���S���T��   �   :��wѾ�2�������i� VX�D�=V�s=YҐ=��=�H�=ۙ�=*�b=&;=��=($�<��<P\�<$��<,�<4��<T�=v�I=�h{=�A�=�
�=p��=dz�=���=n��=��c=h�<n1+�� �DOw���ʾ�����T�#X�������dٿ�m��&��I�&�()��&�*_�0��F��E�ڿ�a���ڎ�6�W��   �    ���̾6]~���
��_���|:2a=.Bp=�<�=�o�=��=1s=FJ=Z�=x��<�O�<`�K<�<pZ<�;G< #�<$��<�w'=6<]=o�=
|�=p��=�1�=�O�=HI�=�b=Ģ�<|�"�4��6�q��ƾ���!Q�����	
���տiY����X���D#�^@&��>#�`����������ֿ�K��FS��� T��   �   {,������l�̊���D���;&\=��e=�&�=�G�=>�c=��5=P��<`��<�l*;x��$��� ����gƼ���zC� :9��v<J� =�zD=�E�=8�=.	�=��=�՘=Ԩ_=l֡<�o��c��a�gӺ���F�/v��z�˿~�d��N%��-� ��x� ����j��XH̿S��Y����jH��   �   ތ�Xf��~�Q���ڽ��� <��= R=�N]=��D=��=�͗<@7���鳼�X+��kr�X��gr���ҧ�*��v����L�P���P���0at<��=~�\=��=O�=���=�/X=��<(�ϼ�jŽ�cH��K������8�4��q���G���z�ۿ�s�����x���.�J��42�)���ɑۿ\����G��&�r��T6��   �   ���E�����/����(�˼�th<�7="�2=�"= ��<���;�$��V�G�]塽��ݽ`���B���)���,��g&���O����ƽ!;���8
��}m�k�<�0=0|c=��n=��I=�'�<0&t�䃝���(�ΐ�t�޾³��|U�Q��������Ŀ��ݿ*��i���J����I��O�ܿl:ÿAx��\��ŴU��a��   �   湾�o�y	��{���;��<J=�=��<�a=����N�����!�V
M�bYs�(����ԑ�Lw���2��rg���8j�Q�A�D��kEͽ:vk��K��h�8<��=�!6=�1=���<0����&c�� ��l��H��K��75�;i��H����������}п�pۿ]�޿��ڿ�cϿBн�G����U����g���4�6���   �   Z鑾$V6���Ľ���ز:���<X0�<��<��׻�<)���� }�2�L�v�����������RվJ�⾗�������Ѿ�[�����s��Vp?��`�����0���;�o�<��=�@�<���;��7����R6����� ׾�n��@?��fl��Ӌ��̞������Ŷ�f���+ ���e���g���l����i��S=���Plվ�   �   ܄V�6����s�`�l���J< .�<�G�<���#�~����� g��m���ɾ�D��X�/��� $���&�-#�+���	�:����¾m����[������I��w;���<(��<(�l<@�e��]x�'���Z��{���侭���:�F^�ft}��ي�p��?Ԕ�)֑���ְz��W[��8�d��y��z���   �   ���R=��<5׼���;�<�M�<��E;����gS��2���Bl��R��}�߾�����(��iA��T�{�`�rd���_��R�"�>�K�%�4�	�lpھ�v��]�c�^���C���F׼���;�
�<O�<`�E;0���N��V��F=l�O���߾���d�(�@fA�!�T�^�`��md�ӗ_���R�v�>� �%�\�	��kھ�r��p�c��   �   q��?� �;���<��<Ȉl<X�e�^ex�&��Z�Z��~��������:��I^�Px}��ۊ�Rr���֔�oؑ� ŉ��z�I[[�8�����"~��؉V�3=����s���l���J<�-�<�L�<�Ő��y#��������g��i��&ɾ)?�U����	$�5�&��)#��'���	�����¾i��(�[����   �   p��X�;�{�<��=B�<P��;��]���V6�R����#׾�p�7C?��il�RՋ��Ξ�ȋ��ȶ�Ʒ���"���g���i���n��I�i��V=����oվ	쑾Z6�E�Ľ���c�:���<�3�<���<`�׻2)�G��Gx�{L�����L�������Mվ��⾰����o�Ѿ�V��V���x��i?��[�T����   �   ��8<��=N&6=F�1=��< ���+c��"�:�l�K��ӥ�95��=i�J��Mè�����п�rۿ��޿B�ڿ+fϿWҽ�)���KW����g��4����蹾ޚo��{	��{���;�0�<�J=H�=��<@�<�Z��gG��o��T�!��M��Qs��Б��r��].��)c���0j�F�A�,��H;ͽ�ek�2���   �   L 0=��c=�n=�I=,'�< /t�0�����(��ϐ�~�޾$���~U�o���G ��_ĿY�ݿ"��7k���K�G���[��=�ܿ+<ÿ�y��^]���U��c�V��%���@�/�����L�˼�mh<48=@�2=0�"=���< 0�;���$�G��ܡ���ݽ���i<��)���,�a&��������bƽ
2��\)
� �l��~�<�   �   ��=�P�=���=�0X=��<��ϼ�lŽ�eH��L��U���X�4�{�q���`�����ۿHu��v��Z���/�6��3�����C�ۿ�����H����r�%V6�����g����Q���ڽ�����<V�=\R=�Q]=.�D=��=�ݗ<@����ѳ��J+�4\r�uO��Ti���ɧ�睽'n��duL� ��� ���`�t<~�=��\=�   �   �
�=��=R֘=��_=֡<�p��d��a�)Ժ�z���F���v��:�˿�~�����%�N.����&���(�����OI̿�S������kH�U-����[�l�.����D��;�[=B�e=k'�=I�=�c=~�5=���<T��<@�*;P�����������PƼD����NC� FD9��v<r� =ȁD=�H�=|�=�   �   �2�=�P�=�I�=��b= ��<��"������q�6�ƾ��H"Q�����O
��e�տ�Y��2�����$E#��@&��>#����֮������ֿL���S��>T�����̾P^~���
��_� z|:�`=HBp=�<�=p�=卉=T3s=(J=ʳ=���<�X�<��K<p�<`p<pQG<�-�< ��<0|'=(@]=)q�=v}�=���=�   �   B��=�'�=T�=�=0�(=Ѕӻ�|��gi*�����9
� �"�&�Z������0��&ɿ��Õ����rb��A�������ɿ������vT]�Ä%�Vd��X����;�x���H�� Hf<N0/=vu=&ʋ=$R�=�$�=;��=�!l=`�Q=�9=v(&=��=��=��=�P,=@VF=l�h=�|�=(�=�D�=I��=�c�=�   �   ��=8z�==7�=qc�=<+=07��|���X&��Ɛ���߾���W�����	X��6�ſ��߿T����� ��,��� �����g�Eƿ��������BY��T"�o���ߗ��6����@���y<�0=�Rs=x\�=UA�=�Q�=D�u=$�X=�:=��=��=4��<<��< v�<@m	=\�$=N~I=��t= ��=��=��=je�=�   �   ހ�=@>�=s��=G��=$�1= ��!������~����}Ҿ����K�S�����~;��!տ~��gJ�������%����迩տ�b��)t��A���pM��ǯ׾�΍�)�(��립�9����<��3=�m=&Ɓ=*r=��h=�wF=��=hE�<�[�<�,<�9�;`�;�F;P��;��x<,�<��=(�W=Cn�=�p�=#$�=�   �   W�=M�=�$�=���=�:=p��;N�R�����r����c0	���9��Eo������&���6ĿLֿ=�῕�忷�ῒ�տ�ÿꬿ�����o���:�&�
�¾ED|����+P��0�S��h�<�y7=��a=�[h=.�S=��*=<T�<��\<����<(�����~70�X�0�fI��輈�n���;x��<��!=�wi=�Ȓ=�   �   �=#��=���=�Ԉ=�B=��c<F��g�ڽ*zM��<��6h�$X#��-S� 2���Ǚ�燮�q���	ɿ?c̿��ȿ4���ѭ��*���ʁ���R�r�#����G�����T��H��dH������<�8=,�M=D�>=H�=�~�< �d
��p8?�D���|ɳ�cѽ���j录Rٽ���l���H�R�(�Լ ��h��<p<=�   �   j1=8/\=�;�=lG{=�[F=T��<0ע������d$�1%��J�Ǿ��	��33�<^�蚃�Ѹ��3ڣ��¬������N��M��oȔ������\��2�-	���Ǿ�ۇ�e(����P켈�%<�	=��2=�.=��= R[<�b>���)� _�� �ݽt+��Z-�M�C��iQ���T��$M��_;��� � > �P���L�[��ȝ��H9<�   �   ��*;4��<(�?=p/Z=�D=4��<��c�0�V�i>���=R��!���޾J���5�h}X��w��{��5����f������������t�d2V�ʥ3����98۾����P����z!`�Hs	��q�<�=.�#=F =��H<�6��b�T��.���W���A��fq���������:��_��P;��.1�����3c�j1���w�����   �   �B� �:����<^�,=Č8==�d<<��ؼ����^�`o��n��ڀ�/b�Ό*��uC��V��%c�-g��/b��#U�A��'�2��+xݾ�쥾��g��N�_ɚ��ɼP�2<�"=��=Lz	=�V�< rT�FX��ҽ;�$��#f��!��i��}UӾ�*��k��ܯ�������q��ξय�*ڍ�4�V�����G���   �   
��lC�@FD;�5�<�"=P=x��<��X��N3��aǽGl'�pv�tڦ�#<Ծ� �K����"��\,�US/�'i+��� �m�WV����;g}��#j����~��:���D;=�<J�"=d=���<@!Y�X3�/hǽ�p'��uv�+ަ��@Ծ� �;����"�`,��V/�sl+��!�G�c[��+�;󀠾�(j�A���   �   &R��Κ�+ɼȚ2<� =��=�|	=�`�<�RT��:X�V�ѽ>�$�gf�������}PӾ]%�Pf������z��:l�ξ����֍�&�V�����?��P7� b2�T��<Z�,=z�8=.�=XT<<��ؼ(��mb�6eo�9r���⾳d���*��xC���V�S)c��g�`3b�W'U�:A���'����|ݾ	𥾇�g��   �   �P����(`���	��l�<��=��#= =��H<h$����T��&���R�]�A��_q�����r��-6������6���,�����0c�m1�
��t������(+;���<��?=�1Z=�D=���<�d���V�,D���AR��$��'޾�����5�{�X�+w��}��! ���h��y���\�����t�S5V�N�3�����;۾����   �   k݇�(�`!���켰�%<�	=��2=�".=��=hn[<�;>��)�9W����ݽ�%��T-�}�C��bQ�^�T��M�$Y;�V� ��8 ��귽��[�����p9<�8=�4\=I=�=�H{=n[F=<��<ᢼ�����g$�C'���Ǿµ	��53��^�n�������ܣ�yĬ������P����ʔ�r���1�\��2��	�4�Ǿ�   �   �����T��K�jiH� ��<$8=�M=>=��=8��<��������**?�����,����Xѽw��`�Hٽ����9�����R���Լ �շ���<<=��=)��=¬�=Ո=(B=@�c<(��<�ڽ�|M�v>���j��Y#��/S�Z3���ș�s�������ɿ�d̿5�ȿ���>ӭ�,���ˁ���R��#�B���   �   i¾KF|����R���S��f�<�y7=�a=X^h=�S=��*=�a�<X�\<�������� � ��(0�H�0��:���輨Mn���;���<\"=�~i=i˒=b�=��=�%�=���=�:=���;��R�\��r�<���1	��9��Go������'��8Ŀ�Mֿ�����#����տL�ÿ"묿�����o���:��
��   �   ��׾ύ��(� ��<��X�<��3=��m=�Ɓ=�t=��h=f|F=0�=dR�<|j�<��,< ��;`X;�9G;���;� y<�$�<
�=��W=q�=�r�=�%�=1��=&?�=믵=O��=<�1=��������p����~Ҿ����K��������]<���!տ���wK��
����&��w�过տlc���t���A���qM����   �   ՘�C���p�6�j	��l�传y<.�0=NSs=�\�=�A�=�R�=~�u=��X=h�:=��=�=4��<���<��<�q	=��$=`�I=��t=���=i��=��=Gf�=���=�z�=k7�=]c�=�+=`B������.&��ǐ�j�߾y��PW�哉�yX����ſR�߿���3� �6-��� ������rEƿ���₊�CY��T"��   �   d꾽X����;����\��pIf<�0/=�u=Aʋ=AR�=�$�=c��="l=��Q=:�9=�(&=6�= �=��=�P,=`VF=|�h=�|�=�=�D�=@��=�c�=:��=�'�=�S�=��=��(=`�ӻ}���i*����s
�D�"�M�Z�����0��:ɿ��ϕ����rb��9������ɿ������RT]���%��   �   ���aߗ�,�6����(��Py<��0=tTs=Y]�=\B�=S�=�u=p�X=��:=��=D�=���<ȡ�<��<�q	=��$=`�I=��t=���=z��=��=af�=ڝ�=�z�=�7�=�c�=+=P0�������&��Ɛ�A�߾���SW�J����W����ſc�߿������ ��,�K� ������࿘Dƿ@��@����AY�T"��   �   k�׾�͍���(��馽3����<@�3=҂m=�ǁ=v="�h=v}F=�=T�<�k�<h�,<@��; \;@<G;@ �;� y<�$�<�=��W=q�=�r�=&�=v��=�?�=���=G��=&�1=�
��������Ӂ���|Ҿ��7�K�ә��y
���:��. տ���hI�������$��}�迳տ�a��bs��a@���oM�-��   �   9¾�A|����:M����S��p�<�}7="�a=�`h=�S=x�*=�d�<H]<����4��P��( �d(0�"�0��:�����Mn���;ĩ�<~"=*i=�˒=��=H�=�&�==:=���;�R�2���r�(��w/	�r�9�lDo������%���5Ŀ�Jֿ���&��F��,�տ��ÿ�謿����?�o�C�:���
��   �   7���z�T��C��]H����!�<� 8=��M=��>=�=`��<@��������(?�~���ҿ���XѽZ��`�Hٽ����=�����R���Լ  շ\��<�<=��=ω�=׭�=�ֈ=B=@d<�����ڽ�wM��:���eﾬV#��+S�1��Mƙ�w���ݼ��]�ȿ�a̿˜ȿ���:Э�\)���Ɂ���R���#�=���   �   Xه�(�������%<�	=��2=�&.=��=�x[<3>�$�)�fV���ݽ�%�YT-�c�C��bQ�Z�T��M�.Y;�]� ��8 ��귽h�[������r9<�9=6\=w>�=xL{=�`F= Ĵ< ʢ������a$�K#����ǾX�	��13��	^����:���wأ�����ϥ���L������Ɣ�}����\�^2�X	�ʤǾ�   �   ^	P���^`��S	�X�<v�=�#=  =��H<����T��%��R��A��_q�z���g��)6������6���,�����;c�n1���Y�����7+;���<��?=B5Z=>D=4��< Lc�@�V��8���9R�S��D޾;����5��zX�zw��y��U���e����������B�t�U/V��3�����4۾#���   �   hJ�Ú�H	ɼ0�2<�)=h�=��	=ph�<xFT�08X�N�ѽ҂$�	f�������oPӾW%�Rf�� ����z��El�ξ�����֍�"�V�����?��p6� �0����<��,=В8=�=��<<�rؼ���Z�$[o��k���|��_��*��rC���V�"c�� g�,b�k U��A�%�'�����sݾx饾N�g��   �    ���t.��?E;lL�<6�"=t=���<��X��K3�i`ǽ�k'��ov�Oڦ�<Ծ� �G����"��\,�[S/�.i+��� �s�aV����;j}��#j����"���8�@�D;�C�<6�"=�=���<�5X��C3�vZǽ�g'�Ejv��֦��7Ծo �s����"�sY,� P/��e+��� ���%Q��_�;�y���j����   �   B*� (���<v�,=*�8=.�=�t<<p~ؼ���.^��_o��n�����%b�ʌ*��uC� �V��%c�5g��/b��#U�A��'�6��,xݾ�쥾��g�dN��Ț�\ɼ��2<>'=��=��	=�p�<�*T�.X�V�ѽ9~$�4f�G������KӾ 꾶`��g���Uu���f�$ξ*����ҍ���V�����7���   �   @�+;D��<��?=
8Z=�D=x��< �c���V�o=��j=R��!��x޾@��
�5�g}X��w��{��9����f������������t�k2V�ͥ3����98۾����P�@��  `�(j	��x�<t�=�#=L =�
I<���f�T�&��`M�B�A��Xq��������1����*2���(���	��c�:1����찚�����   �   �A=�;\=a@�=vN{=aF=���<�Ѣ�����:d$�%��.�Ǿ�	��33�<^�蚃�Ӹ��6ڣ��¬������N��P��sȔ������\��2�.	���Ǿ�ۇ�A(�����8�%<	=�2=�(.=�=`�[<�>�t�)�O����ݽV �PN-���C��[Q�.�T��M�eR;�� �3 �8᷽.�[������9<�   �   ��=��=D��=f׈=�B=�
d<&����ڽ�yM�e<�� h�X#��-S� 2���Ǚ�臮�u���ɿFc̿��ȿ9���ѭ��*���ʁ���R�r�#����A���r�T�,HcH��>�<� 8=�M=��>=��=|��<@q�������?�����綳��Nѽ�y�tU彈=ٽ������:�R���Լ @e����<�<=�   �   ��=��=�'�=�=�:=@��;��R�d��dr�t��\0	���9��Eo������&���6ĿLֿB�Ῑ�忻�῔�տ�ÿꬿ�����o���:�&�
��¾3D|�^���O���S�dm�<,}7=��a=�bh=,�S=�*=�p�<!]< c��\�����켒��0�ts0��+��z輨n� V;l��<F"=t�i=�Β=�   �   ��=�@�=:��=���=�1= C��������l����}Ҿ����K�T������;��!տ���iJ�������%����迫տ�b��)t��A���pM��Ư׾�΍��(�z립 8����<��3= �m=`ȁ=x=��h=<�F=��=�_�<dy�<P�,<`ȟ;`�;��G;@I�;�#y<$5�<��=H�W=�s�=Du�=�'�=�   �   ���=X{�="8�=d�=(+=�1��;���>&��Ɛ���߾���W�����X��6�ſ��߿U����� ��,��� �����g�Eƿ��������BY��T"�p���ߗ��6����X�伈y<.�0=|Ts=�]�=�B�=�S�=Ƞu=��X=t�:=�=��=x��<8��<d��<6v	=��$=P�I=4�t=0��=α�=�=Jg�=�   �   �n�=خ�=j��=&��=��=��<�⼏̽��F�����Ǐ�*!���P�T���r���J�����K1ȿW�˿�1ȿ����W}��)՘�z���hR�i#�iz��{��J�Z�:�����o��B���<B#=$R=p2h=l�m="�h=*�^=�@S=��H=V}A=�?>=a@=2�H=��W=�tm=�ӄ=���=�,�=�X�=���=|z�=��=�   �   ~�=���=~��=<�=o��=���<�Ҽ��Ž��A�X]�� �澁*��L�[D}�ٕ��`��p�����Ŀ�aȿ��Ŀ-�������e(��cO~�p�N��A �E���Ƥ�LIU������d��!#���<��%=�_R=�f=��h=,-a=�T=6yE=��7=�]-=['=2?'=0
.="M<=~3R=]o=;K�=���=�m�=�#�=b]�=^�=�   �   Դ�=��=t��=�	�=�~�=|��<������	4�������پt��B�N4p��G��c⡿(H��a��{q��1���(��Mա��a����p��2C�#��J޾p��n�E��dཀ�D��쓻��<��,=ΉR=�_=�Z=�I=��3=�!=��=�4�<�2�<PD�<`x�<��<�l�<~�=0WG=��u=#;�=v7�=@��=���=�   �   ���=:��=���=��=*��=��=��8�K#�� ��d4���ľ���g1���[��c��⊔��Ǣ�dի�Yி䥫�Y|��LA��Z6��p�[��1�	���Ⱦ�E��d�,��］�h���{;���<�`6=��P=�IQ=�,?=h~ =ؼ�<pi�<��"<���:�hɻp,0�pH�HG&�������;���< ��<��>=Զ}=�=��=�   �   ��=���=-x�=Pۨ=�%�=�!= 	�c��a��a��P���"�Pc�ɊA�L\f�"v���8���O���������Ï��ge�Y�@�w����|�h����A󏽜;�� Jh<�X=��?=�HJ=X:=0k=���<�X<PR�(o������N���s�'���%����h�LN:�`,���3��<0��<�%M=v`�=�   �   �Dp=��=B�=��=��=�@7=~7<d���0ʽ�x6�.����Lƾ4����#�G�C��`�|$v�K��+\�������t���^�K9B��u"����f�ľ�G���[8�ս�y:���F��G�<�d+=LE=��;=�"=�H�<�� ;ୣ�l�4�Y���a#����`���X
��7�6��i꽌տ�ҋ�R %��YA���y<B� =�   �   �� =��U=$��=�]�=��=R�H=�B�<,腼�Z���
��\��A���#Ӿ�~���K7��I��{U�X<Y�J�T��^H��d5����H����ξƒ��G�V�����׋�Ĕ�� �o<,�=F�@= �C=��"=,��<�+�:(6ּ,�n�枾����r�&�2!E�>�\�'sj�Hsm��d�X�Q�R85���5�ֽ�G����@'~;�   �   ��޺ d�<z�E=�s=�_x=hT=��=��;�K#��h��T"�7vo�5���Yξ?"��#��#k���'���*���&����7����8ȾB雾"8c��%�����*��0u�;f=_>=P=�T9=0��<P
�;pƼ�*��j�ڽa��YyQ��:��
ؖ�������C���0������� ���Yq�<_=�/W�_y���� ��   �   ^&�@���&�<��>=l�_=F�V=>M$=`��<`�j�j�e��۽��)��ik��֗��޸�y$־��N�������I��g�
�оl౾'؏��1Z�z���|���&��4��0�<�>=�_=&�V=@K$=,�<�k��e�n۽X�)�rok�Sڗ��⸾�(־�
�S��"����N��2�k�оK䱾vۏ�37Z���������   �   �Ĭ����@E�;j=�\>=�P=V9=���<�5�; `Ƽ#%���ڽ����sQ��7��FԖ������ﱾ޶��㗯�� ����eSq��Y=�|R��q���� ���ݺlq�<"�E=�s=�`x=�T=�=@W;�S#��n���W"�.{o�28���]ξ�&������m���'���*�p�&�/��t9�?��<ȾK웾�<c�d)��   �   ���T܋�`��� �o<��=L�@=��C=��"=|��<���:T$ּL�n�e���d���&�E��z\�(lj�(lm��d���Q�<25�V��xֽ�?�����~;4� =^�U=��=�^�=��=�H=�<�<H󅼻^���!
��\�/D���&Ӿ$�߱�FN7���I��~U�a?Y�B�T��aH�g5����9����ξW���B�V��   �   v^8�Zս�:�@�F�0B�<^c+=BE=R�;=
&=HR�<�c!;������4�>��������4��S
� 2���7_�̿��ɋ���$� (A��z<T� =$Kp=��=�C�=G��=��=?7=(p7<*��5ʽ�{6�B���xOƾ�����#���C��`�U'v�����]������Q�t��^��;B��w"�.����ľ�I���   �   g"h��������C��x?h<6W=6�?=�IJ=d:=�n=���<ht<0综Y��$����N�R}s�������6�h��>:����pT3��5<`��<v-M=�c�=�=W��=Ey�=�ۨ=e%�=F�!= ��^�c� d��a��R��:%��d���A�^f�[w���9��:Q��! ��q���ď�����,ie��@���M��H��   �   �F���,����k��y{;@��<\`6=F�P=JKQ=6/?=�� =���<�u�<�"<���:pɻ� 0�x�G�x&� ���p�;�Ŋ<���<��>=��}=��=!�=J��=p��=���=�=䰆=�=h�8��%�����5����ľ����1���[��d��ꋔ��Ȣ��֫��ᮿ���e}��AB��47���[�L�1����BȾ�   �   0����E�,f�ƛD������}�<"�,=�R=j_=Z=`�I=چ3=�%=޵=T@�<�?�<PR�< ��<��<�{�<��=�]G=��u=�=�=�9�= ��=q��=���=��=���=
�=C~�=���<�!��{��u4������پ�t��B��5p�=H��%㡿�H��5��Or������)���ա��b����p�s3C����K޾�   �   .Ǥ��IU������d��$#�0��<b�%=�_R=Df=��h=`.a=�T=Z{E=@�7=|`-=V^'=�B'=�.=�P<=<7R=�`o=�L�=4��=�n�=�$�=H^�=�=�=��=���=9�=4��=���<T�Ҽ�Žd�A��]������*���L�E}�rٕ��`��߅��U�Ŀfbȿ?�Ŀ����݁���(���O~�ЃN�B �����   �   �{���Z�����b�o��B���<\#=@R=�2h=��m=d�h=|�^=AS=f�H=�}A=@@>=ha@=��H=�W= um=�ӄ=���=�,�=�X�=���=|z�=��=�n�=Ү�=X��=��=��=<��<X���̽F�F��������4*!���P�f���!r��	K�����Q1ȿZ�˿�1ȿ����L}��՘��y���hR� i#�9z��   �   =Ƥ�\HU������d��#�� �<�%=�`R=bf=��h=R/a=hT=|E=��7=a-=�^'=C'=..=$Q<=b7R=�`o=�L�=>��=�n�=�$�=V^�=0�= �=��=���=��=Ԥ�=D��<@�Ҽ+�Ž�A�]�����;*���L��C}��ؕ�9`�����}�Ŀ�aȿc�Ŀ�������(���N~�ւN�JA �v���   �   e���E�=b� �D�@֓� ��<
�,=v�R=�_=�Z=4�I=r�3=0'=$�=hB�<tA�<�S�<��<ܴ�<|�<��=�]G=��u=�=�=�9�=5��=���=4��=��=j��=�
�=m�=|��<�������4�������پss��B�X3p��F���᡿oG������p��_���'���ԡ�Ea����p��1C�I��I޾�   �   nD��T�,�x켽�c� �{;���<jd6=��P=VNQ=�1?=|� =��<�y�<��"<�Ճ:@ɻX�/���G��&����� �;�Ŋ<��<��>=�}=�=B!�=���=���=_��=�=���=��=��8�� �����N3����ľ���?1���[��b��􉔿�Ƣ�Mԫ�9߮�ä��A{��E@��l5��̳[���1�����Ⱦ�   �   �h�S���0��`]h<$]="�?=�MJ=:=�q=���<<`�滸U��v����N�P|s���������h��>:�P��T3�6<���<�-M=�c�=~�=���=*z�=$ݨ=_'�=�!= �빎�c��_�O�a�O��b ��a��A�JZf� u��V7���N��f����	��=���de�k�@���T~�h쫾�   �   X8��ս�q:� )F��R�<�i+=�E=��;=*=xY�<��!;����*�4�#���%���������R
��1���&_��˿�uɋ���$�('A� z<� =�Kp=��=�D�=���=E��=xE7=��7<L��,ʽ�u6�4���;Jƾ�����#��C�e`��!v�����Z��������t��^��6B��s"�ܾ���ľeE���   �   ^���ҋ�T����p<
�=A=�C=��"=���<�k�:�ּj�n���������&��E�^z\�lj�lm��d���Q�:25�V��xֽ�?��,��`�~;
� =��U=��=X`�=�=��H=<O�<�؅��U���
���\��>��g Ӿ,�?��I7�=�I��xU�Y9Y�Q�T��[H��a5�S��8��L�ξ������V��   �   x���
��൧; =e>=%P=X[9=���<�T�;YƼ�#����ڽ"��0sQ�\7�� Ԗ�u����ﱾٶ��ᗯ�� ����fSq��Y=�rR��q��j� ��fݺ�s�<�E=t!s=Pex="T=$�=@";6B#��b��P"�:qo��1��0Vξ������~h�
�'��*���&�к��4�v�� 5Ⱦ曾�2c�p!��   �   
&���|�,@�<��>=�_=T�V=(R$=���<(�j�L�e�j۽a�)�fik��֗�k޸�^$־��N�������I��o��оp౾(؏��1Z�n���|��D&� �~�p4�<��>=�_=�V=�S$=��< �j���e�n�ڽc�)�Kdk��ӗ��ڸ� ־�I��ԇ���D���龒�оnܱ��ԏ��+Z����[u���   �   �1ܺ4��<�E=�$s=�fx=�!T=�=��;�H#��g��xS"��uo��4���Yξ#"���� k���'���*���&����7����8Ⱦ@雾8c��%�����>�����;�=�b>=4$P=,\9=؝�<pz�;�JƼ�����ڽԕ��mQ�24���Ж�x���]뱾�����������N���Lq��S=��M��i���� ��   �   � =��U=��=�a�=��=��H=PJ�<ⅼ>Y��e
���\�QA��s#Ӿ�v���K7��I��{U�]<Y�Q�T��^H��d5����J����ξŒ��7�V�����׋�D�����o<"�=� A=H�C=l�"=��<�!�:�ּ��n�2��������&��E��s\�'ej�em��d��Q�,5���Goֽ�7��м�@w;�   �   fRp=��=0F�=���=���=zD7= �7<���/ʽDx6������Lƾ&����#�B�C��`��$v�N��/\�������t���^�L9B��u"����d�ľ�G��k[8��
ս�x:��vF�pL�<Fh+=fE=�;=�,=b�< �!; ���v�4�����E���������M
�t,�N���T�_¿�����v�$�(�@��?z<@� =�   �   �=���=d{�=�ݨ=s'�=�!= ����c��a���a��P���"�Hc�ŊA�K\f�#v���8���O���������Ï��"ge�\�@�y����z�h������\9��HQh<l[=��?=2NJ=�:= u=���<��< ��,B��ܨ�D�N��ms�֪�����ڛh�$/:����( 3��c<��<�5M=g�=�   �   j��=<��=<��=��=���=��=ء8��"��ي�G4���ľ���b1��[��c��㊔��Ǣ�iի�]ி祫�[|��MA��\6��q�[��1�	���Ⱦ�E��R�,�T］�g� �{;���<�c6=��P=XOQ=�3?=�� =x��<Ą�<��"<�؄:��Ȼx�/�X�G���%��A��`c�;ڊ<<��<
�>=��}=��=�#�=�   �   \��=��=���=�=p�=<��<������4�������پt��B�N4p��G��e⡿*H��d��}q��2���(��Nա��a����p��2C�#��J޾m��a�E�fd��D��擻l��<h�,=b�R=._="Z=�I=��3=�*=D�=dL�<�L�<P`�<���<���<��<��=RdG=��u=a@�=<�=��=��=�   �   ��=���=H��=��=ं=��<�Ҽ��Žj�A�Q]����~*��L�[D}�ٕ��`��p�����Ŀ�aȿ��Ŀ-�������e(��dO~�p�N��A �G���Ƥ�CIU������d�� #�8��<��%=�`R=�f= �h=0a=zT=�}E=��7=Fc-=Va'=�E'=J.=`T<=�:R=�co=mN�=���=p�=
&�=@_�=��=�   �   ���=���=�%�=���=��=zxX=�JA<� 0��v齖P��x����߾�e�V=8���[�ܟ{��N��N�����N���X����{�˅\��N9�����+1����e�Ί�k�����̻�WV<�E�<LU�<�=l=�R=J=�
=`.=��=�20=އE=`\^=Tcz=漌=̭�=4��=,��=��=���=Z��=��=�   �   �F�=�S�=n�=`�=�?�=[=��V<P@'�϶��@K� "���m۾q��o�4�]�W� .w��⇿2����r��y����ㇿq\w�_wX���5�y1��^�:����P`�(F������1�����(Un<�8�<��<�=L=\��< ��<���<�L=Z=7 =��3=B�J=tf=���=+��=�4�=�B�=r��=l=�=p��=pw�=�   �   �N�=b@�=:%�==��=,��=�db=0ډ<���I<Ͻ*9=�&y��0�ξ���e+�e�L�)Aj�׀�qR���ފ�A��Ϳ��n+j�B�L��+��	�ԱҾ�˘���O�d��#2���޼@��:�x�<�`�<�v=��=_�<8	�<��<�!�<�A�<h��<��<���<2=:�'=l�F=ȧj=�~�=:�=:|�=H��=���=Jw�=�   �   P��=�l�=���=|��=H��=��l=��<�"ͼ9��T�'�g���'⺾���.���:�*V���k�u_y��~��y��(k�I�U�SH:�?������2c��
��5Y6�:�ܽМ_����p�<���<�=3=p=`#�<h2�<��<h�d< e$<�h�;���;�D�;�<�p<���<b�=�$0=Vzc=�U�=�/�=1��=ֲ�=�   �   ���=�F�=���=���=-��=Ԝw=��<X�Y�����d�Rna������Mؾol�z�#�WF<�~O���[�A�_��I[�9�N��U;���"�!���׾`g����e����������� �h/�<u=��="�=�o=��<|�<p��;@D�0�C�X���wμ ��d%��yƼp���pwŻ�@�;8��<�4$=�,h=��=��=�   �   ��=N<�=R�=�d�=��=�)�=Ԅ= � �\�E���ܽ��7�8��-ݴ�{c�@
��4��/�_$:���=��9��.�1��B�����,̱�����;6�2I��>g��l~��[<D�=>(=R0=��=�]�<0%�<�[�;�\5��?޼@/��qi���������\J��������k�V�$��ߣ��@�:,��<ޫ7=*;�=�   �   Td=>�=�,�=���=%؜=� �= k,=8�><�K輫R��"d���S���������ę߾>�J���=�x��
q��&�#����jھ������H����n������ [�;z�<��1=��G=8!@=�=���<��<xM�(q���t�Z��uڽ��_��fN��A�>�V����ѽ�f��p)@�t����!*<6=�   �   ���<��N=���=���=׹�=婀=��>=L �<@"%�xO�
�ʽ�����[��ύ�d����Ⱦwݾ��꾀���辅gپ:¾�\���[����I�������E� �9���<\9=��^=��b=��H=P=\��<@Z߻, ��:��՛н��-.���K�s-b�F]o�0�q�ۥh�s�T��8�C���n۽,���4����:�   �    W��}�<PyA=��s=Gu�=R@v=��H=$9�<���;�Aټ׃���۽�i��>N�J.}�xC���G��#������ c�����������i��7����O��VD��L交��< ~A= �s=\v�=6Av=6�H=5�< {�;hNټ�ۃ���۽�m��CN��3}��F��:K�����Ɏ���f��>��7�����i��7�;���V��O��   �   �N� ��9,��<0X9=��^=��b=��H=�=��<�2߻����5��[�н��m.���K��'b��Vo���q���h�j�T�8�U��f۽���(����:d��<F�N=ư�=j��=���=	��=��>=��<�5%�bO�6�ʽ���F�[�_ҍ������Ⱦ{ݾ���ǹ���zkپ�=¾�_��g^��O�I�6������   �   )���d���.�;�q�<��1=��G=v @=&=x��<��<PM�Ri���t����vmڽ � ����II�Z<��7L��y�ѽ�^��Z@��o���H*< >=�d=��=^.�=���=�؜=� �=xi,=��><�V輾V���f���S�������:�߾3�k���?����Bs�)������mھ����������H�Ĝ��   �   �M��Eg�P�~��	[<6�=(=0=��=`�<*�<p|�;`E5�00޼@6/��ei��|�� ���iB���	��������j���$�ƣ� ��:x��<ڳ7=d>�=~�=@>�=��=^e�=:�=�)�=ʂ= �!�4�E�>�ܽ��7��9���ߴ�wf��A
��6�1�/��&:�5�=��9��.�����u�ᾎα�l���>6��   �   �������@J�l)�<�r= �=��=6p=��<�<��; �C���C�PF��Xcμp��X�4aƼ�扼Ż���; ��<:=$=V4h=%��=���=���=!H�=���=p��=B��=�w=���<8�Y��⋽g�&qa�����SPؾ�m��#�/H<��O���[�Z�_��K[�$�N�CW;�J�"�s��I�׾ i��`�e��   �   �Z6���ܽ�_�($��P�<Ą�<��=j2=n=%�<6�<��<�e<�y$<`��;��;���;h�<pq<x�<д=r,0=z�c=Y�=h2�=z��=���=���=�m�=D��=ֽ�=<��=��l=|�<t)ͼ�;��"�'������㺾��a����:��V�E�k�6ay�_~�Zy�S*k���U��I:�W��� ���d��+���   �   ��O�S���3����޼�C�:�u�<d^�<v=`�=�_�<p�<��< '�<|H�<���<4$�<��<�7= (="�F=P�j=e��=��=O~�=��=8��=�x�=|O�=A�=�%�=l��=��=�cb=�։<8��J>Ͻ�:=�z��l�ξ���M+�p�L�QBj��׀�S��Mߊ��A��`���u,j�,�L���+���	�ԲҾS̘��   �   ZQ`��F�S����2������Qn<D7�<8�<|=TL=���<@��<���<�N=�=�9 =P�3=2�J=tf=-��=���=6�=�C�=~��=X>�=0��=x�= G�=T�=Bn�=m�=�?�=p[=(�V<B'����AK��"��ln۾����4���W��.w�ㇿ�����r��˻��䇿�\w��wX�]�5��1�@_ྖ����   �   ��e�����j����0̻xWV<�E�<8U�<�=�=�R=\J=6=�.=,�=�30=X�E=�\^=�cz=��=�=R��=F��=,��=���=h��=��=���=���=�%�=���=��=,xX=�HA<L!0�Dw��P��x����߾�e�p=8���[��{��N��	N�����N���X����{���\��N9�v���1���   �   �O`�~E�����D0�����hYn<�:�<t�<
=�M=d��<ة�<<��<�O=~=`: =�3=��J=�f=K��=���=*6�=�C�=���=j>�=D��=$x�=6G�=>T�=xn�=��=.@�=�[=�V<>?'�!��z@K��!��Hm۾.���4���W��-w�i⇿忏�Er��%���sㇿ�[w��vX�z�5�1�^ྦྷ���   �   �O�9��X0��H�޼�̍:}�<0e�<,y=^�=�e�<��<��<x+�<�L�<��<'�<H��<�8=�(=��F=��j=���=��=j~�=,��=Z��=�x�=�O�=bA�=&�=��=���=�fb=|މ<԰��:Ͻ8=�kx��>�ξ^���+���L�+@j�uր��Q��ފ�i@��2���G*j�8�L��+�<�	���Ҿ�ʘ��   �   $W6��ܽڗ_����h�<$��<��=�6=�=�,�<�=�<���< e<��$< ��;��;`��;0�<�q<��<T�=�,0=́c=>Y�=�2�=���=��=��=@n�=���=���=���=V�l=0�<dͼv6����'�M���຾S�����ߚ:��V��k��]y�� ~��y�'k���U��F:��������a������   �   J��򙫽���@���7�<By=��=�=:u=�<�<�-�;�kC���C��@���^μ��漠
�0_Ƽ`剼�Ż���;���<~=$=�4h=U��=ʎ�=���=�H�=H �=���=���=~�w=���<�Y��܋��b��ka������Kؾ!k���#��D<�#|O���[�5�_��G[�>�N��S;��"�����~׾ie����e��   �   �C⽚6g�@R~�p0[<<�=(=l0=x�= k�<p4�<p��;�35�(޼�2/�ci��{������A��3	�������j���$�tţ� ��:$��<F�7=�>�=��=�>�=��=�f�=��=,,�=�=�R���E��ܽ��7�6���ڴ��`�j>
��2� �/�2":���=���9��.�5��|����ᾗɱ�j��V86��   �   '���$��p��;���<�1=�G=�&@="=���<<��L��d���t�* �� lڽ�� ����H�<��
�L��T�ѽ�^��@��n���J*<�>=`d=.�=4/�=ყ=uڜ=M#�=�p,= �><\;�}M���`���S�B�������`�߾T�5��^;�9���n��$�0���gھ�𲾈�����H�a���   �   t;� +�9<��<�a9=�^=��b=�I=T =�ɍ<�
߻>���3��p�н���.���K�'b��Vo���q�]�h�V�T�8�J���e۽���~(� ˾:���<f�N=���=���=e��=���=��>=L.�<� %��mO���ʽ����[��̍�'���7Ⱦsݾp��>���|cپ^6¾lY���X���}I��������   �   ����<��A=��s=y�=�Fv=~�H=�C�< ¯;�8ټ�ԃ���۽�h�!>N��-}�BC���G����銯��b�����򓋾�i��7����O���C��7交��<�A=8�s=�w�=�Ev=��H=G�<�ܯ;.ټу�8�۽te��9N�b(}�/@��D��`��)���:_��������{i���6���H���8��   �   ��<2�N=���=��=B��=Ϭ�=��>=�)�<�%�tO�4�ʽ����[�Yύ�*����Ⱦ�vݾ���v���辂gپ:¾�\���[����I�v�����E� ��9\��< ^9=h�^=
�b=�I=L!=�΍<@�޻���/����н:�N.�ښK�^!b��Po�7�q��h�L�T�v 8�D��)]۽���b�@�:�   �   �d=��=�0�=��=ۜ=S#�=�o,= �><�D��P��`c�1�S�k���R�����߾.�A���=�x��q��&�&����jھ������H����6���h�㼠c�;,}�<�1=$�G=&@=v=���<� <(�L��]�j�t�Q����dڽk� ����D�7���8B��<|ѽ\V���@��V���r*<�F=�   �   z�=�@�=��=sg�=b�=,�=l�=  �v�E���ܽ!�7��7���ܴ�Qc�@
��4��/�_$:��=��9�	�.�2��C�����+̱����;6�I�6>g�i~�x[<.�=(=H0=H�=�l�<�8�<ྒྷ;5�D޼�)/�0Xi�Nu�� ���:��R��������j�H�$������ ;���<\�7=�A�=�   �   ���=#J�=T�=,��=��=�w=���<`�Y��ދ�~d��ma������Mؾbl�q�#�SF<�~O���[�D�_��I[�=�N��U;���"�!���׾^g����e����x��������D2�<4w=��=`�=|u=t �<��<�I�; C� sC�1��\Lμ��$���GƼ�͉���ĻP��;@��<.F$=<h=p��=W��=�   �   x��=To�=���=$��=���=ܸl=��<ͼI8����'�C���⺾����$���:�)V���k�x_y��~��y��(k�K�U�VH:�?������/c����'Y6��ܽ\�_�`��x�<���<P�=.6=�=4.�<8@�<��<�e<��$<���;�I�;���;8�<X'q<<#�<H�=^40=��c=Z\�=05�=┽=���=�   �   �P�=B�=�&�=P��=��=.fb=�܉<^���;Ͻ�8=�y�� �ξ���a+�e�L�)Aj�׀�rR���ފ�
A��ο��n+j�E�L��+��	�ұҾ�˘���O�Z���1��4�޼ ��:hz�<`c�<�x=6�=f�< �<� �</�<dQ�<X��<�.�<���<D==�(=��F=��j=僉=��=d��=���=Ȼ�=�y�=�   �   �G�=�T�=�n�=��=B@�=�[=0�V<�?'�����@K��!���m۾o��m�4�[�W�!.w��⇿2����r��{����ㇿt\w�`wX���5�z1��^�8����P`� F������1���� Wn<�9�<��<�=�M=ث�<���<���<�P=�=�; =3=��J= f=m��=ּ�=B7�=�D�=~��=4?�=���=�x�=�   �   0>�>���=�=]g�=���=PE3=�'5;��J��*꽑�D�f��$þ������\�,���>�U�J���N���J��?��-��h����ߺǾ�◾��[��_�����:Mh�$��2����,�Ђ�8	)��fH�eX�bG��r�@���0�;��<�@�<$W=M=��{=��=��=`�=���= ��=���=
� >��>�   �   ��>i>L�=|�=p	�=��=r�5=�]�;�aB�y�㽧D@�wa��}B���@�h��:�)��p;�	�F��J��F��q;���)��w�����þlr���4V���y���Z�\����Xx���p �P,�8�2��_H��C>�P��`�?�`��;`�g<���<8�=J@=@n=���=0ۣ=(9�=<a�=`��=r��=T��=r�>�   �   �& >���=�&�=���=.��=�К=�b==P#�;�!*��ѽ�[3�a�������m��
��7 ��31�b<���?�i�;��1��  �1�
���澒;��9y��HF��d��S����;�\N���T��@K��`��̋��*컀,���&���𫚻 �:h <*�<��<�g=lhC=�ho=���=P5�=�̹=�=�%�=�4�=�O�=�   �   X��=��=��=$��=��=��=�G=X�S< ���ĵ����e�n�����bоy��ɳ�&?!��-+�o�.�=�*��� ��,��@���Ͼm����u�fl-��?�X���̞��}?� ��9p~�;0��;`L;��辻(��X��(������������;0�C< ť<p!�<l#=��P=�= J�=|֯=���=ʁ�=�]�=�   �   ��=���=���=�<�=��=D��=r"R=��<,%��������1CM�"���'���ܾ���B����=���P��5�.y����پ?���c鋾�kN����װ�H<��̉��C;�L<�<h�q< ](<�f�; q�0m��OL��}�T`���o�� �p��S2�pR�� �*;@�I<�b�<ܼ=&BO=V-�=Qu�=`�=�/�=�   �   9�=�O�=�5�=j��=,'�=l6�=��Y=���<�e/�d�^�� ٽ�(���j��Y��h����վN�����B ������\�Ѿ�����[�� Ia���!��Խ~o��+�����:��<0�<��<��<�v�<�[< 8�8H��d/��<�ܼ��
�nn ��U-�Ry/�d$%��8���μ�S�@;X	�<r�=$~Y=V،=�;�=�   �   �E�=}�=J��=��=���=N#�=��[=|G�<�� �n������pJ�`q:�:r��	���᫾�����ʾ_R;}�ǾN���ܥ�4���|&a��(����	�� �� ��9�ݮ<p
=�_#=��!=,G=���<��\< ����Fo�T��05���m�ɺ���!�����6ޱ�+Y���3��@.x�T/�X��� 4�l��<|H-=ZQv=�   �   ��W=���=���=V��=ĩ�=	
�=�V=v�=`�;�\���k�@XŽ�}��19�s	c�⃾ 
������[���h���;$��V�v��M�2y�N�⽸ҋ�`7�� ��9���<�&=L�M=0�Y=�M=��-=P
�<H�p<��m���ļ��;�e���H���6���n�Rw�0"��$�����3zɽ�w����5�蔄���)<
=�   �   H��<�q>=�1q=%�=� �=6,s=ƟF=�l=8�Q<��5�� ������g̽����r%���?�R�S��9_�Bw`��5W�\D���(��\�q�Ž�\x��1ۼ sN; ��<nw>=�6q=�=Q"�=j.s=�F=�l=ȏQ<��5�t�U����l̽¾��v%� @�3�S��>_��|`��:W�iD�D�(��`���Ž�hx�Fۼ`�M;�   �    E�9L��<
�&=�M=��Y=P�M=��-=`�<(�p< �m���ļ��;�s���vC����⽈��pj��r���F �!���/rɽ�p��J�5�d����)<�
=�W=6��=���=���=���=�
�=*V=�=@P�;\d���k��\Žƀ��59��c��䃾���x���`���_���'����v��M�2}�	��J؋��I���   �   x�� ��9�Ү<�=�[#=��!=�D=X��<H�\< D�� >o�@��45���m�ʵ��������ױ��Q��e,�� x��F/�P��� �����<*P-=�Wv=qH�=6�=���=�=n �=�#�=��[=�D�< P�"��/����L��t:�>r�F���䫾�����ʾ�U;��Ǿ
Q���ߥ������*a���(��������   �    o�48���/�:���<��<p��<\��<�r�<W< ��8���*����ܼ��
��f �|L-�o/�F%� -�h�μ�{S�`�;��<��=��Y=zی=x>�=6;�=�Q�=O7�=p��=�'�=�6�=*�Y=\��<�r/���^��ٽ��(���j��[��|j��Y�վV��3���� �&���"��Ѿe����]��~La���!�iԽ�   �   ^۰��<�։� ;x�L<��<��q<(T(<�Y�;�{��k��IL�`�}��W���d�� �p�52�����+;�"J<�s�<
�=�IO=�0�=8x�=���=�1�=���=��=���=�=�=n��=N��=�!R=��<�+������f��EM��#���)��6ܾ������@�����JR�7��{����پ)����ꋾ$nN�:���   �   kB㽶���΢�(�?� \�9�g�;`s�;�*; ��ﾻp���|�x��@������@5�;X�C<Dѥ<4.�<�$#= �P=�=�L�=�د= ��=���=d_�=���=��=|�=���=:��=��=�G=��S<(��9ǵ������n�a¢�оv����]@!��.+���.�}�*� � ��-�kB����Ͼ�����u�'n-��   �   �e�iU����;��S���^� dK�`��ڋ��5��/� �&��������'�:�
<�0�<���<�k=�lC=�lo=
 �=M7�=�ι=��=*'�=�5�=�P�=H' >P��=>'�=@��=F��=`К=�a==@�;$*�Z�ѽ�\3�9������o���
��8 �g41�N<���?�O�;�b	1�^! ���
��澀<���y��BIF��   �   v�]�����\����`x����p*ﻀ0���2��aH��C>���� s?����;�h<t��<\�=�@=�n='��=Oܣ=<:�=2b�=>��=2��=���=��>�>Hi>NL�=��=p	�=��=��5= U�;�cB����tE@��a�� C��LA������)�q;���F���J���F�$r;��)��w�|�����þ�r��I5V��   �   �_�����lMh�~��3��x�,�X��X
)�gH��dX�(aG�@q����06�;, �<0B�<�W=�M=T |=�=��=��=���= ��=���=� >Ț>0>��>���=�=Ng�=���=E3=� 5;��J�Q+���D�$f��3$þ������n�,���>�[�J���N���J��?��-��h�����ǺǾ�◾x�[��   �   X�������\�Ȼ�x�H~�`ﻐ'�H�2��XH��:>��~�`U?����;x
h<Ї�<L�=N@=:n=`��=|ܣ=[:�=Pb�=P��=H��=��=��> �>Yi>�L�=��=�	�=e�=P�5=�e�;�`B����.D@�(a��B��@���ߋ)�+p;���F���J���F�<q;�,�)�w�4���{þ�q���3V��   �   �c��Q���;��I��L�`K�@;� ���컸���&�����������:�<$5�<$��<Dm=�mC=�mo=^ �=�7�=�ι=��=N'�=�5�=(Q�=b' >���=�'�=���=��=kњ=�d==�6�;�*���ѽ�Z3���������l�v�
�7 ��21��<���?���;��1�� �q�
����x:��Qx���FF��   �   �<�헆�ƚ�p?� ��9���;��;`�;�F�������g���P��� ���PN�;`�C<@ե<@1�<&#=�P=\�=M�="ٯ=L��=Ѓ�=�_�=���=F��=�=Z��=B��=[��=,�G=0�S<���µ�=��A�n������о������>!�^,+�.�.���*��� ��+��>��R�Ͼ���>�u�xj-��   �   E԰�^<���`�;��L<t��<Pr<Hq(<���;`��P�0L� k}�tM���[��@�p�)2�`��� �+;8(J<�u�<��=0JO=�0�=lx�=��=2�=��=���=F��=�>�=���=�=�&R=d(�<���k���_��@M�n ���%���ܾ������K�����SO�H4��v��Z�پ,����狾�hN�����   �   zo���� ��:��<�#�<���<���<���<�v< `�8|�L�� xܼ.�
�b ��H-��k/��%�+�|�μ�wS�`�;��<|�=�Y=�ی=�>�=�;�=6R�=8�=h��=2)�=�8�=��Y=8�<�J/�4�^���ؽ��(�
�j��W���e����վM��ԁ��� �����꾅�Ѿl���hY��CEa���!��Խ�   �   ��케&:H�<�=�d#=(�!=M=̞�<h�\< 0e��o�X���5�"�m�m�����p���ձ��P���+��x�F/�8��� $����<�P-=^Xv=�H�=��=���=	�=��=�%�=Z\=4T�< �����]���DG��m:��5r�`��0߫��}���ʾO;F�Ǿ�J���٥�����"a�T�(�������   �    ��9���<��&=��M=v�Y=��M=��-=$�<@q< )m�p�ļN�;�o����@����⽜���i�]r�<��������qɽ_p����5��~����)<$
=��W=���=U �=糟=Y��=��=�V=J�=P��;@J��k��QŽ,z��-9��c�W߃�9��y���D���Z���T!����v�M�u�7���̋��#���   �   ���<�}>=<<q=��=�$�=�3s=@�F=�s=ȰQ<�5��������d̽r���q%���?���S�@9_��v`�T5W�0D�w�(�z\�G�Ž@\x��0ۼ`zN;T��<Px>=�7q=��=�#�=�1s=�F=~s=�Q<�5��������`̽���`n%���?��S�:4_��q`�0W�(D�ʨ(�BX���Ž�Ox� ۼ@O;�   �   ��W=��=B�=d��=t��=}�=:V=�=В�;�P��,k��UŽ�|��09��c��ჾ�	��U���:���O���)$��=�v��M� y�$�⽉ҋ��6�� I�9���<0�&=֕M=d�Y=(�M=�-=@�<Pq< m���ļ��;����I<�����:���e�.n�����1����iɽ-i��:�5��h���*<�
=�   �   ]K�=���=L��=Z
�=��=H&�=�\=�R�< ���^��O���`I�lp:�O9r��	���᫾_����ʾKR;p�Ǿ�M���ܥ�/���m&a� �(�������8�� 9�9\߮<�=xa#=r�!=�J=���<��\< �c��o����5�T�m�������\��2ϱ��I���$��Bx� 9/��}�� ���˲<8X-=�^v=�   �   �=�=�S�=N9�=Z��=�)�=�8�=N�Y=� �<�T/�`�^���ؽ,�(��j�}Y���g��e�վ1�����< ������Y�Ѿ�����[���Ha���!��Խo��*�� ��:��< �<\��<Ш�<�~�<�q< ��8�y�����qܼl�
��[ ��@-��b/��%�T ���μ�LS��c;t0�<��=8�Y=�ތ=HA�=�   �   ~��=���=@��=F?�=��=3�=&R=�%�<���r������BM��!��n'���ܾ����9����;���P��5�-y����پ<���^鋾}kN����װ��<�tˉ��O;��L<<�<@r<�i(<��; �@Q�-L��c}�`G��TS��`mp�(2������$,;�HJ<؅�<b�=<QO=4�=2{�=l��=
4�=�   �    ��=,��=��=Գ�=���=b��=��G=X�S<����õ�|����n�����>о`�����$?!��-+�p�.�>�*��� ��,��@���Ͼl����u�\l-�z?�6���^���{?� X�9���;Д�;@p; u��Ⱦ����8g�����t���J��pj�;��C<ߥ<�;�<�+#=h�P=�=�O�=fۯ=G��=|��=a�=�   �   �' >&��=(�=��=+��=pњ=Ld==�/�; *�Дѽ`[3�A�������m��
��7 �31�_<���?�h�;��1��  �2�
���澒;��6y���GF��d��S��h�;��M���R��4K� P�P�����X"�h�&����`������:�<�8�< ��<p=�pC=4qo=�=.9�=pй=@�=�(�=7�=
R�=�   �   '�>vi>�L�= �=�	�=q�=<�5= d�;@aB�)�㽄D@�ga��rB���@�e��8�)��p;��F��J��F��q;���)��w�����þlr���4V���k���:�\����`x�����ﻠ)���2��ZH��<>�H���Y?���;hh<���<�=X @=ln=��=0ݣ=;�=�b�=���=���=���=��>�   �   ��
>"?	>i�>(��=H4�=9F�=7�=�z= |8���=�ެνJ1'�p$m�K󚾿d��}޾�G��ι�(������o��t�޾�;���ʞ� {��*>�B�
�v`Ž卽fj[�.�C�ږK���h��0��Xt��h~��YϮ��i���^1}�:9��yּ��û(�i<H
=�JT=F��=�R�=>#�=�X�=��=���=��>�E	>�   �   PX	>�->��>B@�=��=Q��=�,�=�=��F:<	7�|zɽ�#�9h��՗������پbq�
&����U�Bu�d8ھ�#��S?��fu��*9�4|��V�������-P���8���@���]��������-d���i���um��lox��6��׼0!ڻ��U<nR=F(L=^u�=�=�i�=���=8��=��=g�>I�>�   �   
|>��>
>N��=��=`k�=�Ɗ=�+ =��[;f�#�����F���Z�ێ������*;�v�Zb�!m�����s�̾�D��������c���*�	����ܩ�j�k��m/�p^��q!��=��Id��L�������a�������|k��v1��^ۼ����<L�<��2=�s=u�=g��=���=��=��=�j�=�I>�   �   l��=^g�=�K�=���=d#�=��=;?�=��$=��;���_^�����vrD����c��6����ξ1Bܾҥ��۾?�;#2��ȝ����4�H������νս��:l3������мġ༾����1�POX���w�H�������z�1Z��Q,�l	�@�_�@�:(�<D=�gB=�{=��=�8�='��=�1�=���=TQ�=�   �   ��=���=���=�E�=!�=�Ǭ=�{�=��&=(.<Uм�
�����a�)��`�.0��q������O3��E�¾Jݽ�},��Q��$e���FY��&��7�F���hBA�L�ּP�g�@W#���F����p��9�=�ԖU�fR`�|E\��zJ��-� ������H�!� f>;K�<HE�<6�1=�qi=غ�=��=���=���=�^�=�   �   d�=X��=<��=nm�=��=B��=T�|=4##=�X<|;���^�%0½,����:�c�f�0��������ߞ�6S�������f��.���8X��+�U>��O���<�N��yƼp�Ļ`�;p��;�|�;�AѺ�2����x\��*��ޔ6�6]B��WC��:��*)��3�$�� ��p�뻀k�;X�<��=ԲB=�I}=�ϙ=�u�=LW�=�   �   �ʱ=O��=0�=���=2ި=��=��d=Tp= Sa<��S���0� 5���)�l{��9��CW�rNn��{�QY~��Lu��ra��D���!����+﬽��O�����  �8P|<�~�<0 �<�a�<�w�<`��;���t~��8޼`�>4�TvK��[�ܕb�a��U�X?��|�xQ�H�a�@��:�A�<�=^>T=��=w�=�   �   e�=�֚=�x�=��=�ߐ=b`y=bB=�l�<G9<��/�,N�P�y�������"����$�8�4�;I=� (=��4�ʌ"��!
���ٽ�(���:�p��p��;HQ�<�=2f1=H�5=4N&=�=�i�< `<𭂻$ђ��]�j�6��!h�J􉽳雽Ɖ���X��D��L���$���#^�jM�ܢ��`�q;h.�<d^+=T�i=�   �   :!B=��i=\�|=��{=�%h=(�D=�:=R�<P:�;�J��!����M��+��ͳ�S�ս�����[�Z{���񽜉ҽ����Z�p�t�	�@��0�_<r.=B'B=b�i=D�|=<�{=�)h= �D=:>=�W�<�I�;�J��#��f�M��-��qг�էս9"�,��1_��~���񽓐ҽr��,q���	����`�_<�'=�   �   @D�<H�=�`1=8�5=`I&=��=�a�<�Q<�Ă��Ԓ�2^��6�Hh���"曽R���gS������9�����
^� B�,����!r;�>�<re+=x�i="�=.ٚ=�z�=��=Q�=�cy=�dB=�p�<�J9<�/�8P�P�y���"�������$���4�'M=�2,=��4���"�<%
�]�ٽ�.���:��*��0��;�   �    Ѝ8�{<�s�<���<xW�<�m�<�q�;0.�������޼��4��tK�[���b�*a�ڟU��N?��r�l=���a����:LS�<��=LET="��=�=�̱=b��=�=J��=�ߨ=���=��d=dq=Sa<p�S���0��7���-��}��9�/GW�fRn�]�{��]~��Pu��va�۴D�#�!����]�����O�ԙ���   �   �Ƽ�Ż��;���; S�;��Ѻ3�P����d��h����6�^B�WC��:��&)��.���༴������P��;<!�<��=�B=�O}=�ҙ=mx�=~Y�=�e�=��=���=�n�=��="��=��|=�##=@�X<�?����^�3½*���;���f��������➾nU��ڱ��i������;X��+�oC��������N��   �   `HA�,�ּؕg�Hk#�hG�x��(�^>�*=�<�U��T`��F\��zJ�b-����,���К!� �>;�V�<�Q�<V�1=�wi=���=V	�=@��=���=r`�=l��=���="��=�F�=�!�=`Ȭ=�{�=��&=�.<�Yм������\�)�t`��1���r��귳�X5��Y�¾U߽�l.�����f��ZIY��&��;����   �   W����p3�����lмp����1�\SX�P�w����������z�|1Z��P,� ���_�@o�:%�<�=6lB=��{=�!�= ;�=���=�3�=f��=�R�=���=Zh�=�L�=@��=�#�=�=V?�=�$=��;��=`��V��<tD�������������ξ�Cܾ���Ύ۾�;�3��bɝ�-�&�H�M����ν�   �   �ީ�ܶk��p/��a�@u!���=�:Md�N��Z
��4���a������|k�"v1�h\ۼH��0<��<��2=�s=�=���=T��=Z��=��=�k�=�I>l|>��>T>­�=B��=�k�=�Ɗ=f+ = �[;t�#�8���S���Z��ێ��¯��+;�w侤c�nn��K�.來�̾�E������"�c�ʧ*�����   �   �W�������/P� �8���@���]������������������m��:ox�j�6�T׼ڻH�U<8T=$*L=Rv�=���=hj�=\��=��=���=��>��>�X	>�->��>v@�=��=\��=�,�=8=��F:�
7�t{ɽ��#��9h�֗�������پr�c&�,�����u��8ھ.$���?��u�c+9��|��   �   �`Žb卽k[���C���K���h��0���t���~��UϮ�bi����0}�99��wּ�û�i<*
=�KT=���=S�=�#�=�X�=(��=Έ�=��>�E	>��
>.?	>q�>6��=D4�=2F�=7�=�z= �8��=�4�ν{1'��$m�h��d���޾�G��չ�,������o��m�޾�;���ʞ�{��*>�J�
��   �   V������,P�H�8���@���]�����ع��NU���)���l��\lx���6� ׼Pڻ(�U<lU=+L=�v�=�=�j�=���=��=Ү�=��>��>�X	>
.>��>�@�=.�=ʝ�=-�=�=�8G:�7��yɽ��#�p8h�5՗�������پ�p�%���� ��t��7ھ$#���>���u�*9��{��   �   ۩�Ȱk�Lk/�T\��o!���=�"Gd��J��$���
���^��"���~wk�Hq1��SۼX���'<d�<��2=@ s=��=M��=���=���=��=�k�=J>�|>��>z>&��=֒�=Xl�=�Ǌ=\. =��[;(�#�Ο��#��3Z�Nڎ������);�u�!a��k������P�̾�C������<�c�Z�*�����   �   ����Th3�����м�������1��JX�Z�w�W��[���J�z��)Z�DJ,����h�_����:T+�<
=nB=��{=K"�=d;�=N��=�3�=���=�R�=���=�h�=�L�=҈�=�$�=�=�@�=8�$=@>�;���~[��O��ypD�a��������k�ξx@ܾ��T�۾��;�0���Ɲ��"�H����.�ν�   �   �<A��{ּ�og�F#���F��������3�f=�r�U�lJ`��<\��qJ�f-���������!���>;�\�<V�<�1=�xi=��=�	�=���=&��=�`�=���=:��=���=RG�=�"�=�ɬ=�}�=��&=..<PHм��������)�	`��.��Fo�����=1��)�¾5۽�}*��x��|c���CY�2&��3�ꎞ��   �   (mƼP�Ļ �;�	�;�;@�кx�2�L���$M�������6�dSB�VMC�2�:�v)��(�`�༤p�뻰��;�$�<��=ԺB=�P}=ә=�x�=�Y�=Xf�=~��=L��=�o�=��=���=��|=
)#=pY<x,��r�^�1+½T����:���f�.���z����ݞ��P��h����d��1����4X���+�9��װ����N��   �    X�8�|<ԉ�<�
�<�l�<p��<P��;@Т��m���޼X�^�3��jK�R[��b��	a�ĚU��J?��o��8༨�a�@��:LU�<��=�ET=n��=m�=/ͱ=���=��=��=��==��=��d=�v=�pa<h�S�:�0��/���#� x��9��?W�Jn���{��T~��Gu�dna��D��!�J����鬽��O�8{���   �   H^�<�=�k1=��5=�S&=6�=�w�<�~<0i��콒�JS�ԭ6��h��퉽�⛽Z���Q������ß�����f^��@�X����-r;�?�<f+=�i=s"�=�ٚ=f{�=o�=X�=|fy=�hB=�{�<�g9<X�/�2D�8�y������g����$���4��D=��#=��4���"��
��ٽ�"���
:�����4�;�   �   r-B=��i=��|=~�{=F/h=�D=�D=�f�<p��;X�I���`�M�a'��Cɳ�!�ս�����Z��z�����ҽl�����p���	���`�_<�.=�'B=*�i=P�|=��{=�+h=��D=�A=�a�<P~�;��I������M��%��sƳ�E�ս<����W�Rw����)�ҽ
�����p�v�	�0����_<z5=�   �   �$�=�ۚ=L}�=$	�=��=:iy= kB=\�<l9<(�/��E�@�y�B����������$�V�4��H=��'=��4���"�h!
���ٽ(��f:�p��p��;`R�<č=g1=|�5=�O&=l�=tp�<�q<����>T�h�6��h��뉽�ߛ��~��mL��n���*���(��^�6�xx�� �r;hO�<�l+=ʌi=�   �   Eϱ=� �=1�=~��=��=V��=��d=*x=hra<��S�p�0��1���&�z��9��BW��Mn���{��X~�:Lu��ra�۰D���!�`�����O����� �8�|<x��<,�<�d�<\{�< ��;��t���޼Z�.�3� jK�,[�@�b�xa��U��B?�
g�@&�(�a����:�e�<�=vLT=@Ç=��=�   �   h�=���=���=�p�=��=f��=��|=�)#=hY<4/��D�^�z-½�����:���f�أ��]����ߞ�S�������f��!���8X���+�->��*�����N�yƼ��Ļp�;���;���;�Ѻ��2�<����T����n�6�&UB��MC��:�V)�
%���䓼�p����;�2�<��=@�B=�V}=�ՙ= {�=�[�=�   �   ��=T��=���=0H�=�#�=Dʬ=~�=��&=�+.<�Kмr�����|�)�2`��/���p��ε��,3��-�¾;ݽ�r,��H��e���FY��&��7�)���BA���ּXg��T#�`�F�H��8 弔7�"=���U�vM`�Z?\�NsJ��-�ޮ�Ј�� |!��5?;�e�<�_�<"�1=�}i=x��=��=���=���=>b�=�   �   ���=pi�=�M�=f��=,%�=x�=A�=(�$=�8�;>���\��J���qD�F��,�������ξBܾť�
�۾8�;2��
ȝ����*�H������ν�����k3�����
м��������1��MX���w��	��ȵ����z��+Z�PK,���鼀�_�@�:�/�<�!=NqB=T�{= $�==�=���=>5�=���=�S�=�   �   �|>:�>�>���= ��=�l�=�Ǌ=D. =��[;>�#��������%Z��ڎ������*;�v�Pb�m�����p�̾�D��������c���*������ܩ�6�k�Hm/�^�xq!���=�Id�L��G��(���_��2���<yk��r1�XUۼ����)<d�<�2=�!s=~�=J��=���=���=��=�l�=[J>�   �   �X	>".>��>�@�=J�=杺=(-�=�=�1G:87�zɽ΀#��8h�}՗�쟺��پ[q�&����T�Au�b8ھ�#��P?��au��*9�2|��V������x-P���8�X�@�Z�]�X���L�������������l���mx��6��׼�ڻ��U<bU=P+L=�v�=;��=�j�=���=j��= ��=��>��>�   �   8�>lV> s>�� >p��=M�=e��=�=V=��;;���B������f�-��7\�Z���p��x��'����	��]������� b�q9�n���t㽽(��������2B��������}���� ���4���B�֗G��B�f#4��c�߁ ��ӿ�H�w���� U;/�<B�]=:P�=��=nI�=<��=��>��>X>�   �   �k>Z=
>_>8�=b��=�=�=bi�=}=>s= �P;&�	��Й�U�����)�x�W��?���`��ִ���6��]����j�������v\�#�4���8�۽mm��d���䆽򒽖��Gٽ:~�h+�K0�]�=���B��B>��60���;���^8����s�x�⼀`;|��<�lY=���=()�=�U�=ș�=d( >e>z
>�   �   T�>d�>=>���= ��=�w�=މ�=d%v=<�=`6�;D���)����潷��n�J��q������!��JA��秐�ۆ�9p�QgL��W&�'��ƽ�֗���x��j����K����ý�{��s���"�q-0�l5���1���$�G��GJ�&��X_h�<ܼ���:TH�< L=Z��=�a�=Q�=,��=l��=�h>ke>�   �   7�>� >z��=�\�=8��=NI�=Ʊ�=��h=�=��;��㼨S����н���
:7�^Y��t��d���ᄾ�B���p���T�8_3�P*�@ݽ�磽4r���?�X�1�,WG���z�\@����̽A]��t��	��� �PN����c��"�׽�У�~�Y��|ؼ r��q�<��3=Ps�=�=~��=��=X�=r6�=  >�   �   ~�=���=n �=~��=\��=��=Fޏ=֛R=��<��y;�˼�f�ÿ��g���ho��S<�.�R��`��Yc���[���J�ڢ1�ҩ����ǳ��\p�"r#�D���qӼ���^*,�o��W����Ž�i� ��2����i���u�`%�������M���ਸ਼���y<&h=�U=�.�=Xͧ=�N�=�X�=���=���=�   �   "��=~k�=F��=>��=���=�|�=��w=�V0=�-�<��::x�ü�6N�􅟽��׽+V���z3.���7���8��1�b!�ԁ
���߽lB��~�f����������M��`�"�hˤ��^T�����"P��Ӌǽ��ֽ��ڽM ӽ�l��nѧ�o���zgK����8>d��}s;Dv�<�'=T/W=���=�z�=�P�=�_�=�=�   �   �ý=V3�=��=^��=�%�=Ʋ|=��A=x��<(5Y<�»��ּ��A��l�������nݽ����@/
���� ��h����0gĽ"�ĒK�Hs�xL����;8�`<4��<��C<`�A;H�#�$�ϼ��)��Eg�Lc��`����b���g��톣����V��N�Y�$�&�d"߼ �T� �:�<�v=
�@=fy=���=���=�n�=�   �   �?�=5��=��=5b�=��h=Z/6=��<�Sv<�e�H�����0�F�f݁��̝��ʵ��Ƚ,�ҽo7Խ1M˽�㷽v�l;m�:���e���8�:8ي<���<L=��=�^
=�H�<pBi< ʣ9`p�PZ�
f.��[�N0|���������S;��B.���x}��b�D=>���`2���S
���;���<L�=��T=�]�=��=�   �   ��g=:�l=:,_=��A=�= ��<0p<� ��lS��D��xC7��;a����E����嘽}-�� ����p�����0_[�4�!�t��������0A<@��<��(=8�P=V�g=�l=2_=��A=�=���<h�<0Ъ�\H�����
@7�$:a����1����瘽=0�������t��s��th[�n�!�8���>���A<0��<,�(=&�P=�   �   =��=xX
=l;�<'i< =�9`#p�|h�l.�r[��4|�R�������;��!-���t}��b��6>�����"���3
��$�;8�<�=�T=z`�=S�=vB�=���=J!�=�d�=�h=�46=h��<Pgv< d����������F�ށ�sΝ�_͵�_Ƚ`�ҽ5<ԽWR˽�跽����DEm�^�(v���F�:\ˊ<���<�   �   ��`<h�<��C<� A;x�#�h�ϼΎ)�pMg�g������ke���i��3���o��VV����Y�&�&�<߼P�T����:D,�<^}=4�@="y=@��=��=0q�=ƽ=�5�=2��=���=�'�=�|=�A=��<XAY<0 »��ּ��A��m��#ö�"rݽ�����1
����|��k�B��hlĽ����p�K���i�P{�;�   �    %������"�d٤�p!�&T��䍽)T����ǽ>�ֽ̋ڽ�ӽ2n��Eҧ�t��� fK���(/d���s;X��<�,=�4W=!��=6}�=2S�=�a�=�= ��=Rm�=��=��=Z��=�~�=��w=BY0=�1�< ;:�üp8N�����2�׽�W����5.���7���8�u1�(!�m�
�q�߽�F��>�f��������   �   ��뼸}Ӽ8����0,�o�|[��m�Ž��H� �|4�e��l��=w�^&��`�����M�@�В��`�y<l="�U=�0�=Vϧ=�P�=^Z�=$��=��=��= �=��=���=���=�=cߏ=��R=8��<@�y;�˼V�f��������(q�V<���R� `�A\c�=�[�B�J�H�1�
�����R����bp�8x#��   �   ��?���1��\G�j�z�pC����̽�`��%�G�p� ��O����!���׽+ѣ���Y� zؼ�|q�w�<��3=�t�=��=���=��=lY�=�7�=� >��>*>|��=�]�=(��=)J�=~��=��h=2=�;,���T����н���;7��_Y�	t��e���ℾ	D���p���T�a3��+�Cݽoꣽ>9r��   �   ��x��
j�7���TM��i�ý[~�Bu���"��.0�6m5���1���$�����J�3&���^h��ܼ��:TL�<LL=���=	c�=R�=2��=`��=i>�e>��>��>�>L��=���=wx�=J��=�%v=D�= 2�;����*��-�潵����J�nq������"��$B�������ۆ��:p��hL��X&�?��!ƽ�ؗ��   �   ����k冽��'����Iٽ�@,��K0��=�,�B�FC>��60���0���8���s����w;���<>nY=w��=�)�=�V�=h��=�( >be>�
>0l>�=
>L_>��=���=�=�=�i�=(}=s=��P;�	�Rљ�Q���U *�0�W�Z@��a��L���.7��Й���j��J ���w\�ʌ4�L��_�۽�n���   �   K�������B��M������֊�� ���4��B�ؗG�ȩB�0#4�Uc��� �=ӿ���w���张j;|1�<Z�]=�P�=��=�I�=|��=��>�>�X>H�>~V>1s>�� >���=S�=\��=�== �;;���SB�������-�8\�m���%p�����1����	��b������� b�q9�{��2u�)���   �   �����ㆽO�i󯽨Gٽ~�+��J0���=���B��A>��50���<���e6��0�s�x����;x��<PoY=߻�=8*�=�V�=���=�( >qe>�
>>l>�=
>\_>��=���=4>�=�i�=J}=�t=�Q;��	��ϙ�_���,�)�عW��?��>`��k���E6��똚�j������Dv\���4�2�s�۽�l���   �   r�x��j�����I����ýMz�s���"�<,0��j5�2�1�<�$����G�#��lYh�4ܼ@S�:�Q�<\!L=G��=�c�=�R�=���=���='i>�e>��>��>�>���=(��=
y�=��=(v=�=�O�;X���'��|��}���J�q����� ��n@�����@چ��7p��eL��V&�$�3ƽ�՗��   �   �?��1��SG�
�z�O>��M�̽�Z������� �BL�i��<����׽�̣���Y�(nؼ�Jp��~�<��3=�u�=l�=���=d��=�Y�=�7�=� >��>N>Ա�=8^�=���=�J�=���=��h== .�;��㼸P����нޠ�	87��[Y��t�\c��q����A��tp���T�X]3��(��=ݽK壽�/r��   �   ���$iӼ����%,���n��T���Ž
�<� �j0�i���d��Tp�B ������M����0e�� �y<zo=��U=�1�=
Ч=HQ�=�Z�=���=n��=B�=l �=D�=d��=b��=�=���=&�R=���<@�y;@�˼h�f����������l�NQ<�\�R��`��Vc���[��J�V�1�������N���Vp�m#��   �   ����$����"�p�����f	T��܍��K����ǽf�ֽ4�ڽ��ҽ�f���˧��|��v\K�x�`d� t;���<�/=�6W=᥈=�}�=�S�=5b�=d�=X��=�m�=���=���=&��=��=��w=0]0=�;�<��<:ܺü�-N����P�׽WS���X0.���7���8�w1�k !�
���߽>����f�d������   �   ��`<��<0D<��A;{#�\sϼ�~)�D<g�,^��٬���\��ua������� ���P��wY�X�&��߼�~T�@E�:�1�<r=� A=Vy=���=u��=�q�=xƽ=�5�=���=&��=�(�=R�|=�A=ܭ�<�VY<0�����ּ��A�%g��1����hݽ�����+
����f���e���콣aĽ핽ЉK��c�1���;�   �   �#=(�=\d
=�T�<�\i< ��9��o��G�[.�t [�z$|����������4���'���k}�b��0>�������`)
�p4�;,�<&�=ƢT=�`�=��=�B�=#��=�!�=`e�=p�h=�66=��<�vv< �b�p���T�F��ׁ��Ɲ��ĵ��Ƚ��ҽ�0Խ�F˽|ݷ��욽�0m����0T���-�:��<���<�   �   ��g=2�l=l7_=p�A=l�=��<��<P���t4��Г�p47��-a�W����������W)�������m������[[���!�������x4A<̯�<R�(=��P=��g=��l=�2_=��A=��=���<��<0���$?�����v87��0a����T����ߘ�_'��ۚ��vj������S[�b�!��齼 ����PA<���< �(=��P=�   �   �D�=.��=�#�=xg�=̢h=N;6=P��<��v< �a�L芼�����F��ׁ��ǝ��Ƶ�XȽH�ҽ$5ԽmK˽[ⷽy��9m�$���c��@N�:tڊ<���<�=V�=�_
=|J�<�Gi< ��9h�o�4T�b.�`[��)|���������X5��d'��zi}�<	b��+>����$���
�0k�;0�<:�=R�T=Wc�=�	�=�   �   HȽ=�7�=j��==f*�=�|=��A=��<�bY<�����ּ|�A��g��Ƽ��rkݽ���.
�������Lh��콞fĽ���K�0rἐJ�p��;0�`<L��<��C< �A;0�#�`ϼ �)�Cg��a��<����_��"d��������Q��~vY�2�&��߼HmT�@��:�<�<ބ=A=Py= ��=���=|s�=�   �   ���=o�=��=	��=���=��=��w=�_0=@�<�&=:��üv.N�1���Q�׽�T�d��2.�1�7�2�8�21�!���
�\�߽$B���f����䊒�`
�J�� �"�<ʤ�B�LT��ߍ�#O����ǽ��ֽ��ڽ��ҽ>i��yͧ��}��>]K�rw�d��@t;���<p3=�:W=駈=��=|U�=�c�=��=�   �   d�=~�=V�=~��=|��=#�=��=�R=X��<��y;��˼��f������Zn�S<���R��`�&Yc�>�[�u�J���1����|�罜����[p��q#����(qӼ����),�f o�\W���ŽH�� � 2����g��s�_"��������M���ἀ`���y<�q=D�U=�2�=zѧ=�R�=\�=Ċ�=���=�   �   J�>�>���=�^�=���=�K�=F��=��h=�= 0�;��oQ����нС�L97�w]Y�vt�bd���ᄾ�B���p���T�(_3�=*�a@ݽ�磽�3r�J�?��1��VG�F�z� @��_�̽�\��3�O	��� ��M���������׽aΣ��Y��pؼ _p�\�<��3=�v�=H�=���=\��=�Z�=�8�=> >�   �   �>�>�>��=���=�y�=���=�(v=��=`P�; ��T(��b��,����J��q������!��7A��ڧ��
ۆ��8p�EgL��W&���ƽ�֗���x��j������J����ý�{��s�r�"�<-0��k5�S�1�V�$�����H�$���[h�Xܼ 7�:Q�<�!L=���=d�=S�=��=$��=fi>)f>�   �   Nl>�=
>p_>��= ��=l>�=2j�=�}=�t=�Q;��	��ϙ�����s�)�?�W��?���`��ȴ���6��W����j�������v\��4���+�۽dm��Z���䆽p򒽊��Gٽ0~�\+��J0�F�=�p�B��B>�N60�\������7��<�s������;Ц�<�nY=���=2*�=�V�=���=�( >�e>�
>�   �   ��>��
>�$>�">�G�=��=�q�=V�=<Bm=4=�
,<�댼�(?�g蜽k�׽���.�.'���+��;'�s!��T	�A\�t���]���Qa��XΈ�˚��]½�h���%�N�Q�j�h����[��<Ʊ��Ƶ��Ǳ��"�����dEz��G��O����|
A� Oӻ��<$�k=�h�=���=�	�=�F�=��>�
>�   �   �
>z	>M�>�C�=X�=`��=^7�=E�=0h=X3=�|#<xΌ���<�k)��emӽS�����=N#��i'��"�����U�:������>3��L�������o���b��){��Z#!��}L�|cy�������z����������h���9���Z/u�* C��A�aO�� �;�P���4��<��j=2�=,�=�5�=�P�=p�>e�	>�   �   �C>Ɵ>��>R+�=�p�=���=�M�=���=��W=��=��<@����5�'���<�ǽ|����J0�Jn����W�
�u��>W̽���q���Z$g�B-b��'��+l߽"��("=��g�2쇾�C�������������똾bP��V�f��U7�����P���e-�П��.�<f=�W�='<�=N��=�M�=׍>T>�   �   �$>��=���=F��=(��=��=��==�=xq:=�J�<p��;Ҙ���.��\��,p���Q޽Ҧ��$H��	�0��=� �Ͻ)���nӆ��S��l/�2�*���I�|:���L������*%�`�L�ğq������!�����(��Չ�Uv�j<P�
�%�m��ջ��<7�����/�<6�\=�-�=m�=���=���=~(�=4� >�   �   ���=8�=�"�=QF�=��=�|�=J��=P�P=�=�5�<���x഼�,��}�t���;�½�wٽl�q"彽�ؽ�.��OG������#>���Pм��Ƽ������<�s.���ɽ0���6*�`uK���f�H�y�Pŀ���}�K3n�.U�;�4��Q��Խ�戽v������L��<�L=j��=��=�#�=tw�=�$�=xe�=�   �   `�=:��=9��=4j�=V��=�`�=��H=|�=<�<@1;��Y����6�*�q���������/������3d�����Y��j�_�l��0
ȼ(�N��_��鍻�7'��0���A1�Xq�Ƚpj�"� �^:9��oJ�yR���P��4E���1�F��v���:���Om��a��,�`=�<$�0=�f{=���=��=���=0��=�&�=�   �   �ɻ=�K�=X�=�ƌ=�se=�+=0+�<x�><@�G�,����Y��)�>�R�h"v�]���$��SO��\7������n�c�&�1��f���r�������<�u�<��<�C< �O:�܄����i��l���5齁M
�,�_�"�`#��Z���|���;�ʽ����YS��2缰�ƻ��m<=F�L=Ń=-��=�#�=!��=�R�=�   �   q��=bȌ=�lr=d�>=p�=�D}<���������	0��,W���s�Q��z�J������P%u��YY���3���`�������<<`f�<�@�<��=n�=f�=t��<p�.< |���<�bpP����F���2eؽ}D뽆4�w��a޽��ƽ����NK��(�I�6��`tg���G;�"�<�@=.�G=.�w=0��=\�=L'�=�   �   ��b=<�C=��=`6�<@RS;�(���b���Q�a҅�J4��UH�����I^���7���Ւ��N����T�#��2ۼp�O� W�:��<Ԓ�<��+=�FQ=~ch=��n=��b=��C=��=xF�< �S;����X���Q�^ͅ��/��0D��)���[��6��WՒ��N��
�T�~�#�$<ۼ�O����:��<$��<<�+=�@Q=�]h=ơn=�   �   ��=��<��.<P���`P� {P�/������jؽ�I�m9��{�e޽�ƽ󑩽�K����I�����eg� 1H;�,�<�E=<�G=2�w=���=�^�=�)�=*��=Pˌ=�rr=l�>=�=Xe}< ��􂉼t���f0�&W���s�cO������k�������(u�r^Y�j�3�J�`,���ū�#<�Y�<\4�<�~=:�=�   �   ��C<��M:�턼l������q���;齦P
�&/�Z�"��b#�]���5�����ʽ߼���YS��/�psƻh�m< "=|�L=Fǃ=L��=(&�=P��=�T�=F̻=N�=�Z�=�Ɍ=�ye=~&+=�8�<غ><�*G��y��HP�`)�b�R�4"v���������Q��,:��­��F�c�"�1��t��s�@;�x�<\i�<���<�   �    S'�@��:J1�󌽿�ȽZm�>� ��=9��rJ�!|R�n�P�7E��1����r���;��lPm��_케��B�<J�0=Lj{=���=��=§�=���=�(�=T�=V��=v��=�l�=୛=/c�=�H=ġ=��<@]1;�tY�����6��q�����t����1���Ĺ��g���!��.]��j�_�" �ȼ8�N�P���@���   �   ������<�y2��uɽ����9*�\xK���f�U�y��ƀ���}��5n��/U���4��R��Խa爽���˟�L��<JL=í�=��=%�=�x�=&�=�f�=(��=��=�$�=0H�=��=�~�=Q��=2�P=D!=�;�<�m��޴�h�,�,}�셣�U�½,zٽo彸%� �ؽ"2���J��� ���)>�����м��Ƽ�   �   t�I��=��sP�����5-%�ղL�b�q�K���
#����()��։��v��=P�Ѧ%�H������6�����2�<*�\=�.�=n�=���=���=�)�=Ȓ >�%>�=���=���=���=x��=��=l>�=�s:=<N�<@��;�ј���.��]���q���S޽5���xI�	����$���Ͻի���Ն��S��q/�j�*��   �   "򁽴��o߽����#=���g�7퇾�D���������с���옾�P��
�f�>V7�ۈ��P��e-�����1�<�f=�X�=�<�=��=vN�==�>yT>YD>4�>�>D,�=rq�=���=�N�=���=��W=��=`�<ı���5����w�ǽ	��r�N1�\o����j�
����BY̽v
��P���8(g�d1b��   �   ,q���d��.}��|$!��~L��dy��������� ��4���B������b���x/u� C��A��N����;� �����<H�j=�2�=�,�=H6�=0Q�=��>��	>M�
>]z	>��><D�=��=���=�7�=��=�h=�3=�|#<Pό�V�<�*��/nӽ������N#�nj'���"�T���V�]������f4��QM��U����   �   �˚��^½j����%���Q��j������[��UƱ��Ƶ��Ǳ��"������Dz�bG�O�����A�PAӻ��<n�k=(i�=��=�	�=G�=ػ>)�
>��>��
>�$>�">�G�=�=�q�=P�=(Bm==�	,<�쌼)?��蜽��׽���..�2.'��+��;'��!��T	�v\齻��������a���Έ��   �   �o���b��%{��P#!��}L�@cy�١���������7���J��ź�������-u���B��@�/M��&�;��w��H��<v�j=03�=-�=�6�=`Q�=ĵ>��	>X�
>iz	>��>bD�=�=��=8�=	�=�h=�4=x�#< ˌ�̂<�u(��clӽ�������M#�@i'�t�"�0��sU�h��-����2���K��Ǿ���   �   �G��-k߽���a!=��g��뇾,C������������꘾JO��9�f��S7�܆��M���_-�w��7�<  f=WY�=�=�=���=�N�=]�>�T>pD>L�>)�>�,�=�q�=7��=BO�=P��=��W=�=�<����$�5�����ǽ/��Y�/�m�z��B�
�{��U̽�����""g�d+b��   �   ��I��8��K��P���)%�ĮL�؝q�����} ������&���Ӊ�z v��9P��%���򽩷���/� ��L;�<F�\=�/�=�n�=x��=P��=�)�=� >�%>P�=,��=���=��=��=��=w?�=tv:=XU�<`ǐ;�Ƙ���.��Y���l��WN޽m���nF��	����+�N�Ͻ����-ц��S�ri/���*��   �   P}��L�<��+���ɽr���4*��rK���f�A�y��À���}��/n��*U��4��N�Խ	∽�������T��<L=&��=��=�%�=ry�=�&�=Pg�=v��=.�=�$�=�H�=B�=t�==��=��P=�$=$D�<��PѴ�>�,�v}�L����½Jsٽ�g�L彽ؽ+���C��`��J>���\�ϼ��Ƽ�   �   $'��&���;1��ꌽq�Ƚh�n� �P79�SlJ��uR��P��0E�T�1��������4���Dm��M�����M�<Z�0=`m{=���=d�=\��=t��=�(�=��=���=߷�=m�={��=�c�=�H=��=$�< �1;@]Y����4�6���q��𒽞���.*�������_�����sU��_�|����Ǽ��N�P6�� ��   �   h�C< <Q:Є����-
��g��10�XJ
��(���"�D\#��V�N��2���`�ʽ����NS�8�p9ƻ��m<&=��L=bȃ=%��=�&�=Ƚ�=@U�=�̻=}N�=<[�=eʌ=
{e=(+=8=�<�><��F� p��pD��)�\�R��v������y��J��@2������ �c�l�1��V�X�r��,��0�<Ѐ�<(�<�   �   ��=���<8�.<�A���+뼦fP� �����t^ؽP=�-�8p�lZ޽��ƽɉ���D����I����Jg���H;|4�<�H=b�G=ʦw=G��=	_�=E*�=���=�ˌ=�sr=V�>=<�=hk}<@Ň��}��������/�j W���s�K���뇽�������u�POY��3����D���R��Y<0s�<0L�<l�=��=�   �   �b=^�C=�=hT�<�_T;@��~N���Q�ǅ��(��;=�����T��/��Β�NH����T���#�(&ۼ(wO����:���<���<\�+=�GQ=Vdh=>�n=`�b=��C=��=(H�< �S;���W�(�Q��˅��-���A������W���1��В��H���T���#��ۼ gO��, ;t �<��<�+=*LQ=�hh=��n=�   �   ���=�͌=�xr=��>=X�=��}<@׆�n���x��D�/�\W���s��H��	ꇽ� ��?����u��RY�B�3����$�� ��xC<�h�<TB�<��=�=��=���<8�.<0v���:�,oP����A����cؽ�B�[2��t�^޽��ƽ&���$F����I�8���Bg� �H;8;�<�L=F�G=��w=; �=�`�=8,�=�   �   fλ=`P�=N]�=�̌=0�e=�-+=XI�<x�>< �F�$d���9�)�H�R��v� ����z���K��r4��@����c���1��b�x�r��ܽ���<8w�<��< �C<��O:�ۄ�Z��	���k��45�M
�{+���"�+_#��Y����.���m�ʽз���PS��缐5ƻ��m<d(=>�L=�Ƀ=���=\(�=f��=�V�=�   �   �=4��=���=�n�=���==f�=��H=n�=��< �1;8NY�P��6�L�q�L�ﮧ�$,��7���gb������X����_�\���ȼ��N��[���卻 6'� 0��LA1�#�Ƚ@j�� �:9�FoJ��xR��P��3E��1����q��>7��hHm��Q� ��dN�<��0=o{=���=��=���=���=:*�=�   �   ���=T�=(&�=J�=��=3��=��=D�P=
(=HJ�<@�� δ���,�}�3�����½\uٽBj�!���ؽ.���F�����J#>�z���м@�Ƽ���j�<�A.���ɽ���6*�8uK�h�f���y�ŀ�t�}��2n�J-U�A�4��P��Խ䈽Z���)��l��<ZL=���=���=�&�=Pz�=x'�=Ph�=�   �   &>�=��=��=0��=F��=�=�@�=�x:=�Y�<Ԑ;�Ę���.�Z���m���O޽F����G�	�ڹ���ŋϽꨪ�;ӆ��S��l/��*���I�]:���L��a���*%�E�L���q������!������'���ԉ��v��;P�>�%����̹���2� ��,9�<��\=�/�=Ao�=���=���=�*�=C� >�   �   �D>��>n�>"-�=xr�=���=P�=��=T�W=`�=�<����$�5�h�����ǽ<����/��m�j��4�
�<��W̽b��Q���($g�-b����l߽��"=���g�'쇾�C���������ꀣ��똾6P���f�RU7����O���b-�����P4�<*f=.Y�=�=�=���=O�=��>�T>�   �   e�
>{z	>��>�D�=Z�=l��=u8�=p�=�h=�5=�#<(ʌ���<��(���lӽ��N��N#��i'���"�����U�&������43��L��澂��o���b��{��R#!��}L�qcy�
������t����������X���%���&/u���B��A��N����;�����4��<d�j=�2�=�,�=d6�=RQ�=ĵ>��	>�   �   �>sp>�>���=V��=r��=|��=�z�=�e�=�^=T�=��<��(;�	{�b~�T?� m��Є��t��6���X�r��&T��M7�"�&�0�-���V�'蔽�ֽDE��+S�"l��r����ԾX?����AE�%L��F��~������1ӾX����4����>����6�t��&�d,�<�R�=�H�= 2�=0��=�>�h>�   �   D�>F�>��>���=��=���=�y�=aE�=�Y�=ڬU=��=>�<��:`�������;�(�g�m+����������h�Z�I�� -�ȵ�^i#�8mK�����G�Ͻ&����M�p3���F��`оGE�r���o�m��x������Ͼ�?��"v��<g:�h��ʵl�����<��=��=,F�=��=��>�V>�   �   ��>�4>
��=b�=@0�=��=@®=�S�=2�s=��8=���<x�h<����6�����*�3�ƬX���m��Oq���d��UK��6,����hg���$��+�\y�Rp��4$��]>��}��,���þ=��	��#7��	��Y��r��O��þ�N��Zu�r.���۽��U��ڸ��x=�(�=�m�="O�=�o�=�C�=�>�   �   V��=̊�=���=�Q�=d��=X:�=!��=qs=\z==�"=�ڛ<PϬ;XP�tQ��(���)���C�ĸO�N=L�$�:����4�� Wü����|<���f�@��1���l轿4&��`��������]`̾����S���z������;n���J����\�#9�}	½�4��`e���=�,�=.O�=X��=���=H��=޹�=�   �   ��=.��=�
�=��=ڪ�=��=SX=r"=���<x�f<�;�b���4_⼪���
$�X/��.�
� ��A��:мdZ���*�0����=ƻ��[��Z]�����F|�P�;���s�A3������N�ľƊҾ��׾6�Ӿ�Ǿ=��˚���
z�<?�*�����Z����;*=r=I��=*��=�r�=��=�"�=�   �   8�=6��=��=�ʏ=��f=*=�p�<��K<����	D��r��Hy�D�� ���e(���(�D� �6��8��X��(5����P�;H�0< B2<���;���hr��xw��Rɽ�����B��s�����F��	h��B��g]�����1|���?����P�����ܽ�肽H�˼п<b�=d�u=��=[F�=���=��=���=�   �   �۫=Aϗ=�%z=5:=��<@F)<0��t-���j�6�>��\�\�k��-o���g�~ W�ȵ>�\�����������[
�`>;��\<�^�<M�<���<�;�<@lT<�5��<6���Y��|�̽�q���8�}^��u}��K��w퍾�;���|���!o�Z�M�A'�T��􀯽�5K�w���<<P�= Ld=��=��=n�= �=�-�=�   �   P;�=�^U=t�=0�~<P�Ļ���v�G�����D��Yܹ��ý%!½-��6Ҧ��鏽Zrj��i0�����Z� )�:Xhy<��<C=��3=N==�1=z=���<@Δ��W��In����������o9�D`K�LxT���S�O\I���6��"��g�6�Ž�������wE�آ;<��=�H=��=��=帝=�=��=�   �   �2=�j�<g�;𾝼��<��╽��ɽ�[����
�4�.��;�4G���齲z½�f���EV�B��0�ذ<$ �<��!=f�P=�q=��=N7{=�ka= 2=<{�<���;ب��z�<��ە�3�ɽ*T����
�b��������D���齫w½e���CV��A�� 0���<�<�!=Z�P=&q=��=�1{=�ea=�   �   ��< ��l�Vn�����������9��dK��|T�ήS��_I���6�B%��i���Ž��������uE�(�;<
�=�H=�=��=��=��=��=p>�=�eU=ң=h�~<@_Ļ4�伴�G�F��>���չ��	ý�½�(���Φ�Q珽�oj�i0�t�缈�Z� Ȯ:�Yy<���<�>=��3=�==�1=Zs=�   �   `v��`I��t_���̽@u�.�8���^��z}�&N���>���~��%o��M�C'�W������V7K�|w��؜<<�=rNd=o�=K�=J�=�=�/�=>ޫ=Zҗ=-z==:=��<�m)<�L�����_��>���[�V�k�d'o�6�g��W���>�ҏ�T���l���Hj
���=;P�\<U�<�B�<���<@/�<HPT<�   �   ������w�<Xɽ���b�B�:�s����I��~j���D���_������}��BA����P�<���ܽ�邽h�˼��<��=\�u=C��=�G�=@��=f�=� �=>:�=Ď�=n�=�͏=�f=�*=T��<X�K<���h�C��d��|m�����:d(���(��� ������8���-5��z����;p�0<�+2<�V�;����   �   `b]�<������;���s�O5��������ľ�Ҿ;�׾I�Ӿ�Ǿ�������z��?�
 ��������;"+=
=F��=D �=�s�=|��=v$�=p�=$��=�=7�=���=�
�=^YX=�"=���<H�f<�R;�R����[�0���$�(/�:.�n� ��E�,CмXc��`=������gƻ��[�8#��   �   >5��!q�67&���`�L⏾ф��Pb̾�����T��K|�G���;n���	����\��9�
½4��Ae���=�-�=�O�=2��=���=Z��=��=���=P��=N��=�S�=j��=�<�=`��=�us=�~==�&=��<��;�I��O��d���)���C�X�O�z@L���:����(��<_ü(���E���p�@��   �   5s���%��_>�L�}�.��r�þ��⾛
���7�?	�)Z��s��"�hþO���u�Pr.���۽
�U��Ӹ��y=�)�=�n�=�O�=zp�=�D�=j>�>]5>4��=Pc�=�1�=���=�î=iU�=֫s=��8=���<8�h<@��|6��t��N�3�~�X���m�Rq�L�d��XK��9,�̞�Dn��X(��+�>y��   �   _�Ͻg��O�M�D4���G��aо?F����p�xm��x�L������Ͼ�?��v���f:����V�l����<���=l�=�F�=t��=�>W>��>��>��>H��=���=���=�z�=F�=bZ�=�U=��=�>�<�
�:��������;�P�g�,��Q��_��^�h�8�I��"-����k#�,pK�t����   �   M�ֽ�E�,S��l������Ծ�?��=��TE�'L��F�|~�<���:1Ӿ챬�64���>�U��Ȱt��&��/�<dS�=,I�=r2�=���=+�>�h>:�>�p>�>���=z��=���=���=�z�=�e�=��^=&�=h�< �(;p{��~��?��m�ф�"u��l�����r�|'T��N7� �&�\�-���V�%锽�   �   �ϽG����M�r3���F���_о�D�:��Wo��l�>x�������Ͼ�>��Hu���e:����b�l�(��@�<U��=��=G�=���=2�>W>��>��>��>l��=���=���=�z�=XF�=�Z�=̮U=��=�A�<�A�:���,����;�p�g��*��������T�h�L�I�" -�H�� i#�>mK�ٮ���   �   �o���#�]>�,�}�-,��P�þZ������6��	��X�Iq����PþJM���u��o.���۽Z�U�౸��|=�*�=Yo�=pP�=�p�=E�=�>6�>v5>d��=�c�=�1�=���=Į=�U�=:�s=��8=��<��h<�m꺼.�� ��R�3��X���m�<Lq�X�d��RK�>4,�h���c��#�$+�y��   �   90��)k轜3&���`��ߏ�ށ���^̾���L��#Q���x�����;����� ����\��6��½:4� �c��=)/�=Q�=��=l��=���=h��=���=���=���=T�=ª�=�<�=븓=�vs=t�==)=��<��;�7�,E��0���)�&�C�l�O�J8L�p�:�x���	��0Pü`����6��<a��@��   �   RV]�����z�_�;�x�s��1������Y�ľ��Ҿ��׾ӺӾ}Ǿ�
������z��?�(��������pG�;\0=�
=���=@�=�t�=���=�$�=��=z��=d�=��=��=�=�ZX=z"=4��<�	g< �;�@�X���N����H$�*�.��.��� ��;��/м�P���� t���ƻ�[�<��   �   $h��rw��NɽF��ΡB���s����rD���e���?���Z�����y���=��c�P�����ܽ�₽��˼��<r�=��u=ʈ�=�H�=��=��=X�=�:�=��=��=WΏ=ʞf=�*=$��<��K< 
���C��\���c�ܐ����:\(���(�ܿ �L������ ��@5�@2�`@�;��0<�S2<p��;`���   �   ���()���U����̽�n���8�$y^�Nq}�RI���ꍾI9��;z���o���M��<'��L��Bz���)K��b��h�<<�=�Rd=��=q�=�=��=b0�=�ޫ=�җ=�-z=�=:=��<�q)<@A�4���]���>���[�x�k�r!o�,�g��W���>���l��������>
��m>;X�\<�i�<W�<8��<E�<8�T<�   �   ෡<�����G�R@n�����Y
�����(�8��[K�lsT�ĥS�cWI�&�6�P��c���Žp�������ME���;<��=L�H= �=��=λ�=�=E�=�>�=�fU=��=(�~<�XĻ��b�G�f ���<���Թ��ý�½�%���˦�x㏽Rgj��_0�h���Z�@�: �y<���<vH=��3=&==�1==�   �   |2=��<�;������<��Օ�+�ɽZL��j�
�����"��)@�1���o½�]��
7V��*����/���<x*�<v�!=*�P=�q=�=Z8{=�la=�2=x|�<���;������<�nە���ɽeS��'�
���������NC����6t½ a��T;V�|/��(�/��<$-�<z�!=��P=tq=J�=�;{=�pa=�   �   �@�=�kU=��=�<�Ļ`��F�G�`����6��ι��ý�½� ��jǦ�3����bj��\0�X��0�Z� �:Pzy<���<pE=��3=�==�1=�z=���< ����V�:In�I������l��9��_K��wT��S�q[I���6��!�.f�ֵŽb������@VE���;<
�=z�H=�=��=2��=��=�=�   �   |�=�ԗ=�2z=D:='�<�)<���p ��HS���>���[���k��o��g��W���>��������h����G
� @>;��\<�b�<�O�<���<=�<�nT<p1��05���Y��=�̽_q�ը8��|^�zu}��K��A퍾�;��t|��� o�O�M��?'�SQ���}���.K�i����<<��=*Sd=��=H�=/�=��=�1�=�   �   <�=ᐽ=��=�Џ=��f=�%*=���<�
L< ���C��M��pV�2�����HY(�R�(��� �T�����8���5� ��p$�;��0<E2<���;����q���ww�TRɽl��p�B�փs�����F���g��YB��5]��T���{��z?����P������ܽ�傽�˼��<>�=J�u=��=XI�=Π�=��=��=�   �   ��=ؽ�=
�=�
�=H��=��=4`X=P"= ��<� g< �;�-�p���HI�*���$���.�D.��� �x>�(6м,W��&����� 9ƻ��[��JZ]�p���2|�<�;���s�73������?�ľ��Ҿ�׾�Ӿ�Ǿ�������E
z�j?�>��������/�;�.=
=���=��=u�=���=�%�=�   �   ���=���=���=zU�=^��=�>�=库=&{s=��==-=,�<��;8-��A��N���)��C���O�j:L���:�(�����|Uü\����;���e�Z@��1���l轱4&�	�`���������V`̾��
��S��yz��侜�;;�����@�\�~8�½�4���d���=�.�=�P�=��=���=4��=���=�   �   h�>�5>��=`d�=�2�=���=ZŮ==W�=ޯs=V�8=���<(�h<�8꺘,��~��l�3�ƩX�8�m��Mq�$�d��TK�6,����f��b$�Z+�0y�?p��*$��]>��}��,����þ7��	�� 7��	��Y��r��8㾪þ�N��u��q.���۽��U�pʸ��z=�)�=�n�=@P�=�p�=.E�=�>�   �   ��>��>�>���=X��=H��=u{�=�F�=`[�="�U=(�=D�< `�:\�������;���g��*����:��&�h� �I�� -����8i#�mK�����@�Ͻ����M�m3���F��`оCE�p���o�m��x���x��Ͼ�?��v��
g:����̴l�ذ�4 �<���=T�=�F�=x��=%�>W>�   �   � >�~>���=�i�=`7�=���=BԺ=�=�k�=�b{=��Q=j#(=�R�<�4�<��^< U�;�X�: x�� N��y�� �� �޹�ԅ���]�>� ���w�)Fӽ�.%�Lfq�1���T�ھ���l$�.c<���O��>\���`��?\��O��(<�q#�����־����f	]�3��o���E��i=ȍ=�-�=�v�=dJ�=mu>�   �   [�>&!�=��=���=X�=���=�q�=�0�=���=�6l=�vC=Nk=���<lS�<��F<���; b�:��A�@��� �����: ܘ:@����<���Jl�̽>� �x�k�s���[־�-��� ���8���K��4X��w\�"=X�$�K���8��b ��(�I^Ҿ����X���¨x��⾻
�=h�=���=���=t��=�G >�   �   p��=Jv�= ��=��=�8�=��=��=��=��e=H�==�=tf�<�5�<([<`��;`GN; �: 
O���V:��@;�~�;Э�;��:;�Q��lԶ�v�J�A1��^��Z�]O���Ⱦ����b��>�.�R�@��yL�s�P�*�L���@�H�.�����R���*ƾ,����I���?]�@	׺�� =���=��=���=J��=lg�=�   �   :��=��=��=w�=D#�=U�=��l=
*>=�1=|��<�Ж<�+=<���; d�:@(�� ���!�� � ���R;@q�;H�/<[M<~0< �`;��>�z���o���E��]Y@�����灴��>f	��y� H/�P):�_>�Qg:���/������	�3侊J���{�� 4�"�ԽB�3��͖;�:.=ʑ=h��=���=P��=x�=�   �   ���=@W�=�֭= �=ʀo=��4=�>�<��< ��; (3�p����`�L���pq��H)m��::��d�@S��<�;y><���< [�<,Ǩ<�t<�R ;����0Y�IwȽ���7ce�N���)�ľ%���
�G'�[�"��r&�=Y#����S%������ƾ"���URd����kq���wD<�<=�ƒ=P��=&�=B_�=\0�=�   �   ���=n̝=�y�=~�<=8��<�%< �����`��@0�`�C�JMH�?�4f*�"��XѼ>�������}�;0�y< ��<�f�<�U =��<Lp�< �������}������5�	�z��塾k�ž�o��> �i�����m	�H�����ʾ0L���w����;��T����L㖼���<�LI=�ˑ=��=�_�=�,�=J+�=�   �   7]�=�U]=��=�T<��)���	�v�a�8���岽,)Ľ?�ɽ��ýt'���h��z
~�l�<�x�� �S�@�6;�;�<P��<�=n�+=��'=�	=|L�<�ū��oϢ�ޅ��2>��L{��ʛ������̾�{۾�!��cݾ]�о_���l��0��
�M��l�PU��f9�P�ƻ���<\�P=Ǎ=b�=�^�=�ɰ=ZҤ=�   �   ^�@=<��< Ւ:�p���k�0���2�������*J&���&�\� o�������ɽV]��HI��ϼ O[��#�<dh=2�4=+S=��Z=�&I=��= �< .�`�)��D���&�*�4�A�e�1;��&;��S���a������fo���ѐ��\y�$�K����^۽HM��(
� Ԍ;@��<��P=��=��=�ݛ=�2�=�:�=�   �   H��< ����K�� ���$�$ �F�>���[�ٷo�Z�x�*�v�Էi�
HS��5�,���Q�͙�~/���]��BA<�=ЦG=ħs=.,�=l�=��e=$�+=��<`J��*?�$����6��>��[��o���x���v��i��CS���5�U��wMཐʙ��	/�(�]��CA<�=ҤG=�s=U*�=�=2�e= �+=�   �   �z��)��K���*��4���e�>>��^>��\V��e������.r��SԐ��`y�a�K�7�b۽�O����`͌;,��<�P=��=M�=�ߛ=<5�=>�=��@=���<@7�:�V���k�����)������XE&�$�&�;�ik�����.�ɽ�Y���I��ϼ�A[��"�<�f=��4=�'S=j�Z=�!I=h�=p�<�   �   <��բ����z7>��Q{��͛���� ;G۾L%�FgݾZ�о�a���n���1����M��n��W���h9�p�ƻ ��<n�P=ȍ=��=�`�=�˰=դ=q`�=�]]=Ŀ=BT<��)�ƍ	���a�f���ݲ�g!Ľ�ɽ#�ý�!��d��<~�@�<����S���6;�9�<4��< �=��+=�'=�	=?�<����   �   ����4���5���z�P衾{�ž�r澂@ �2��p��#o	�Ā�'��ʾ�M���x����;��V��u���喼���<�MI=�̑=$��=ga�=�.�=v-�=>��=�ϝ=r}�=.�<=��<(=%<�(�4����(0��C�&CH�l?�6_*���8Ѽ:�� ����x�;��y<4��<t`�<R =���<e�<�m��D���   �   O|Ƚ���ge�������ľ��h 
��(��"��t&��Z#�1���&�����ƾH����Sd�����r��&��vD<��<=Rǒ=3��=Q�=�`�= 2�=��=�Y�=�٭=_�=^�o=B�4=�P�<�	�<`?�; �2��x���`��򁼌g���m��1:��\⻀V���3�;�q><���<�T�<���<0�t<@��:�)���8Y��   �   iJ��1\@�r���򃴾[侊g	�.{��I/��*:��>��h:���/����n�	�a�dK�� |��� 4��Խ��3� Ж;�;.=�ʑ=&��=���=r��=��=���=���=��=�y�=&�="X�=�l=�0>=<8=(��<�ܖ<0@=<���;���:���@����� �"�@�R; b�;��/<xOM<0p0< o`;��>�f�Js���   �   �_�<�Z��P����Ⱦٗ��k��U�.�l�@��zL�r�P��L���@��.����9S��!+ƾa,��4�I����&?]���ֺ� !=M��=v�=V��=(��=fh�=���=�w�=���=`��=�:�=��=���=<��=�e=8�==��=�l�<�:�<H/[<p��;�NN;��: �O���V:��@;Pn�;���;@�:;0l��hܶ�h�J�V4���   �   �� �5�k�|���� ־�.��� ���8�M�K�$5X�#x\��=X�u�K�3�8��b ��(�;^Ҿ�����X��(�x�`־���=�h�=���=X��=��=DH >��>�!�=���=���=Z�=���=�r�=�1�=���=�8l=�xC=�l=���<�T�<��F<���;�S�: �A��׊� �� �: ��:���X�<���TNl�n̽�   �   �/%�Tgq�Ơ����ھ3���$�mc<���O��>\���`��?\�µO��(<��p#�����־���f]�U�����2��k=�ȍ=P.�=w�=�J�=�u>� >�~>���=�i�=�7�=���=`Ժ=�=�k�=�b{=��Q=&#(=�Q�<�3�<��^<�P�;@H�: ����`����� �� %߹�݅�p�]� � �,�w��Gӽ�   �   �� ���k�����c־�-��� ���8�S�K�4X�w\��<X��K�P�8�'b ��'� ]Ҿ����HX���x�`ľ��=Hi�=���=���=F��=VH >Ɣ>"�=��=���=p�=��=�r�=�1�=ɥ�=29l=\yC=�m=���<hW�<0�F<���;���:�-A�@���  ��@/�: �:��� �<����LKl��̽�   �   �]�n�Z�O����Ⱦ<�������.���@��xL�z�P� �L���@�7�.����P��)ƾ�*����I����L9]��dֺ�!=g��=?�=��=���=�h�=���=�w�=���=���=�:�=��=��=���=γe=`�==�=$p�<�>�<�9[<���;��N; f	: �K� �W:��@;���;P��;��:;�H��lҶ���J��0���   �   9D��FX@���������� �re	��x�G/�(:� >��e:��/�m��^�	���}H���y��7�3�j�Խ��3����;@.=2̑=>��=���=��=8�= ��=8��=/�=�y�=J&�=jX�=ޗl=�1>=r9=<��<���<J=<p��;�;�: �~� m��{��  � �R;���;(�/<@fM<��0<��`;��>�<��Tn���   �   �tȽ��(ae�����}�ľ�
��%���"�^q&��W#�+���#����S�ƾУ��jNd����l��V���D<ҽ<=-ɒ=���==�=Za�=�2�=G�=Z�=ڭ=��=��o=��4=@R�<��<�J�;@z2��o�`�`��끼@_���m�x:� .�@����g�;h�><$��<�b�<�ͨ<��t<�� ;(�� -Y��   �   �z��
��5���z��㡾�ž�l�:= ��������k	��}�/���ʾdI��;u����;��M��U���Ж�P��<0SI=�Α=���=kb�=v/�=.�=���=�ϝ=�}�=��<=D�<@%<�!���j��*0���C�@H��?��Z*�����ѼX-���m�����;�z<���<�o�<�Y =���<�w�<�������   �   ���dˢ�J���/>��H{��ț����t�̾^x۾G�d`ݾԭо�[���i��<-��,�M��h�^N���Z9�0�ƻ��<>�P=ʍ=4�=�a�=r̰=�դ=�`�=2^]=p�=�DT<��)��	���a�Ȋ��Oܲ�f Ľ��ɽ��ý����a���}�b�<�<��gS��q7;�H�<T��<��=��+=��'=.	=�U�<P����   �   ���8�)��?��^#�L�4���e��8��-8���O��g^��R���l���ΐ��Vy�ڢK� ��V۽}F��L��@!�;���<��P=��=��=���=�5�=�>�=��@=��<�J�:�U�V�k�u��&)����F���D&���&����j�������ɽ"W���I�|	ϼ �Z��0�<&n=<�4=�/S=��Z=\+I=p�=� �<�   �   H�<����5�:�����>���[�8�o���x���v�ܬi��=S�1�5�����D�#Ù��.�`�]�hiA<>=��G=r�s=�-�=S�=B�e=�+=�<�E���>����������>���[���o�;�x�;�v�B�i��BS���5�8���J��Ǚ��/���]�^A<� =ΫG=8�s=N.�=��=��e=h�+=�   �   ��@=���<�K�:�A�d�k�y��-!�^���~�@&�֢&���df�I�����ɽNR��B�H��μ��Z�p4�<�n=��4=J.S=��Z=�(I=��=��< )�أ)��D��j&��4��e�;��;���R���a������"o���ѐ��[y�3�K���>\۽�J����p�;8��<��P=��=M�=��=a7�=q@�=�   �   �b�=�c]=@�= fT< r)�b�	�~�a������Բ��Ľ�ɽb�ýF��\����}���<�l�� YS���7;DJ�<��<��=$�+=p�'=L	=TN�<P�����0Ϣ�Å��2>��L{��ʛ����~�̾�{۾�!��cݾ-�о�^��pl���/��(�M��k�&S��~a9�@�ƻ��<��P=�ɍ=x�=Vb�=�Ͱ=$פ=�   �   V��=(ҝ=���=��<=<�<Pe%<`��0ڵ���� �/�ʩC��4H��?�R*������м�%�� [�� ��;Pz<���<�l�<X =��<Xr�< }��p��}������5���z��塾a�ž�o澺> �c�����sm	�6�c�龴ʾ�K��Uw��.�;��R��(��\ۖ�$��<QI=1Α=���=�b�=T0�=@/�=�   �   ��=�[�=8ܭ=="�= �o=�4=b�<��<���;`�1��L��``�݁��R����l��:� ⻀c���j�;Ȋ><4��<�_�<pʨ<��t<@_ ;���x0Y�wȽ���&ce�G���!�ľ���
�D'�W�"��r&�6Y#����D%������ƾ㥛��Qd�"�� p������D<V�<=zȒ=S��=n�=�a�=�3�=�   �   ��=d��=��=�{�=|(�=�Z�=��l=�7>=�?=���<��<�`=<p��;@��: �}�`E��J�� @���R;P��;��/<�aM<��0<��`;P�>���zo���E��PY@�����ၴ���;f	��y�H/�M):�\>�Mg:�~�/������	��aJ��Z{����3�#�Խ�3�0��;h=.=cˑ=���=x��=@��=��=�   �   D��=tx�=���=���=<�=l�=���=���=ʷe=n�==�=�w�<|E�<hD[<��;��N;��	: �K� �W:��@;���;�;��:;PM���Ӷ�0�J�&1��^�رZ�YO���Ⱦ���a��>�.�Q�@��yL�s�P�(�L���@�B�.�}��wR���*ƾ�+����I����2>]���ֺV!=���=��=���=���=�h�=�   �   Δ>2"�=\��=4��=�=���=�s�=�2�=���=8;l=Z{C=|o=T��<dZ�<�F< ��;@��:�A�@��� ����/�:@�:�����<����|Jl�̽:� �t�k�r���X־�-��� ���8���K��4X��w\�"=X�"�K���8��b ��(�>^Ҿ�����X�Z��x�ݾ�п=oh�=j��=@��=��=NH >�   �   � �= 1�=bc�=@��=c5�=D��=d��=��=�Ʌ=�o=,�W=J�C=�h3=�A'=�=�=6�=:j=@=��=li=$��<�Dw<��߻�m&�Hp��0� ���z��õ�O���7!���G��zm��r��s������,��S��D����P���l�}�F����������g�{��Ze��� ;�A9=�=�=�=B��=��=�   �   hc�=�b�=�x�=|��=��=�h�=Y��=;��=2�u=�Z=�B=�!0="=Z=��=�Z=�:=re=�^=pB=��=���<��<@����v�fʰ��(���t��ٱ��K����/D�v*i��������\���?���a���������h�,SC���c��$`��5�b����b�[�`	`;VU<=�ۜ=|��=���=�_�=�   �   �=~��=��=�&�=jU�=͕�=֙|=[U=�N3=�=(�=��<T;�<���<���<���<�1�<Ԋ
=|�=�=��=�n=�[�< �9<����w���6�v�c�=������f�c^9���\�#|��n��wi���0��{�����!|��{\��8��	5�󠾵LS�`l�?���;&�D=���=�A�=��=� �=�   �   ���=�
�=e��=��=X ~=0�G=��=L��<�7�<��<�n�;��J;�8v;�<�;�0-<P �<��< ?�<
�	=�=
8=bv= 6�<��<�W��Ft~�����ȺH��Д��ξ�>{(�FI�Ff�}�_���}������f�}���f��ZI��{(�֐���˾|Ð�r�;�s�Ͻj9� �d<jQ=N@�=.��=~�=���=�   �   �=k�=���=�I=�=жp< ���бy�@�Ӽ�������� �����`�� P��: <pi�<��<HY=�c%=�a$=2�	=Կ�<@�Ż�k1��½�&���|�Fk��!b꾓��-0�o6J��^��6l�%�p�מl�u�_�AK��1�*��뾺 ����x�`3�䢦��D���L�<j _=���=�t�=H��=�c�=�   �   ��=�)f=��=��s<h��TC �FyV�(@��Lz��"�����]���ߝ��P��Z�B�����(I��]�; O�<�=��&=��4=��(= ��<�J<K���1�����VJ� ��(;¾�����*���<��EH�2|L�9�H�6�=���+�q��1���]�ľg�����K�Z���N�r������<�)k=�=�i�=Fu�=4��=�   �   �EH=�2�< �:D���6v�D������n��!� ���(�(�x���Z����g�����\A"��s�`��;���<��=E@=�>E=X;*=X��< Da9`|�gA��\���E_�}����þ���	����$�"�A{&��#��T����a��Ⱦ�����h�jl�=z����`��;Hy=ƿr=���=z�=苙=�w�=�   �   d�<��	���2���������c(���M��$l�]��h߄��E��حw���^��m>��o�!t彮����e&�Ȃ'��x<�o=�'D=T�\=��T=�Z*=�̳<�E��fe@��)Ž���t`�����?��ԾF��x���|�����15�پ����Dj���Bp��.��L㽮�s�Շ�X��<�a/=P�s=E��=��=\iu=�D5=�   �   hc3���K�"�ý;+�aM�bh�������7��s9��o{��؊��kȱ�Y����L2a��,����*��bo�@֏:p�<��>=�hl=|Dy=�@d=�r,=���<p73��K���ý&�e M��d��Ʃ���3��Z5��bw�������ı��U����-a���,���2'���j�@%�:��<Ψ>=zfl=Ay=�;d=Tl,=l��<�   �   �q@��1ŽY�Tz`�N���C��?Ծŭ����ċ�o���.9�پ�����l���Fp��.��P���s�ۇ����<�a/=�s=�=��=ou=RL5=d%�<0z	���2�ߵ������](�6�M�0l��Y���ۄ�<B��ԧw�7�^�i>�l�en�p����_&��t'��x<�o=F&D=��\=��T=DU*=0��<����   �   �G������J_�������þ-����	�a����"��}&�N�#��V�����d򾡩Ⱦ�����h��n�}��!���;>y=��r=ٳ�=>�=U��=�z�=�MH=�F�<��:���J&v�⥹�}������� ���(��(�����V�4��a�����:"��rs��
�;���<r�=PC@=�;E= 7*=|��< rY9����   �   ����jZJ��"��a>¾����/�̬*�(�<�PHH��~L���H�K�=�� ,��������N�ľ� ����K�����j�r�С�l��<�*k=�Ú=�j�=Hw�=ǲ�=��=�1f=D�=��s<����4 �$iV��7���q��w��돺��U��ٝ�PK��@�B�4����I�0w�;@R�<H�=��&=z�4=��(= ��<�2<[��+7���   �   4�&���|��m��=e�a� 00��8J�L�^�9l�`�p��l�Y�_��K�X1�D�������^�x�w4�$���<G���L�<D!_=u��=$v�=��=�e�=���=<n�=��=��I=�=��p<@��p~y�4�Ӽ���ʰ�Ц���� ݻ� `���O�HH <�m�<��<�X=2b%=�_$=ޗ	=ж�< ƻ|s1�߄½�   �   ϽH��Ҕ�7ξm��|(�I�.f�}�Y���l�������}��f��[I��|(�v����˾Đ�$�;�"�Ͻ�9���d<kQ=�@�=&��=E�=,�=���=N�=* �=P��=�~=L�G=��=t��<�I�<(<P��;�hK;@�v;�j�;�B-<��<T�<HA�<,�	=�=�6=t=�/�<��<�b��z{~�/����   �   �c�ف����侍��_9��\��|�uo��0j���1���{�������!|�k|\���8�h�r5�J��LS�Rl�f~?�`%�;J�D=G��=�B�=޽�=�!�=t�=��=
��=�(�=�W�=v��=��|=�`U=zT3=֪=��=��<�C�<���<\��<d��< 4�<4�
=R�=4�=�=�l=4V�< A�9�����z���8��   �   ��t��ڱ�FM���0D�f+i�T	��f��$]�� @��7b�������h�8SC���7���_����b�&����[�@$`;�V<=�ܜ=0��=N �=�`�=Jd�=�c�=z�=���=(�=?j�=ط�=���= �u=�Z=��B=�#0=�"=�[=��=:[=�:=Ze=^=�A=��=���<���<`���Nz��̰�L*��   �   ��z�?ĵ��O��08!�^�G�,{m��r���������/��E��(����P����l��F������������g��~�fWe��� ;�C9=��=h>�=Ƶ�=�=B!�=~1�=�c�=���=�5�=���=���=-��=�Ʌ=�o=�W=
�C=&h3=|A'==��=��=�i=�=6�=�h=��<x>w<�
�p&��q��.� ��   �   8�t��ٱ�L����/D�O*i�������t\��m?���a�������h�MRC��� ���^��Kb�����[� F`;VX<=.ݜ=���=� �=�`�=ld�=�c�=z�=ȇ�=8�=Nj�=규=���=v�u=Z=&�B=�$0=�	"=h\=��=V\=�;=�f=|_=C=P�=��<���<P����w�˰�%)��   �   �c���������]9��\�L
|�4n���h��T0��hz��G����|�bz\���8��	�3�|�'JS�Uh�x?��E�; �D=D��=LC�=\��="�=��=H��=.��=�(�=�W�=���=ڟ|=paU=U3=��=r�=��<hF�<���<��<���<�8�<��
=�=�=�=&p=x]�< d�9$���Cw��^6��   �   ιH�Д��ξ[�az(�/I��f��}������������z�}���f��XI�"z(�r��}�˾����d�;���Ͻ�1���d< oQ=aB�=��=��=��=���=��=^ �=���=~=��G=�=���<�K�<
<p��;��K;��v;@}�;XM-<��<��<0H�<އ	=�=�:=�x=�9�<��<�S��r~�����   �   l�&���|��i��T`�o��,0��4J�#�^��4l���p���l�6�_�K��1�\���	����k�x��/�����4��LZ�<&_=$��=Iw�=���=Pf�=��=�n�=��=P�I=R=��p<@����{y�h�Ӽ���R�����X���׻���_��xO��W <�u�<`�<�]=0g%= e$=��	=<Ś<��Ż:h1��}½�   �   _����SJ���9¾w���|���*���<��CH��yL���H�Ϟ=���+�S��l����ľ����R�K�G����r�x����<�/k=eŚ=@l�=$x�=d��=c�=t2f=��=��s<���4 ��hV�D7��q�����!����T���ם��I���B������I�@��;�[�<j�=<�&=t�4=v�(=��<�Y<LB��5/���   �   q=�����iB_�P���,�þ����	������"��x&���#�R�ʼ��]�X�Ⱦӥ��8�h�h�2s��t�A�;�=b�r=ǵ�=��=<��=K{�=�NH=4H�< !:����%v�����0��ȕ�L� ���(�f(����U����`��-	��|6"��`s��1�;���<
�=tI@=�BE=:?*=���< f9Jv��   �   `]@��$Ž2�Lp`�I���<��_ Ծ4�����/��r����0��پϛ���f���<p��.�zD��s� ������<Hi/=*�s=�Ċ=5�=�pu=�M5='�<�w	�r�2�����N���](��M�l��Y���ۄ�B��c�w���^�jh>�Ek��l�t���p[&��a'���x<du=8,D=��\=�U=_*=�ֳ<����   �   �3�\�K�Y�ý2"���L�b��|���!0��d1��@s��΂������R��d쉾�'a�E�,��	���@^� t�:`�<b�>=rml=�Gy=�Bd=tt,=���<x43���K�i�ý&�J M��d�������3��E5��Ew��Ԇ���ı��U���;-a��,��?%���f�@��:��<L�>=�ll=�Hy=�Dd=�w,=���<�   �   H3�<�V	��2�����+���
Y(���M��l�9V��t؄��>���w���^�
c>��f��d�a���.R&��F'�H�x<(x=�-D=��\=�U=�\*=�ϳ<P>���d@��)Žv�vt`�����?���Ծ9��g���p������5��پ�����i��Bp� .�K���s�͇�,��<tf/=�s=�Ċ=��=�su=�Q5=�   �   �SH=�U�< Y:d}�\v�����!{�Ȑ��� �,�(�� (����'Q�%��X�����,"��Cs��[�;̞�<�=,J@=�BE=�=*=���< Zb9�{�$A��>���E_�u���ٮþ����	�����"�:{&���#�zT����a�֦Ⱦ�����h��k��x��j�0�;t}=��r=���=
	�=Z��=}�=�   �   m�=�7f=
�=��s<���p' �HZV�j/���h��O������~L��YН�>C���~B������H�ǘ;dc�<��=t�&=��4=�(=��<@P<PI���1������VJ� �� ;¾����{�*���<��EH�/|L�4�H�/�=���+�`��	���+�ľ*���3�K�!�����r������<�-k=�Ě=|l�=�x�=ȴ�=�   �   ���=�p�=��="�I=�=�q< ����Ly�x�Ӽ�������� ���Ļ�H�_��
O� m <�}�<��<F_=�g%=e$=d�	=�<`�Ż�j1��½Ո&���|�>k��b꾐��-0�o6J��^��6l�&�p�՞l�q�_�;K��1����뾏 ��F�x��2�١��\@��R�<�#_=���=@w�=*��=Qg�=�   �   ���= �=V�=쳙=�~=|�G=��=X��<]�< .<@�; 
L;�@w;���;�d-<`�<$��<�M�<��	=�=6;=�x=9�<��<8V���s~�S�����H��Д��ξ�<{(�EI�Ff�}�`���~������e�}���f��ZI��{(�ʐ���˾XÐ� �;���Ͻ�7���d<ZlQ=�A�=���=&��=:�=�   �   <�=(��=X��=b*�=�Y�=���=��|=�fU=�Z3=J�=�=��<�P�<��<���<���<�=�<��
=@�=Э=��=jp=�]�< m�9P���dw���6�j�c�9������d�b^9���\�#|��n��xi���0��{�� ���!|��{\��8���4��򠾃LS��k��}?��'�;��D=s��=�B�=D��=\"�=�   �   ~d�=4d�=�z�=X��= �=@k�=���=
��=�u=�Z=��B=\'0=,"=�^=�=$^=t==�g=l`=�C=��=X��<��<Ј��jv�Nʰ��(���t��ٱ��K����/D�v*i��������\���?���a��������h�)SC���[��`���b�����[�@`; V<=_ܜ=��=@ �=�`�=�   �   X��=��=Lv�=Q�=4��=���==#�=.�q=�IW=��C=P8=N�3=�5=(==n�H=dW=�e=j�q=�dw=0$q=x@X=x4$=��<�G��y����)�n�m� ﵾ����)/���`��%��g΢�����&�ɿ��Կ�ؿ��ԿB�ɿ~h���l��i���5e_�R-��n���;��Ҍ\���� T#�ȃ�<<�c=&�=HA�=��=�   �   V�=X.�=_�=�h�=�^�=WÏ=Rhx=�V=�:=�	'= �=��=�+=�'=��6=H=�	Z=,]i=*�q=�Yn=�W=r&=���<�rg�����Fh����x��h�+�n�\�"�������u���^ƿ<ѿ��Կ�Bѿ�\ƿnT��R���\2��o[�5�)�j�������noW�!�彜��(I�<�e=���=`�=(��=�   �   i��=S$�=���=�R�=C��=h�W=�L)=$\=h �<쨜<���<�!�<(�<�V�<���<ZF=hZ6=lNO=��`=Dae=h�V=�|,=@�<0��c�����b~W�t���}j�,"���P�ƕ��Lʗ��O��{����ƿ�ʿ��ƿH���4]�����J����O�&� � E�=���H�-�ѽK�`�<�?j=:��=���=��=�   �   l�=�]�=��=L�]=t�=��<�< ���`�Y�dЗ�<���<����s>� mQ�з�;��<���<nt!=,B=(�T=�jR=nT4=��< 1���/���ӽ��=������׾<�hB>���j�t���L���G��\��� ��Iڶ�qL��9G�� ��,�j���=��2��վ뵐�bt1�����Dn��d��<\�o=�΢=V\�=�[�=�   �   0�=��s=:�*=p��< ���P���K)���j�����o���D���B����
q�L�7��U輘�0��\�;�<$=��8=ЊH=\;=��=x�#<�.޼N7������}��E��%���l�&���N��1u�L���WC������Z��d@�����m<���v��*O���&�k���ո���w�/D����h:'�
p=
�t=
�=d�=R�=�   �   ��P=��<p��;�꽼�FY�˕����޽�h�����u����r�����qѽ^����O�<�ʼ �`�D�<ʈ=��5=օ==< =42�<+�~a�����QK�6ᘾ��Ծ%���r.�P���m��΂��t���4��=Ɗ�^��eUo�9vQ�b�/�y��{5־�4��B�I�RP��S@� �*;�=�^u=��=u�=&��=�   �   �2�<�ӻXX)�2Z��i���<�$�z�I��]g�S{�B܁����|p��W�{"6����,;ӽk1��R��`�&����<�=�8=�3=NV=�#
<ؿ�0R���=���l��]����߾^�|D)��B�ȇV���c��Bh��=d�J�W��6D��-+����r�㾎r��xNq���������м�x<~:/=~�o=R9�=�|p=�7=�   �   hA��S�rʽ���X�R�^Ƅ�~����[��f���ٱþ!}���E���2��S���c��m-�������L����C;���<��)=j@=�4+=(��< �8���3�Iɽ�b)�X4z�(����ؾo����Jc(��3�Z7��3�|�)���A���=޾�V�� ?��ý2��ؽ��I�p��Li�<��==\Jb=[=�)=L�<�   �   �hV���ֽ�*�3q��V��'\��'��w���{T��	��3�a��œ澦UǾn!�����9����#��L9���{F<�O=x�C=�YK=��&=�]�<��'��ZV���ֽm�*�jq��R���W��������Q�.�	�1����o���QǾZ����1�9����x	��<0��ȄF<P=ڨC="VK=b�&=N�<8�'��   �   $ɽ�g)��:z���[پ�q���Kf(��3�h	7���3�.�)���Q��ZA޾0Y��A����2�$�ؽ�I�����g�<��==$Mb=�[=��)=��<��@��qS��ʽ����R���>|��W���{��3�þ�x���A��M/��(��եc��i-�`��f�����@~;���<��)=4@=�0+=���< �9�p�3��   �   B�,�l�Ta���߾��AG)���B���V���c��Eh��@d��W�	9D��/+�}��<�㾪t���Qq����������мx<0;/=��o=F;�=<�p=d�7=�F�<аһ�H)��P��~�����$���I��Vg��K{�}؁����Pup��W�S6�p��h4ӽF,����� k&�4��<��=�8=�|3=�Q=H
<��鼞X���   �   SVK�䘾4�ԾK��Uu.��P���m�BЂ��v���6���Ǌ�w_���Wo�JxQ��/����7־F6��;�I��R罔V@���*;J=�`u=���=^w�=A��=��P=H��<`#�;tͽ�n5Y�����޽c��}�p�"��@����iѽ������O�P�ʼ p_�|�<��=�5=\�==, =d(�<�G�އa�2���   �   J�}�\H��N ��&��N��4u������D��K�������A��W����=���v�O,O��&�$���Oָ�^x�.E�����='��p=��t=V�=<�=��=^�=��s=��*=ƭ<���D3���;)���j�ݙ������𰘽������p�h�7��A輀�0�P��;8�<�=��8=`�H=�;=R�=h#<�<޼&<�� ��   �   ���G�׾��ED>���j������ ���������W��g۶�pM��H��� ��K�j���=��3��վq����t1�8���Pn����<��o=�Ϣ=�]�=h]�=��=�`�=�=~�]=��=�/�<�!<����HcY������������XM>�@�P����;@�<��<w!=�B=^�T=�iR=lR4=���< �����/�K�ӽ��=��   �   &����l�l-"�B�P�����9˗��P��
|����ƿ��ʿ��ƿ�����]��|���dJ��c�O�o� �rE�`����H���ѽ,J���<RAj=%��=���=^�=��=V&�="��=UU�=Z=B�W=�S)=�c=�<D��<<��</�<�<a�< ��<�I=�\6=�OO=�`=�`e=Z�V=�z,=H�< "��c�q�����W��   �   N	��z��[�+���\�����(����u��h_ƿ�<ѿS տ?Cѿ(]ƿ�T��m���d2���n[��)�"���g����nW�
�彔���L�<��e=S��=�`�=��=W�=�/�=��=$j�=�`�=%ŏ=lx=bV=�:=�'=��=��=�.=*�'=t�6=VH=d
Z=|]i=�q=.Yn=��W=Dp&=x��<��g�����Mh��   �   �ﵾ��*/�=�`�&���΢�Ӛ��Q�ɿ�Կ�ؿ��Կ�ɿKh��Yl��$����d_��-��m��/;����\�����P#����<$�c=��=�A�=���=���=��=�v�=lQ�=���=ꃛ=s#�=��q=JW=��C=.8=�3=��5=�==��H=�W=V�e=��q=�cw=H#q=J?X=�2$=4��<�L������*���m��   �   P���x����+�y�\����s����t���^ƿ�;ѿj�ԿZBѿP\ƿ�S�������1���m[�J�)�݄��t���vmW���ړ��P�<صe=Ƅ�=@a�=J��=>W�=�/�=��=0j�=�`�=0ŏ=6lx=�V=�:=�'=��=<�=(/=��'=�6=H=>Z=b^i=�q=DZn=<�W=�q&=��< wg�o�����h��   �   B���!j��+"�G�P�r����ɗ�cO��hz���ƿʿ��ƿW���C\��'���>I��u�O�� �C뾑��X�H�/�ѽ�D�'�<�Cj=���=6��=��=Z��=�&�=C��=tU�=v=v�W=&T)= d=��<<��<\��<�0�<��<<c�<p��<K=4^6=�QO=��`=ce=ƥV=d},=H�<8��c�W���2~W��   �   :����׾���A>���j���r���J ��A������ٶ�2K��F������j��=�p1�mվ𳐾Rq1������_�� ��<>�o=Ѣ=�^�=�]�=*�=a�=@�=��]=$�=D0�<�"<����`aY�ܶ��\����~��xH>� �P� ��;�<��<py!=,B=b�T=FmR=\V4=@��< n��L�/���ӽս=��   �   �}�CD��U���:�&�/�N�0u�6���B��s�������>������;��Pv�w(O���&�����RҸ�g�w��@�L����'��v=��t=��=4�=i�=��=J�s=>�*=�ƭ< ���2��l;)�F�j�����e���}���������p���7��=輈�0����;�#�<�=�8=f�H=P;=>�=�#<�(޼b5��v��   �   �OK��ߘ���Ծ���q.��P�9�m�L͂�zs��h3���Ċ��\��`Ro�osQ��/�T���1־�1��ĘI�XI��H@�@I+; =Veu=>��=mx�=���=��P=���<�'�;�̽�5Y�የ���޽�b��}��o����������3hѽ�����O�ܤʼ �^�D��<b�=z�5=��==�! =9�<x�ya�6���   �   F;�N�l��[����߾��RB)�1}B���V���c�g?h��:d��W��3D��*+�F��?��o���Hq�z��$���8�мX7x<B/=t�o=�<�=\�p=̈7=�H�<`�һDH)��P��L����$���I�kVg��K{�g؁�z��up�tW��6���23ӽ�*������3&�왪<0�=J�8=��3=JZ=�5
<��鼃N���   �   Fɽ�_)��/z�W���U�ؾ�l�C���`(��3�O7���3�z�)������\9޾�R���;����2���ؽ��I�`����z�<��==�Qb=�![=��)=P�<��@�qS��ʽБ���R�|�4|�� W���{���þ�x��sA��!/�����Y�c��h-������h��� �;���<�*=�@=�8+=���<@�8��3��   �   (QV�~�ֽZ�*�Bq��O���S�����:���O�o�	�R.�!��X��LMǾG����h�9���������ЬF<�X=��C=�]K=��&=|a�<�'��YV�v�ֽR�*�Wq��R���W��������Q�'�	�1�i��L���QǾ%�������9�=����|)����F<�T=ЮC=�]K=��&=i�<��'��   �   X�@��fS��ʽi���R�A���|x���R��8w����þ�s���<���*��7����c��c-�^��)�������/;\��<�*=�	@=d8+=��<��8���3��ɽ�b)�B4z�����ؾo����Fc(��3�T7��3�r�)�t�/���=޾JV���>��5�2�͛ؽ��I��찻�q�<�==BQb=,#[=�)=��<�   �   �U�<0eһ�<)�bI��e�����$�r�I��Og��D{��ԁ����mp��W��6�����*ӽ�#������%����<�=t�8=>�3=lY=�+
<4���Q���=���l��]����߾Y�yD)��B�ƇV���c��Bh��=d�E�W�~6D��-+����H��]r��Nq�`��ڐ��0�м@"x<�>/=b�o=>=�=̆p=�7=�   �   ��P=���<�q�;�����&Y�����<�޽�]�!x�j�!��g��l���^ѽ�읽��O�8�ʼ �\���<��=b�5=,�==�! =D7�<�$��|a�5���QK�-ᘾ��Ծ#���r.�P���m��΂��t���4��=Ɗ�^��`Uo�/vQ�V�/�i��W5־�4��ڜI�`O罄Q@�`�*;�=�cu=N��=Cy�=���=�   �   ��=��s=>�*=�ح< ������(-)���j�F���ф��𧘽�~��<�p��7�&� z0����;�0�<h=h�8=��H=r;=z�=�#<`,޼�6�����}��E�����j�&���N��1u�K���XC������[��d@�����m<���v��*O���&�R����Ը�s�w��C������1'��r=Ќt=��=��=���=�   �   q�=�b�=��=�]=��=�A�<�J<�B���2Y�̞��pr���g��@>��4P��?�;p��<��<~!=�B=΅T=�nR=VW4=��< ���4�/���ӽ��=������׾:�eB>���j�t���L���I��]��� ��Iڶ�sL��9G�� ��'�j���=��2��վе�� t1���� k�����<"�o=�Т=�^�=�^�=�   �   
��=�'�=Ï�=^W�=�Ą=��W=nZ)=k=��<pȜ<�Ċ<D?�<���<�o�<|�<�O=b6=�TO=j�`=�de=�V=h~,=��<��Dc�\���V~W�n���zj�,"���P�ƕ��Lʗ��O��{����ƿ�ʿ��ƿG���3]�����J����O�"� �E�,��ŕH���ѽ�I� �<�Aj=j��=��=�=�   �   XW�=�/�=[�=�j�=�a�=kƏ=ox=�V=��:=�'=��=��=�2=��'=�6=�H=pZ=D`i=��q=�[n=`�W=�r&=���<0qg����	�?h����x��g�+�l�\�"�������u���^ƿ<ѿ��Կ�Bѿ�\ƿmT��R���[2��o[�2�)�c�������ZoW������hJ�<Ƴe=��=�`�=*��=�   �    d�=6��=�ڶ=�ڣ=x[�=6(q=��H=F<'=�z=: =���<\N=O=��*=B_F=��c=�t=tK�=�͎=�߉=~�n=�$=�7<�O���ֽZ.L�^���v���'0�4�j�C��������ԿOh��#�l9
�$���8
�����xGԿ	�^A���h�%�-�����fР��=�5��pϒ���=M�=��=4w�=�   �   ��=P{�=�í=�ژ=5v�=V�S="a(="?=���<�K�<���<���<��<�2=D�-=qO=�o=��=�e�=
,�=D�l=�'%=`�.<����н�G�`d���p����,�&�f�P���w���Iѿh�T� �`��Z
�L���� ��3���п��������%zd��w*�4��m��F89��L���8���=���=Ԭ=���=�   �   �Y�=I�=��=ءn=*4=<��<\L�<p!�;��ú0��� ��� 9����;x]<H��<h�=
==j�a="�y=6�}=�te=��'=@cb<<��[c���t8�ߘ����~#��3Z�-������+�ƿR���J���E����@Y��z�������ƿz@���l���X��3!�<e�t����+��5��H�<���=���=�C�=�8�=�   �   `�=tف=�?E=�c�< 0<��PKѼ0"���I���\�l�Y��A����l,��pp��H<4P�<\�=�GJ=L�_=��W=^*=P��<����6杽N�!��~���.оv���F��U~�Ӑ��^���f�ο,��K��R>�i/�
�cϿB�������G�}���E����i�̾�A�����ȃ��m����=p�~=���=�g�=�   �   B$]=D?=�Mk<`�7��U�iF���	���dܽ����$E��W��v�=�ʽ窠�f�`������ѻ�u<̯=�1=&�@=��(=H��<0��wo�����g��}��m� �"H.�!	`�k���O��������ȿ|�ӿ�׿1$Կ�`ɿ�b��ԥ�������H`�/.��9 �Jo����a�s����E� ��;�h=��q=+��=�Q�=�   �   ���<��A:� �湉��׽FT��\3�/�N�?�`�4Xh��^d��U�~]=��1�f���M���I�4����<t?�<n|=�� =8��<�%_;����7ɽ69�uC����־���Z�=�9j�����{���m��<�����������0���`��xc��Λk���>�	�	�־蜒��6����^���rV<�z%=�[=�B`=L�9=�   �   �����9�u��I��D�� y����/��_x���O�����:���Ø��g���OR�\�O|׽�zx�أ�����;Զ�<��=H�=p!u<t����ꆽj$	���c�-�Yj�����`?�.�c��避a���㖿�㙿�W��t��M삿Ϸe��EA��n�������S�e��	�+��8[S�� �<��$=x�:=U=pI�<�   �   �LP���ѽq'��?l�zb��۽�ͼݾ�;��r��H!����^���&⾿8þ�]����x�ܰ3��6꽾�~��Ĩ�@$<���<�=̽�< �6;�,��`���]#�
g}��y��A�� w�43�.�M��yb�)p�u���p�d�D�O�/g5�C���.��(�� Ɓ� &(��ܻ��� �X;@��<��=�T=�ѕ<�)��   �   6н�!.��9��3𭾽�ݾ�2�����+���6���:��t7��U-��>�K����6-��E6��N7��m��8[���9��D�<�=t=��<@ϻ�@�O-н .��5���뭾��ݾ�/���H�+��6�s�:�Sq7�zR-�"<�׮�� ��)���3��^J7��h�:2[���9��F�<��=�=( �<�[ϻ�'@��   �   �b#��m}��}��>��z��3�҄M�o}b�p��u���p��d�a�O��i5����_2�+��ȁ��((�J໽� �X;���<��=�Y=��<H�)��=P�xѽd�&�z8l�^��ֽ�I�ݾ�5��h��A����Y���!⾌4þ/Z���x���3��0���~�����X/<���<��=ȴ�< '6;,7�3h���   �   ��c������n뾮���c?���c��끿g���喿�噿�Y���u���킿��e��GA�ep�������2�e��	�R���bS�L�<�$=��:=�[=�[�<����9�Gk��C���D��y�9��i���os��
K������5������Yd��=JR���>u׽Hpx�����@��;���<\�=��=�u<����g���t(	��   �   HF��L�־	���=�B<j�ŉ��}���o��E����������|2���b���d����k�t�>�m
���־=����6���xb��hsV<�|%=��[=6H`=Ȥ9=h��< �D:���������ֽN��U3�ΰN���`��Ph�9Wd�D�U�VW=�V,�����)���I����X�<�E�<h}=�� =؛�<`�^;f��>ɽk#9��   �   a���8� �[J.��`�𓉿���q�����ȿ_�ӿ��׿�%ԿEbɿd��������`J`�O.��: �ap��
�a� ���P�E�Њ�;dj=ةq=R��=�T�=�+]=�H=0}k<�O7�ZE�=��v����Yܽ9����?�M��W� �ʽ����"�`�����@�лطu<��=�1=X�@=�(=D��<P.�|�o�����g��   �   T1о��F�X~�,���ؼ����οɪ�����?��0�M�w Ͽ&�������^�}�j�E� ���̾5B��H��ȃ��h��h�=��~=[��=�i�=>�=݁=�HE=�w�<D0<���h.Ѽ�"�8�I��}\�T�Y���A���p���&��� <�[�<^�=JJ=D�_=J�W=��)=4��<����?Ᵹ$�!������   �   ���#��5Z�%������T�ƿ���.L���F�@���Y��{��r��W�ƿ�@���l��G�X�4!�oe⾀�����+�H5��(�<�H�=� �=�D�=�:�=�[�=���=��=��n=�$4=t��<�^�<�o�;��º@Y���j�� ��0Ő;�"]<���<��=d==��a=\�y=n�}=te=��'=�Ub<D���f��8w8������   �   Nr����,�\�f�����5����Iѿ�h쿴� ����hZ
������ �4�
�п��������zd�pw*�4�{m���79��K��\4��֤=���=!լ=���=D��=�|�=jŭ=�ܘ=@x�=��S=�e(=D=���<(U�<���<���< &�<�5=��-=�rO=,o=O�=�e�=�+�=�l=�%%=��.<ج��н�!G��e���   �   �w���(0���j�nC��,µ��Կ�h��#�|9
�&���8
�����'GԿ��A��_�h���-������Ϡ���=�3��Tɒ���=3�=@�=�w�=�d�=���=j۶=ۣ=�[�=�(q=��H=�<'={=F =x��<N=�N=Z�*=�^F=��c=�s=K�=m͎= ߉=�n=�$=X.<�R���ֽ�/L�7���   �   	q����,�I�f�W���m����Hѿ�g�(� �$���Y
����<� �
3�+�п���꽑��xd��v*��2�l��V69�J���/��v�=9��=~լ=��=n��=�|�=xŭ=�ܘ=Jx�=��S=�e(=$D=���<xU�<��<<��<�&�<6=0�-=lsO=�o=��=
f�=B,�=8�l=,'%=X�.<.���н4 G��d���   �   ���E#��3Z����7�����ƿ���J��uE�$���X�uy����࿬�ƿn?���k��J�X��2!�c�Η����+��1���<�\�=�=�E�=;�=�[�=쁧=��=��n=�$4=���<$_�<Pq�;��º�V���h�� ���ɐ;`%]<P��<��=r==��a=Ьy=$�}=.ve=l�'=hdb<��\c���t8�ߘ��   �   �-о���:�F��T~����w���S�ο������<��-�w��Ͽ�󶿦�����}���E������̾�?���
�ă�06����=��~=L��=tj�=��=E݁=�HE=tx�<�D0<(��.Ѽ�"��I��}\�؎Y�^�A�J����� �� &<p^�<�=
LJ=��_=:�W=P*=p��<����K坽��!�<~���   �   g|���� ��F.��`�u���&��F����ȿȿӿ�׿U"Կ�^ɿ�`��-���;FF`��.�'8 ��l��m�a����F�E�pǈ;�o=P�q=t��=�U�=�,]=�I=�~k<�N7�E��<��\����Yܽ���h?��L��뽱�ʽv�����`�������л��u<�=��1=��@=��(=���<0��to����N�g��   �   B����־a����=��6j������y���k��]��Ò�������.��_���a����k���>���d�־���s6�9꾽LJ����V<z�%=l�[=�J`=j�9=���<��D:���b�����ֽ�M��U3���N���`�zPh�Wd��U�W=�,�ϐ��Z��,�I��󑼀�<�K�<L�=�� =P��<@`_;j��5ɽ)9��   �   [�c�奄ug�!��2^?�l�c�Z聿����ᖿ�ᙿ�U��r��bꂿG�e��BA��k�������ʈe��	������1S�@�<��$=��:=:^=h_�<���l�9�k��	C��D��y�4��c���hs���J������5������6d���IR�b�Ut׽ nx�|���P�;���<��=|�=�2u<D{��C熽&"	��   �   �Z#��b}��v������t��3�~M�$vb�sp�$u���p�8d���O��c5�S���)�$����� (��Ի�L�`�Y;4��<Z�=�]=t�<{)��<P��wѽF�&�g8l�^�� ֽ�D�ݾ�5��d��;���yY���!�k4þZ����x� �3��/꽎�~�г��x><|��<r=,��< �6;�%�2\���   �   c'н.�X3��~譾u�ݾ-���$�+���6��:��m7�O-��8�ޫ���⾂%��0��zD7�L_ག#[�H�9��Z�<��=�=��<p�λh@��,н�.��5���뭾��ݾ�/���F�+��6�o�:�Oq7�sR-�<�ʮ�� ��)���3���I7��g཈/[�Ȧ9�P�<޴=8=��<��λ�@��   �   :3P�qѽ��&��2l��Z���ѽ�m�ݾ{0����:����S��6�/þ�U��u�x�N�3�l&꽺�~�����PZ<0��<z=���< �6;�*�5`��|]#��f}��y��;��w�43�/�M��yb�(p�u���p�d�>�O�%g5�5���.�(���Ł��%(�{ۻ���@:Y; ��<P�=�^=��<xa)��   �   Ъ�b�9��c��Z>�,�D��y�C�� ����n��F������0��5���>`��CR����j׽\_x��y���L�;���<�=�=�0u<�����醽.$	�`�c�"�Qj�����`?�.�c��避a���㖿�㙿�W��t��K삿Ƿe��EA��n����|�����e�p	�� ���MS��	�<2�$=V�:=a=�i�<�   �   ��<�G:���������ֽ�H��O3��N�?�`��Hh��Od��zU�QP=��%�.���^�����I��ܑ��
	<�X�<��=:� =T��< V_;���b7ɽ	9�fC����־���Z�=�9j�����{���m��=�����������0���`��vc��ƛk���>�	��־Ĝ��l6��ﾽ�Y��؁V<>�%=T�[=�L`=`�9=�   �   �1]=*P=�k<�!7��7��4��>���mOܽT����9��A��?뽡�ʽa�����`�����Piл��u<��=��1=F�@=��(=@��<���vo�x��іg��}��j� � H.�	`�j���P��������ȿ~�ӿ�׿1$Կ�`ɿ�b��ԥ�������H`�(.��9 �-o��`�a������E��;�l=��q=���=�V�=�   �   2�=�߁=0OE=��<�j0<p���Ѽ��!��I�n\�ZY�P�A�8�����`���XL<Hn�<f�=�PJ=d�_=��W=*=T��<L����坽(�!��~���.оt���F��U~�Ґ��^���i�ο+��M��R>�k/��dϿA���􋛿C�}���E����V�̾�A�����ǃ� ]����=��~=p��=Jk�=�   �   �\�=F��=��=��n=�*4=���<o�<`��;@v��	�� ����p�;@F]<���< �=�
==2�a=<�y=։}=Hxe=�'=pib<<��c���t8�ߘ����}#��3Z�-������)�ƿS���J���E����BY��z�������ƿx@���l���X��3!�0e�c�����+�E5���<���=K�=jE�=\;�=�   �   ���=E}�=0ƭ=�ݘ=�y�=��S=�i(=0H=��<�^�<���<���<�/�<<:=��-=�vO=�o=��=!g�=0-�=�l=�(%=x�.<,���н�G�\d���p����,�&�f�O���x���Iѿh�T� �`��Z
�N���� ��3���п��������$zd��w*�x4��m��.89��L��d7��ԣ=d��=լ=ȶ�=�   �   gܰ=n,�=��=O��=�U=Z�#=̫�<��<�+`<0< �7<h�u<���<��<��%=�pP=�Cw=�"�=�-�=���=��b=�=��껋�������ዾ�k޾��#���c��.���A����F��~����$�h?.�l�1�2=.�N�$�ļ�FD���㿉໿W���n�`�D!�W=پˮ��Ů�:�a��H�;�;=�(�=�ѩ=�   �   i�=��=�=~�l=JQ6=���<��<`(< �2; Ĺ ��9c�;�D<�D�<�(=�6=
Rb=��=�E�=ȅ=�_=��= �ĻW����{�,�����پ�� �&�_�o�������;�fz��p��*"�~8+�j.�n?+��$"�6G��!��5�vи��<���\��F���Ծ����P����X��+�;��:=ҿ�=�l�=�   �   ���=�J�=�v[=R�=$�<`��;��.��ں����d��z��ܺ�����@Ȝ��z#<���<�;"=2ZR=�Yp=v�s=xS=`F= �3��j�Ә��d� �̾���1�S��닿���i+ֿ�����n���"�l�%��"��1�<+�������տ�௿#튿IhQ���TxȾ�sv������?��<	8=�A�=���=�   �   ^�i=�>4=d��<`]w;@z���&-������J��tŸ��½����:̫�镎��qQ� ���H���M<���<n�1=r{J=�>=�=��:�l?�����GDc��W����	�ı@�����!��L�Ŀ'�b�����Z�v �������� �yp��ĿIʡ�J�~��O?�E������6�[������ �I<f1=��q=ੀ=�   �   *�= �@<p�}��e?�:�����(�d�'�N�7���=�� :���,�������ķ��am���� (�̒�<�Y=�=\B�<�0�;��
���ƽ��?�g���X1���(���a�����ٮ�p�̿M?翽=��F��0o�|>�*-��p?�:�Ϳ;V��ݨ��pGa��/(��b�K���s:�x๽�Sؼ4i�<bd#=I=>�<=�   �    �u9����3��BF�n&�V/U�q8��o��ɀ��ƽ��Ĝ��咾����]��V0�R��O���/��(��X<�-�<�M�<Pn<<���p���n�A�����ƾ+���	?�_�t�MÕ�����'ǿspٿ(O�ѣ�+�忂�ڿ�eȿ7$��������u�D�?�����Pƾh�����k_���p��w�<�=�`=�o�<�   �   >�+��ﴽ�o�y S��󊾰�����Ⱦ3q�^�ﾇ����7�Q �+�̾6���̏��]��Q�E�ǽ@�O��o�@�<��<��h< >�JC�xཛྷ�G��C�� �㾻��CH���v�����s��$��5��B�¿������JĦ����P�x�v�I��9�g:�	ԝ��G�wݽZ9���r�$%�<(��<�ރ< �ڻ�   �   �%���g"��jp�-����Ѿ~���U��(�"�1�,�y�0��-��
$�������վoZ���-y�(X*��<Ͻ��K�U�P�<x<k<�bs;�{ȼ�������j�ͭ�@���[�B�b�g����[���p^��s������\��d6j�X@E�?���b����Sm�y���M�� �ż01�;��<@�K<���l3��   �   �� �`�x�A��ˌ�ѻ�O�/���I��t^�9�k�{�p���l�9`�:L�wX2��+����峾�~���%��Լ��#%�p�»��:<��D<����n[�뺴�K� �R�x����O�龖����/���I�Op^���k��p���l�5`��L�cU2�X)�}��s⳾U�~���%�Zм��%� �»��:<0zD<�4���f��´��   �   �$j�ѭ�E�;����B�~�g��������`���u��l𙿹���^���9j�%CE����9f�Q ���Wm�ڝ��P����żP5�;�<�K<x���^3�����a"�vcp�����]Ѿ@}����y�"�d�,���0�@�-�J$�������վ�V��:(y�T*��6Ͻb�K��U���<p4k<�s;܌ȼ�������   �   *G����㾀�GH�|�v�$���su������!����¿{��� ��DƦ����*�x���I�R;�=��՝���G��yݽ�\9���r�*�<H��<L�< Nڻ`�+�8洽�i�S�Q����E�Ⱦ6k�*��V����1��'�̾�	���ȏ��]�&M���ǽ�{O���o�x
< ��<`�h<Pm�ZTC��མ�G��   �   ~�ƾv���?�Ʃt�Bŕ����k)ǿ�rٿ�Q�D��~�忣�ڿ�gȿ�%�������u��?�����Rƾ�������`���p��{�<�=4g=T��< ��9D��y*���:��g&��'U��/�>k���{������y���eᒾ���D�]��P0�zM��H���.��b(�pX<1�<�K�<X`<<�,��%u���r�߯���   �   �4�,�(�T�a�����oۮ��̿�A�@��r��Tp��?�/��A迣�ͿcW��ȩ���Ha��0(�Ud�L���t:�\ṽ�Sؼ�l�<�g#=
$I=0�<=Z�=��@<��}��T?����彀"���'�<�7���=���9�V�,�L�����y����Sm���ༀ2�P��<�\=~=t?�<��;��
���ƽO�?� ����   �   8�	�ѳ@�^��j#����Ŀ� �\�����[�p!�v�����`!��q���Ŀ�ʡ�H�~�;P?����!�����[���F����I<(1=��q=���=*�i=,G4=@��<`#x;|]���-�����BA������	½N���ië�񍎽dQ��i��Pc�88M<D��<�1=}J=�>=�=@��:�s?������Gc��Y���   �   ���S��싿C����,ֿV��T �8�`�"�(�%���"�v2��+�~����տ ᯿^튿�hQ�%��gxȾ�sv����t�?��<x8=XC�=���=\��=M�=�}[=v�=��< �;@q.��º�����*������� 䐼�����#<H��<X@"=N]R=�[p=
�s=bwS=2D=`"4��j�����g�6�̾�   �   �� �m�_�-�������<��z�lq�.+"��8+�hj.��?+�%"�\G��!�6�qи��<����\��F�B�Ծ�������"�X� >�;� ;=���=@n�=�j�=Ə�=��=��l=4V6=t��<|(�<`@<��2; �� g�9���;�D<hL�<�+=��6=�Sb=�=�E�=�ǅ=�_=��=��Ļܘ��[}�b�"�پ�   �   3�#���c�_/��fB��(�z�������$�z?.�n�1�"=.�.�$����D�z��໿񽔿��`�vC!�Q<پ���������a�p^�;.�;=o)�=�ҩ=ݰ=�,�=n�=˵�=ҘU=$�#=��<��<8-`<P0<p�7<0�u<���<X�<>�%=�oP=�Bw="�=O-�=N��=L�b=�=��q������~⋾�l޾�   �   �� �`�_���������;�Tz��p�x*"�08+��i.��>+�j$"��F�.!�5࿩ϸ��;����\��E�%�Ծ̽�����D�X��M�;.;=n��=�n�=�j�=Ꮱ=�=��l=JV6=���<�(�<x@< �2; �� r�9@��;�D<�L�<@,=؞6=$Tb=B�==F�=Qȅ=�_=��=��ĻN���>|�������پ�   �   ����S��닿�����*ֿ7�� ����"���%�L�"�&1�~*�o���X�տ�߯�&슿�fQ����GvȾ�pv������?�p#<�8='D�=��=���=�M�=0~[=��=�<��;�p.��º����� ��~��\��P㐼 ��� �#<���<A"=<^R=�\p=��s=jyS=G=��3��j�ۘ��d��̾�   �   #�	��@����F!��i�Ŀ濸����Z������������n�k�Ŀ�ȡ���~��M?����/�����[�P佞���I<�!1=��q=9��=�i=�G4=���< 'x;0]��|-�����1A�������½+���<ë�����tcQ�@h���_�X<M<���<��1=2J=l>=�=@H�:Rk?������Cc��V���   �   �/���(�#�a�"���dخ��̿�=��;��8��n�T=��*��C=�3�ͿgT��D����Da�a-(�~_�I���o:��ڹ�LAؼ�x�<�k#=�&I=ڥ<=f�=H�@< �}�NT?������}"���'�8�7���=���9�>�,�+�7�������Rm�l�� ����<<_=�=I�< H�;��
���ƽ<�?�j����   �   ,�ƾ���'?�/�t�����
���1%ǿVnٿ�L�c�鿱���ڿucȿ"��Ƞ��(�u�s�?�s��GMƾ������KY����o���<��=j=��< G�9���>*���:�g&��'U��/�;k���{��򸟾q���Yᒾ����]��P0�3M��G��l�.��Z(�X X<�8�<hV�<~<<���|m��m�����   �   �A��m����fAH���v�F���$q����������¿����h������� ��q�x� �I��6��5從Н�J�G�#oݽ�M9��r��7�<|��<4�< ?ڻ4�+��崽�i��S�J����E�Ⱦ4k�&��P����1���̾�	���ȏ��]��L���ǽ�yO���o��<���<�i<���DC�����G��   �   �j�Xʭ�y<������B��g����?���*\���p���뙿8����Z��E2j��<E�#���]����Mm����@F���tż���;l�<��K< ���\3����a"�`cp�����YѾ>}����x�"�d�,���0�=�-�F$�|����v�վ�V���'y��S*��5Ͻ��K���T� �<�Qk<�s;oȼ����D���   �   �� �h�x����)������/��I�kl^���k���p�B�l��0`��L��Q2�&�����ݳ��~���%��Ǽ��%��E»0�:<p�D<�؈��X�(���� �.�x����J�龔����/���I�Pp^���k��p���l�5`��L�]U2�M)�c��S⳾�~�3�%�1ϼ�L%��|»��:<��D<@ǈ��S������   �   4��|]"��]p������Ѿ�w��ڠ�}"���,��0�u�-��$�	�����վ,R��� y��M*�-Ͻ�K�P�T��<�\k<�s;�tȼ�������Sj��̭��?���[�B�c�g����\���q^��s������\��\6j�O@E�4���b����Sm����dL����ż�_�;x�<x�K<xy� U3��   �   v�+�ߴ�e�!S��늾T���N�Ⱦ�e�;��*����+�㾂�̾���mď�2]��F�\�ǽ�kO�P�o��6<���<�i<���GC���Y�G��C���㾷��CH���v�����s��$��7��C�¿������JĦ����I�x�m�I��9�L:��ӝ��G��uݽ�V9� tr�t3�<���<���<�ڻ�   �    �9Н�#��j1�b&�� U�(��f��aw��0��������ܒ�j��V�]��I0��G��>����.��-(��AX< D�<�]�<@�<<����n��pn�+�����ƾ'���	?�^�t�LÕ�����'ǿspٿ(O�ѣ�+�忁�ڿ�eȿ5$�������u�<�?�����Pƾ@���,�^����o�h��<R�=Zl=���<�   �   �=��@<�}��F?���������:�'�t�7���=���9�x�,�����������Am�l�ༀ	�l��<�e=h=�N�<@R�;8�
���ƽW�?�X���S1���(���a�����ٮ�q�̿M?翿=��F��0o�|>�*-��o?�8�Ϳ7V��ۨ��jGa��/(��b�K��Js:�o߹��Mؼ8r�<�j#=�'I=H�<=�   �   ��i=FM4= ��<`�x;�E���-�����|8��E���H½�~��ع��섎�tSQ�L��h/�hdM<��<ܘ1=�J=�>=x�= t�:�j?���� Dc��W����	�ű@�����!��L�Ŀ'�d�����Z�v �������� �yp��ĿGʡ�F�~��O?�>�������[��佬����I< 1= �q=>��=�   �   �=XO�=��[=z�=d&�< P�;�I.�䬺��������`����� ͐�P.��P�#<H	�<�G"=�cR=8ap=
�s=&|S=:I=��3���j�����d��̾���/�S��닿���i+ֿ�����n���"�l�%��"��1�<+�������տ�௿"튿DhQ����DxȾ�sv����~�?��< 8=�C�=���=�   �   �j�=f��=��=v�l=ZY6=$��<l1�<xT<`T3; )�� d�9�;�,D<TW�< 1=�6=�Wb=��=�G�=Ʌ=�_=�=`�Ļ����{�&�����پ�� �&�_�n�������;�hz��p��*"�~8+�j.�n?+��$"�6G��!��5�wи��<���\��F���Ծ󾃾4����X�P4�;& ;=���=Zn�=�   �   ��=��=�\x=�?E=�
=�9�<�>�;���e@�Ȥ)�0O����z;Ȳy<T��<�<)=��Y=��}=@[�=�|=~�A=e�<|����νr!S��״����.�L�ج�������s�T�>�"���8�T�J��JW�&�[�JFW�d�J��28�"�JH
���俼+��N	����I��\
�j���*�K��;��<���|��<2�`=�s�=�   �   ,�=��=��^=��%=4�<��"<�x���q�����tͼ���0+��0O��p��;$ќ<t 
=�@=�j=t.~=R�r=�<=p7�<�� ɽZ5N�����
�4�H��1���ش�������F��DI5�%G��4S�d�W��=S��G�F
5��a�"����3������IF�1���
����F��ٺ��ꦼ��<΋[=Ze�=�   �   ��p=N^L=�=tq�<�~'��ų�f,!�>#Z���,V��b΂���e�`�1��ݼP;�@�*<��<�-=ƶQ=^U=�E-= �<��¼�n��@�� ��I�s�=�0�������|׿N����4�+�΁<���G�P�K�B�G���<�v�+�|�����q`ֿ����rǁ�b�;�
" �����>j9��n��������<�J=v�s=�   �   P�!=H��<�+;!���`P��1����н����F��V���x
������)ٽq����7i�����б��0>�<�=�!=�a=�y�<h?��{S��t6*�]+���z��,�qko�p���}ƿWp�*�������,��k6�&:�º6��-�
1�V���c�ӫſ�ל���m��Q+�rz辘R��L�$�l��`�S�$��<�5,=��==�   �   ��6<0f��Z>��g��w����G%�H�H���d�FQw��M~��y�s>h��^M�+��`����)Z����@t�;(,�<x��<�=p<иX��ွ�����C̾�4�ʺR��^��}����*տG����V��+��!�2�$�p"�����+����տi)���:���R�cP��Lʾ�{�_�
��eo�����ģ<��<T��<�   �    _�9�@�罠�*��Td�V�������ڻ��ɾ��;F'ʾ�佾�j��H����Kk��1�l���FՓ�*(�� ��P�<HM<�u��lA��i⽎TP��Q��@���MH2�E}m�`ǖ��`���~ֿ��~���,�4��V�� ��S��~�׿�x��/p���n�X2�{���Z����M��ܽ@�3������^<0�k< �28�   �   ᓞ�܍�XgM��D��8����@ݾ�[ �b~����c"�dg�h��4��ᾬ�������Z,T����)����!���;� .(9p.ɻ���Dx�����yg��x2˾���SB�R�x�6�����g�ɿ�uܿ���N�쿁T鿫�ݿ|�˿Z-���\���xz�(�C��,��˾gS�����E��,��� `�@Sc;P���N��   �   S��_�Q螾��Ӿ�f��; �48��@K�n�W��:\���X���L��O:�l�"����ϥ׾xI���d������@e�PEY� fܻ�â�nH]��{㽴�E�l�����߾�!��uD�2#r����/f����������qS���[��)���������t���F�M����Oś��#G�rm�n9\�|I��`���(�5�ھ�Į���   �   �U\�b���Ĝ�S)�8[8�k][�&wz�����h��� }��5��U���6}�^���:��C����5!����_�d�	�7擽PM ��3��J.��g���`����O\����V��&�SW8�Y[�Qrz����ǆ���z����������
}�h^���:� A����N����_���	�"㓽�J ��3��].��x���g��G��   �   &���z�߾%�lyD��'r�8���h��t�������JV���^������Y񣿛�����t���F�l��H�ᾉǛ��&G��p�v<\��H�� ���`l5���������M��_��㞾�ӾNc��7 ��/8�<K�ݡW�S6\�R�X���L�L:�1�"�؛�o�׾F���d���|���B`�(@Y�`wܻ�Ϣ��R]�c��(�E��   �   �6˾���#WB�R�x��������3�ɿ�xܿ���G��WW�I�ݿԩ˿`/��w^��y{z�L�C�.�&�˾�T������F������`�_�`�c;����A�
�����`M�\@��䲵��:ݾ#X ��z�ٳ����c���&
���7��� ����&T�Ŏ��#��P�!�0�;� v(9@GɻT���}�����zj���   �   ����K2���m�hɖ��b��,�ֿ�����P.�������F�����k�׿yz��xq���n��Y2����T\��`�M��ܽ��3����� �^<X l< \88C�*놽��罯�*�FLd�_Q��U����Ի�(ɾ�;�!ʾ�߽�(f��&����Dk�n�1������Γ�2��Ԯ���<xJ<���*tA��o�YP�U���   �   �6�z�R�9`��n���-տ����4X�-���!���$��"����	�����m�տ�*��X;���R�<Q��Mʾ:�{���
�"fo�P���ˣ<$)�<\��<��6<H�e��I>�-]��J���A%���H���d��Hw��D~�6y��6h��WM��+��[�c�� Z��������;�3�<���< 8p<8�X��倽��d���F̾�   �   ��,��mo�놝�:ƿPr�D��"��
�,��l6�j:��6��-��1�����d￞�ſs؜���m�R+�{��R����$�'��h�S�T��<v:,=�==4�!=4��< �;���jOP�3(���{н����\��m��;s
�,����ٽ�쩽J)i��y��@j��@K�<l�=>�!=�a=�u�<�H��UW��_9*�x-���}��   �   >�7���9«��}׿����,�+�Ԃ<���G�F�K��G�8�<� ,������`ֿІ���ǁ���;�" ������i9�n��𥍼8��<��J=��s=�p=eL=:�=���<��&������!��Z����N��Gǂ�b}e�n�1�DsݼP�H�*<D#�<�-=&�Q=�^U=:E-=L�<��¼9r���
@��"�����   �   t�H��2���ٴ���⿊������I5��%G�N5S��W�\>S�G�t
5��a�*�����2�������IF��� 
��
�F�;غ��妼��<|�[=�f�=�-�=��=�^=&=�'�<��"< �w�h�q�p���`�̼������@#���ş;�؜<n#
=,�@=Lj=�.~=��r=��<=x2�<� � ɽu7N����
��   �   ��L�M���_���bt濘���"��8���J��JW�&�[�4FW�8�J�f28��"�H
�t��B+�������I��[
�t�����K�u9����|��<&�`=^t�=���=5��=�]x=�@E=�=�;�<�D�; ����d@�P�)�pR����z;��y<���<�;)=��Y=j�}=�Z�=��|=��A=`�<@���ν�"S��ش�S���   �   �H��1���ش�������,��I5��$G�H4S���W�X=S�G��	5� a�����32��\����HF�?��.	����F��ֺ�8ᦼ��<z�[=$g�=�-�=��=F�^=&&=�'�<��"< �w�`�q�t���H�̼�������@"�� ǟ;\ٜ<�#
=��@=�j=�/~=��r=��<=�5�<��3ɽ!6N����
��   �   I�=��������|׿ �F����+��<���G�Z�K�@�G���<���+�������_ֿ^���sƁ���;��  ������g9��j��@������<b�J=��s=��p=teL=v�=���<@�&������!��Z����N��Aǂ�D}e�<�1��rݼ �@�*<x$�<��-=6�Q=Z`U=bG-=p�<��¼�n��"@�� ��8��   �   z�,��jo�ӄ���ƿIo�~����,�\j6��:�z�6��-��/�D���a�'�ſm֜���m��O+��w�tP��$�$����X�S�0��<=,=��==6�!=p��<@�;\��LOP�,(���{н����[��j��2s
�����ٽ�쩽�(i�\x���c��`M�<ܳ=J�!=�d=8~�<�;���R���5*��*��Az��   �   �3���R��]��b����)տ�����U�v*���!���$� "�:����������տ�'���8��	R�QN��IʾJ�{��
�>[o����hգ<@/�<(��<X�6<��e�tI>�]��B���A%���H���d��Hw��D~�/y��6h��WM��+��[���>Z�(���0��;�8�<���<�Lp<ЫX��߀���S���B̾�   �   ����F2�<{m�Ɩ�_���|ֿ�
�8��h+����֛���������׿�v��.n��tn�`U2�<���W����M��zܽį3�������^<�l< �d8�@��ꆽ��罠�*�=Ld�_Q��V����Ի�(ɾ�;�!ʾ�߽�f������Dk�>�1�6���,Γ�T�@��� �<a<`d��gA��f�zRP�XP���   �   0˾L���QB���x��	������ɿ2sܿ�}�]�쿄Q鿼�ݿ��˿�*��vZ���tz��~C��)�ǥ˾LP�����=��d���`f_� d;����?�f������_M�U@��ವ��:ݾ$X ��z�ڳ����c� ��!
���$��������&T�s���"����!���;� ..9�ɻ���t��.���e���   �   ���`�߾���rD��r������c��#��������P��Y��Z���c죿'���<�t�6�F�5��2��~���0G��d�h+\�x1�� `��X5�n��ɥ��PM�`_��㞾�ӾNc��7 ��/8�<K�ޡW�S6\�P�X���L�	L:�*�"�Л�X�׾�E��ȣd����@����\�H*Y��6ܻ����,A]��v�\�E��   �   �J\�%���i�⾁#�=T8�ZU[�!nz�����J����w����j���}��
^���:��=�G������_���	�ۓ��= �h�3�`..�d^��e_����N\����O�� &�SW8�Y[�Srz����Ȇ���z����������
}�c^���:�A����,��f�_�(�	�wᓽF �H�3�2.�8Y��8\��^��   �   �I�_
_�[�����Ӿ�`��4 �G,8�8K���W��1\�ŀX�5�L��G:�c~"����ƛ׾tA����d�<��m󨽶Q��Y��ܻ`���tD]��z�X�E�S�����߾�!��uD�3#r����1f����������rS���[��'���������t��F�B����&ś��#G�l�5\��<���n���Q5�4��#����   �   ����̃�jZM��<��}����5ݾ U �jw�B����`�`����l�Γ��l�GT����1����!���;� �39p�ȻJ���v����Vg��e2˾���SB�R�x�7�����h�ɿ�uܿ���O�쿁T鿩�ݿ{�˿W-���\���xz��C�w,�Ʃ˾9S��,��GC��X���`�_��d;����Z8��   �   �.�Z䆽 ���*�hEd�JM�������ϻ��ɾ:�;�ʾ�ٽ��`��^���N<k�N�1����;œ����n��
<pr<�\�|hA�:h�/TP��Q��4���JH2�C}m�aǖ��`���~ֿ�����,�4��V�����Q��{�׿�x��,p���n�X2�c���Z��F�M���ܽ�3��Ӝ�H�^< l< �z8�   �   �
7<(�e�~<>��T�����;%���H���d�@w�w<~��y�g.h��OM�� +��U�����H
Z�۩�`
�;4H�<���<XZp<8�X�
���b�����C̾�4�ɺR��^��~����*տG����V��+��!�2�$�r"�����*����տh)��:���R�ZP��Lʾ��{���
��bo����ӣ<2�<��<�   �   ��!=���<��;x쿼RAP����Krн���������Xm
�����3ٽ*㩽�i�D[��p���`�<��=$�!=�h=��<�8��]R�� 6*�F+���z��,�pko�p���}ƿXp�*�����,��k6�&:�ĺ6��-�
1�V���c�ҫſ�ל���m�{Q+�_z�{R���$�B
��H�S����<X=,=��==�   �   &�p=XiL=Ԫ=Ȓ�<�B&�4���!��Z�"���G������oe�ԇ1�<Zݼp���+<h4�<V�-=|�Q=�dU=�J-=�#�<��¼n���@�� ��F�s�=�0�������|׿N����4�+�΁<���G�P�K�B�G���<�x�+�|�����q`ֿ����pǁ�^�;�" �}���j9� n��|������<ؗJ=��s=�   �   3.�=��=X�^=&=H/�<��"< Qw���q�h���t�̼�쿼����������;��<�(
=�@=h j=�2~=~�r=D�<=�:�<X༳�ȽB5N�����
�4�H��1���ش�������F��DI5�%G��4S�d�W��=S��G�F
5��a�"����3������IF�/���
����F�Uٺ��覼\��<$�[=�f�=�   �   �yz=i=�>=��= ��<�>�:P<U��Ƽ�� ��A�����Ѽ �u�@X��h�c<d4�<�1=��[=m=�CZ= �=`(];$T����(��K�ݾ%	*�x�t�>����ؿX�J�#�P�@�Z�\�Ʋt������������V�t� \� �?� �"��7���ֿ⤿ݴq�@�'�C5ھ^\��
+�*�D�`!�;<d#=��g=�   �   �~i=� R=th!=��<к�;P3���׼�3���>��dK��,B�9$����[���b;(�<�c=:�D=�!\=��N=B�=��W;�XN�Gc��J���\پ'�&��Gp��֣��տ��� ��.=��^X�X�o���� Ă�H��z�o�NX��<��  ����#ӿ�&��h�m���$���վI3����?�p[�;Y=�^\=�   �   �5=
=D��<��Q��hҼ\�C�ja������8����ǽkm��C���1����N�H뼠Gѻ��i< D�<TJ(=|5,=,��<��8;$>�"����t���̾��9�c������ʿ�.�����@H3��\L�|�a��ap�\�u���p�:�a�$oL�L3��^������"ɿB/��lDa�:��f�ɾEo�)�����/���;�f
=�M9=�   �   �<औ;ؚ��~M��:�����@��)H&�L5��{:��6�HQ(��o����3��tT[��ü���:ޜ<�
�<�!�<�>�:,�&���4�Z�ݴ��F�;�O��y��$�����(���Z$�@�:�� M�N�Y��x^��7Z�½M��;��$�ʋ��v�<]��<����N���)\���V���ٽLG��M�;ܛ�<h4�<�   �   X]%��� �8L��=���Ο)�<bW��8��ϗ��`D���2��'����鑾�����f[���-�N�������`�.�Y�p�;H�!< �R��꽽E;��ȟ�f���0]6�N�{�^4��SgϿSl�����%��4�Y?�fEC���?�֥5�p &�����.��[�Ͽ#��H�z��z5������"��8��\��"a� B�9��N<�?<�   �   X_��@˽0,�C+^�-Ð�����VFϾ���a1�����`+���辱�Ѿ^Q���_���c��|"���ҽT�k�T9ϼ�&�p��<*����n�o����о���uV�5b��z]��Q�׿G������&�#���&�ZE$���\�m����7ٿ������V�q����Ͼ\��Bm�k���@4��ֻ`Ά(޸��   �   ���5�X��㙰�v�*�����U,��
7�"�:�G�7�Փ-��w����_�z����υ���9�o�z΅� ��Ҡ�K޼��l��u�ƣO�����J���%�.�A�h�Tғ��Գ��_ҿ�d�o��y������N�}iￇAԿS��0ڔ�j�i��R/�!��Ԓ����N��U�Οg��'Ҽl���`��������   �   ��=������7ž���"�!��+A�
]��s�\���YZ���1����t�3_��oC�+�#�[��ȾA���H�@��6�ℽ�����z�2���0����|�����Ti�<�7��Lk����=l�������`ѿ��ܿL�	�ݿ��ҿ����c$��v����~m��&9��V	�������}�@/�$���0o0�$�߼���C�������   �   ����:�ʾ�G
��3��E]�����锿����L������{񬿪>��:S���`���_�;"5����Ȱ̾���>+5�7�ս��h����jD��f�wӽ&e3�ٸ��8�ʾ�D
��3�A]�_G政����I��������;���P���^��m�_�H5����[�̾D��(5���ս��h�����I���f��~ӽ�j3��   �   ���0l�ԫ7�@Qk�K��o���¿��cѿ!�ܿ��2�ݿ��ҿg����&��i�����m�[)9�~X	�V�����}�P1������n0� �߼r��ߌ��e��S}=�x���:2žJ��F�!��'A�A]��s������W��f/����t��._�lC���#�tX���ǾK����@�x1�߄�P�����"�2��������|��   �   ���C�.� �h��ԓ�2׳��bҿ�g�tq��{�\����DP�3l��CԿ�T���۔�� j��T/��#��������N��W�.�g��!Ҽd���l���E���~�H�5��S������4�p&����WQ,�#7���:��7�ۏ-�Ft�����Y�?���J̅� �9�Jh�ʅ�����Р��Q޼��l�F|뽱�O� ����   �   U���	V�/d���_����׿L���������#���&�G$���������9ٿ��C����V������ϾX��7n������/���ֻ0���tƸ�D�^� 6˽�%�&#^�[���k���-@Ͼc�澊*��>����$������Ѿ~L���[��Xc��w"�\�ҽ��k�L,ϼH�ؘ��2����Nr���2�о�   �   �_6�k�{�C6���iϿ�n��B�� %���4��Z?�2GC�D�?�N�5��&����O0����Ͽ����z��{5�����#���8��\��@_��( :`�N<Pd<X,%��� �VB��2�����)�ZW�^4������X?���-��D���呾����|_[���-�������.�(�X��9�;X�!<��<�'ｽ�;�3˟�����   �   |�O�{���%�����P��
\$�:�P"M� �Y��z^�P9Z��M��;��$�d��w��]�������N�z���\��Y�V�H�ٽbE�i�;���<B�<�<���;�~���M��0��5����zA&�`�4��t:��6�K(�:j���{+���F[��ü �:h�<��<�"�<���:R�&�z�ཛ�Z�S������   �   #�c�.���Q�ʿ]0�����XI3��]L�Լa��bp���u���p�$�a��oL��3��^�4���F#ɿs/���Da�J��^�ɾ8Eo�M�����/��&�;�j
=�R9=&�5=�=أ�<`"Q�OҼ��C��Y��3�������Uxǽ!e������9�����N����Pѻ��i<,M�<M(=�6,=ܯ�< �8;"!>�/����t�̾a���   �   ]Ip��ף��տ��z� ��/=�z_X�2�o����[Ă����ީo��X� �<��  ����#ӿ�&���m�B�$�1�վT2�6���?�`r�;\=b\=��i=L%R=�m!=<�<0��;��2�$�׼D+�2�>�L\K� %B��1$���0�[��#c;$"�<*f=��D=�"\=B�N=��=��W;]N��d�L��G^پM�&��   �   b�t�Ĵ��w�ؿVX���#���@���\��t��������������t��\���?�ҥ"�l7� �ֿ�᤿��q���'�#4ھ�[���)��|D��7�;lf#=x�g=~{z=�i=F�>=&�=D��<�]�:9U��ƼV� ��A����ȳѼ`�u��r����c<02�<��1=��[=�m=BZ=̤=��\;�'T�9���)��v�ݾ�	*��   �   AHp�ף��տ��� ��.=�h^X��o�4���Â�~����o��X�L�<�H  �`��"ӿ&���m�w�$��վ�0�:��,?���;4]=�b\=�i=�%R=�m!=h�<`��;��2�,�׼Z+�6�>�P\K�%B��1$�����[�@&c;�"�<jf=�D=#\=�N=�=��W;JZN��c�PK��#]پ|�&��   �   �c�͂����ʿ:.��<���G3��[L���a�x`p��u�8�p���a��mL�<3��]�'����!ɿ .���Ba�ʰ�B�ɾ^Bo�������/��@�;�l
=T9=�5=*	=`��<�Q��NҼ�C��Y��9�������Uxǽ&e������,���|�N�\�꼠ѻ��i<�N�< N(="8,=X��<@�8;>�D����t���̾Ս��   �   ��O�y��a#����迈���Y$�6�:�bM���Y�Dw^�&6Z�&�M�0;�̞$�����t迖[��ݟ���	N�g���Y��d�V��ٽ|>����;���<�E�<,�<0�;�}��dM��0��6����}A&�f�4��t:��6�K(�0j���I+���F[���ü �:4�< �<�(�< ��:>�&��ཊ�Z�V������   �   &\6�ڵ{�`3��
fϿ�j�����%���4�ZW?��CC���?��5���%����1,��.�ϿI
��:�z�ox5���� ��8��V���V��:(�N<�l<X'%��� �&B��"�����)�ZW�b4������\?���-��F���呾����m_[���-�G����綠��.���X��M�;(�!<������载 ;��ǟ�����   �   ����V�	a���[��w�׿�����j�v�#��&��C$�����r���5ٿI��(����V����B�Ͼ���i��󔽰� xֻ ���������^��5˽w%�#^�Y���l���0@Ͼg�澍*��?����$������ѾtL���[��2c�dw"�ƭҽ��k��&ϼ�P��l ����m�<����о�   �   ����@�.���h��Г��ҳ�K]ҿ�a�<n�Px���V��M�@fￎ>Կ^P���ה���i��O/�G��5���.�N�EM�b�g��Ҽ|�������������5��S������4�q&����YQ,�&7���:�	�7�܏-�Bt�����Y�-���0̅���9�jg��ȅ�����Ġ�0?޼p�l��q��O������   �   ���sg���7��Ik�����i������]ѿ��ܿ	Ώ�ݿ��ҿ�~���!���2zm�E#9��S	�B���ƃ}�&*�-����a0�d�߼������S��}=�a���02žH��F�!��'A�C]��s������W��g/����t��._�lC���#�lX�s�Ǿ(�����@�70�-݄�f����漠�2��	��h��È|��   �   O�����ʾNB
��3�}=]�B삿�㔿)���F�������묿�8���M���[����_�d5�i��B�̾T��"5�B�ս��h�`��d<��f��uӽ�d3�����(�ʾ�D
��3�A]�bJ政����I��������;���P���^��f�_�B5����=�̾���'5�ϘսJ�h����p=��f��qӽ~a3��   �   �x=�r���<.ž���%�!��#A�]�s�0���U���,����t��)_��gC��#�&U� �Ǿ����j�@�'��ք�f�����x�2�������C�|�����Ni�9�7��Lk����>l�������`ѿ��ܿM�	�ݿ��ҿ����`$��s����~m��&9��V	������}��.�Ҩ��h0���߼��������   �   
��K�5�uP��p��� �_#�o��pM,��7�f�:���7���-�Ip����S�想��ǅ��9�>]�[���Z��ķ��H9޼��l��s�:�O�x���9���#�.�A�h�Tғ��Գ��_ҿ�d�o��y������N�{iￃAԿS��,ڔ�b�i��R/�� ������ �N��S�ޙg��Ҽ������ŝ���   �   l�^�>.˽h ��^�V��������:ϾI���#��r������!���Ѿ�F���V���b��p"�U�ҽ�k�xϼp��l���'��n�=��h�о���sV�6b��{]��R�׿I������&�#���&�ZE$���\�k����7ٿ������V�g����Ͼ"���l�����%�@{ֻ`i�������   �   �%�� ��:������)�SW�T0��x����:���(��E�:���.�GW[���-�<����夽<�.��X��;�	"<������载�;�qȟ�V���.]6�M�{�]4��SgϿSl�����%��4�Y?�hEC���?�֥5�p &�����.��[�Ͽ!��C�z��z5������"���8��Z���[� (:��N<�~<�   �   X#�<�A�;,i��"�L��(�����v��T;&���4��m:�6�\D(��c�^��i!���5[���ü�x�:���<�!�<�2�< ��:@�&����ګZ�Ŵ��A�:�O��y��$�����(���Z$�@�:�� M�N�Y��x^��7Z�½M��;��$�ȋ��v�=]��:����N���\����V�G�ٽdC�P|�;���<$K�<�   �   5=�=԰�<��P�;Ҽ&�C��R����������oǽ�\��?쭽f���@�N���`�л��i<�]�<BT(=�<,=��<�9;�>�Z����t���̾��9�c������ʿ�.�����@H3��\L�|�a��ap�\�u���p�:�a�"oL�J3��^������"ɿB/��kDa�5��V�ɾFEo�f���^�/��,�;.l
=6U9=�   �   ��i=
'R=p!=$�<��;��2���׼Z$���>�DTK��B��)$�����[���c; .�<vk=r�D=�&\=F�N=��=��W;DWN�c��J���\پ'�&��Gp��֣��տ��� ��.=��^X�X�o���� Ă�H��|�o�PX��<��  ����#ӿ�&��f�m���$���վ,3�����?�`j�;�[=Nb\=�   �   T
L=��8=�	=��<�(:����L�fY5���U��Ca���V���7�h>���� F�4@�<�G=�c6=̲I=ڣ4=��<p�A��Q��;�-�ܙ��8����D�@K��� �����F��r;��;^�X������s^������Y��)ď��Q���D]��9������.���⊿�B��( ����$�*��ۓ�`/��:�<�;7=�   �   r59=�N=���<8�<��3�����B�@���w���Q+��~��Rvz���C�4���A� �;T��<��=P�6=�'=�^�<�C�I�� �)�2]��;��	�@�j։�<ͺ��� /���7���Y�~�{�o���o�������%���Hx{�N,Y��6��� ���Є��?�js��Zu��`Q'�ʼ�� ~1���<�*=�   �   ��<���<@T�:d����?��C���S���㽷3��tC�c,��l��O������ oD�0Ӻ� k�9p4�<R�<F� =���<�hM����T-��	��/��@�6�β��
���5濊��3.�.�M���l��ۃ��$�������F��m����l��M�X�-�"���俎-��^�����4�3Y�[��2��*��� �;�0Z�<b�=�   �   �;��X�X�(�T����ཛྷ��]�3�W M���]��uc��@^��hN��t5�����I��Y��^�-���i��ݾ;x�r<X�<�Cj���|��������Jپ�0&�o��좿��ӿ�D����l�;���V�>�m� �}��ǁ��+~�t{n�MW��<�������ӿ���:�m�%�$��m׾�T��
�zw���Y��u(<x�<�   �   8��<
� ֽ����Q�.���֙�xI���D��i���и�RE��������c9T���c�ٽ�^��������#��2������<	a�������c�+��~���R��S��&f�����40��B&�8�<���O��\�dsa�<]���P�Ƽ=�� '�N��V���=�����>�Q�*�� л�'�a�!��hr\�0����������   �    /�������D�x���UԬ�%Ҿ����(�����$�����}���+Ծ����|G��6dG�������y5���μ��ӼB�J�!fͽ��<�����L���V�2��`v�tġ��)˿%S��\�D�!�p�0�
;���>�n�;��1�ֻ"��������˿����qv�JE2��������W;� B˽�F��7ͼ�Ǽ�21��   �   ���ܨ_�^���/Ѿ�g����$�4�~}G�vS��W�� T�	�H��a6������EӾ?\���+b�T��LP��`pY���ln?�:������Ƅ{�/'žM)��#J������U�̿�����N�����B��>�������2[οh	��YZ����J�.W�8ž��z����XV��8�<����d�U��贽�   �   ��g�����U�/O��;��_��k~�Б��&���g{������d���:��p2a���=�������i���6�i��2�������f� �D��J��
��H�>�Jl��ſᾡ���RT�Z:��a夿=5���.ڿ���K������ݰ���v���ۿ��¿!S��'F��U�U�_��|���ŗ��>��r�ﻅ��dC��jd��,������   �   �ᦾ�N!�>O�Ͼ~�u&���?�����kWĿ�ȿ�Ŀ�<����������v����Q�Gh"���ﾵ䧾�9]�R%	��ۤ��^�R�]�oQ��l��\\��ݦ�,I�!��9O���~��#��n<��^��TĿsȿ��Ŀ�9��=���%���j���0Q��e"�����᧾6]�6#	��٤�^�4�]��V������\��   �   �������VT��<��2褿e8���1ڿ>��
�������n����y���ۿ!�¿PU���G��#�U�{��|���Ǘ�|�>��t�ܻ��X`C��ad��%��x��b�g�����O�|K���;��_�f~�펋�/���qx�����b��$8��/.a�b�=����0�����y�i��/�|�����f���D�rN�����D�>��o���   �    ,�d'J��ą����M�̿����D�����0�����L��/�d]ο3���[���J��X�@žd{�����V����<�h����U�sഽ���>�_�����6�оqd������4��xG��zS��W�T���H��]6������
AӾ�X��l&b�t��TK��@kY�J��$r?��������U�{�(+ž�   �   %�2�udv��ơ�9,˿+V���0�!���0�H;���>�v�;���1�b�"��������˿A���sv��F2����� ���X;�kB˽��F�D,ͼ�~Ǽj%1�&�����j�D�ޣ���ά��Ҿ���D�H����N �D��Qw���%Ծ󵮾�C��e^G�>�������q5�ܑμ��Ӽ�J��jͽ�<�����x����   �   ԤR��U��Dh��-�뿬1�tD&�,�<�̰O�X�\��ua� >]�h�P�>�=��'�8�����?������b�Q����ѻ���a�a��\p\�0v���d��`��ԙ��~��	ֽ����Q������Й��C���>�������ʸ�%@����������2T�@�įٽeX������#�P$�������a�������c�������   �   �o�-��ӿF�����;�\�V�L�m�"�}��ȁ��-~�}n�bNW�� <��������ӿN����m���$�An׾&U���	�l	w���Y���(<��<pU�;�X���(��J�����9��O�3��M���]��mc�X9^��aN�(n5���A@�3R��v�-��qi���;�r<P�<�Mj�J�|�,�������Lپ�2&��   �   ೂ�]���C7�z��:4.���M�B�l�Y܃��%��[���OG������l���M���-�h����-��z�����4�+Y�y[�����������;��b�<��=��<���<���:�K����?�w;���J��6	��)���>�#�����l���%����cD����� ��9�>�<tX�<�� =\��<@tM�����/��������6��   �   ;׉�7κ����/�^�7���Y���{��������e���J��d����x{�r,Y��6��c ���������?��r���t��vP'�)����q1����<~�*=�99=�S=̰�<@<H�3�����`�@���w�B����&���y��>nz���C�������A��"�;��<b�=�6=��'=\[�<@�C������)��^���<��S�@��   �   �K��^��C������;�d<^���������^������Y��ď��Q���D]���9����}��.��.⊿J�B�( �"�����*��ٓ��S/��?�<�=7=
L=R�8=r�	=$�<�i(:����K��X5�P�U��Ca�
�V�n�7�?�`��� L��=�<�F=Jb6=&�I=�4=D��< �A�T����-�ښ�����֓D��   �   �։�iͺ���$/���7���Y�.�{�.���������o������Hw{�l+Y�"�6�v�h��������?��q���s��VO'�����0j1��<>�*=:9=T=��<�<8�3�����p�@���w�H����&���y��@nz���C�����H�A��#�;|��<��=��6=��'=�]�<p�C�O����)��]���;��i�@��   �   �����~��P5�B���2.���M���l��ڃ�$�������E�����~�l���M�D�-�<�#��I,��U����4��V��Y�����(�����;�dg�<@�=D�<���<@��:DK��r�?��;���J��D	�*���>�#�����g������LcD� ��� 1�9�?�<xZ�<(� =(��<peM����i-��	��,��+�6��   �   Fo�	좿��ӿ\D����r�;�<�V���m��}��Ɓ��)~�pyn�PKW�<������ӿ9��Îm�@�$��j׾�R�����w��Y���(<��< _�;h�X�>�(�rJ�����:��U�3��M�ɂ]��mc�\9^��aN�&n5���$@�R����-� ni���;�s<h<(9j�r�|�'��Y���{Iپ0&��   �   �R�S��e��;��F/��A&���<�ڬO�
�\�.qa��9]�|�P�ں=��&�ޖ�����;��V�����Q���ͻ���a�T��2g\�Lj��@F��@��,����~��	ֽ�����Q������Й��C���>�������ʸ�'@���������x2T�&�x�ٽ�W�������#�����야Ja�o���.�c� ������   �   �2��^v�%á��'˿Q�����!���0�;���>�B�;���1��"������X�˿���nv��B2���������R;��:˽��F�Tͼ�vǼ�"1�`%�����P�D�ڣ���ά��Ҿ���G�K����O �E��Nw���%Ծ鵮��C��7^G����	����n5�8�μ��Ӽ؀J�1cͽ�<�6���N����   �   �'��!J�@���7��%�̿�f��������>��J�����6	�;Xο���1X���J�uT�!ž��z�����N����<�֢���U�1ߴ�����_�x���3�оqd������4��xG��zS��W�T���H��]6�������@ӾmX��+&b����I���fY��}��g?�Ĥ�������{� %ž�   �   ��ᾂ�� PT��8��7㤿�2���+ڿZ������3���$����r�W�ۿa�¿NP���C��F�U�!��w���h�>��i�{����VC�t[d��#������g�����O�zK���;��_�f~��1���sx�����b��$8��-.a�]�=������蠪��i�E/�r���f���D��F��n��*�>�j���   �   �ڦ�?E�w!�s6O���~�7!���9��a���PĿȿf�Ŀp6�����F���܍���Q�b"�3�ﾄݧ�`/]�	��Ѥ�\^���]��N������\�dݦ�I�!��9O���~��#��q<��a��
TĿtȿ��Ŀ�9��=���$���i���+Q��e"�����᧾�5]�M"	�פ�*^���]��L��v��?\��   �   [�g�a��K辚H�)�;�c_�Ra~�I���[����u�����3_��j5��3)a���=�?����*�����i�*�X���,vf�`�D��F����⽉�>�l����ᾛ���RT�Z:��d夿@5���.ڿ���P������߰���v���ۿ��¿S��%F��L�U�U��Y�⾨ŗ�V�>�2p�����XC�^Yd�% ������   �   �����_�˕��u�о�a�'����4�LtG��uS�+�W�T�ŕH�Y6�t�0���:Ӿ�S���b�F|��A��r[Y�hv��d?������/�{�'žC)��#J�����W�̿�����N�����F��>�������/[οf	��WZ����J�W�žR�z����!S��f�<�����U�Oڴ��   �   z��c����D�)���Jʬ�TҾz�������B��t����Pp���Ծm���?���VG�������a5�wμx�Ӽ`~J��cͽ+�<�Z���0���P�2��`v�uġ��)˿'S��\�D�!�r�0�
;���>�n�;��1�ֻ"��������˿����qv�BE2���������V;�w?˽4�F�P ͼ�oǼ�1��   �   ��D�~�7ֽ���@�Q�����R̙��>��x9������ĸ��:���������i*T�\�P�ٽ	O��lu��p{#��˛��㕼,a�����	�c���v���R��S��'f�����40��B&�:�<���O��\�fsa�<]���P�Ƽ=�� '�N��U���=��
���:�Q� ���ϻ���a�:��fl\�dm�� 8������   �   ��;(�X���(��B��}������3��M�K{]�fc��1^�2ZN�g5�����4但H��2�-�`;i�`g�;�#s<�<*j�H�|��������Iپ�0&�o��좿��ӿ�D����l�;���V�@�m� �}��ǁ��+~�r{n�MW��<�������ӿ���9�m��$��m׾�T��^	�<w�X�Y�P�(<p�<�   �   x�<���< ��:9��>�?��4��4C��� �� ���9�{��_�你z�����UD����� Z�9�P�<h�<�� =���<(XM�����,��	�� ��>�6�Ͳ��
���5濊��3.�.�M���l��ۃ��$�������F��n����l��M�X�-� ���俍-��^�����4�$Y�[�����������;�f�<��=�   �   �:9=�U=���<�<��3�����v�@���w����1"��u��"ez���C�����h�A��W�;���<��=��6=�'=|d�<��C������)�$]��;���@�j։�<ͺ��� /���7���Y�~�{�o���o�������%���Fx{�N,Y��6��� ���Є��?�cs��Mu��,Q'�����u1����<ܡ*=�   �   �\$=8�=�&�<`��;h'S��� ���D��iz�:\��/H���W��Dz�D�ر���I��H�;���<��=��(=V
=�M{<P�̼W�����I�ِ��F���Z�<���_�пF���)�hO��ux�����8���z��,ʳ�Nu��!��>ΐ�6�w� �M���'�6��0Ͽ?����X����/o����H�^��\�м��m<��=�   �   (=�!�<�g<�:��( Ѽ|�<�܃��|�� |�� ��ǈ���u��%����u;�,ͼ�+��x�u<$_�<�S=XJ=�g^<�μ����E�!���0�$+V����u?Ϳ���+&�*8K��cs��������Nt��ӯ��fz��v��|���ԩr��HJ��3%����4�˿z	����T�Z>�����2�D��깽��Ѽ�Q<�5 =�   �   K�< m�;�J�!��.���ɺ���� 	����������I	����^ƺ�e����F�`�?���<�ɪ<���<��<TpӼ�\���:��إ��H���J�\���-ÿ9�������U@��!e��������� ��;����!���#��I�����d�\�?��<��L���¿&����I�Nz�r뤾�H9��@���׼�*�;4��<�   �   �3ֻ��漜 p�?�������=/��Q��mm��0�����͈���m���R�'�/����V���v�n����Ϳ� �;�M��,f�|t��n(�+���	���9��?��0i��K���1��0��%P�^�o�����A���~���A��v��vBp��lP���/������翎���֩���8�|���s��m�'�<m��К�`g(��pP;�   �   ��;�����r���<9��r��Õ�����:þe?о%�Ծ��о��þhί��r���t��9����Ħ��/:����|���г�������E����4վ,�"��i��E��i(Ͽ�`��C�\e7��JQ��pg�P�v�VX|��Dw�6Zh�@4R��8�l��<z�(Ͽi����h��!��gԾ�1��������B����������   �   �̽�� e�7@��_ľ��~���M�ʮ ��$�r� ����Vp	�sN<ž���^f��i�ų̽F�w���"�6�%�7l��[(���Z�m沾O8	�ؤF�PW��_K���O߿D��TL�B$2��|C�@?O�`�S�<�O�.oD�T)3�J'�XL���߿����w^��2xF�u��px��HZ�����w�� e&���#�^x��   �   �/��*��p����l�n0�ޒI���]��j�$co��9k���^��J�%%1��[��J�j��l�����/�������V�\����ϽD 0�����rS޾�@"�R�`��铿?���6��R�8���!��*�X	.�.3+��"����+��⿨���c��ca�b"��G޾\ʏ�|�/���ν�����A]���������   �   �������� ���9)�)Q��w�1׌��<���ޢ�����P?��皿O����By��R��L*��n�F������Ђ0����X����Ą�����l���]��A������f1���k������ҵ���Կ���L����	��@�
��Q�CO�-ֿD ���h����l�r�1��n��t����]�����㫽��-����Rཐ0��   �   /c�����l�3�dUf����Х����_�̿��׿��ۿ/gؿ��Ϳ�ż�������g�v�4�=z�(����q~��m"�,\ͽkʒ�a̒��NͽA"��}�{^��o����3��Pf��
���̥�������̿��׿��ۿ�cؿ_�Ϳ�¼�������+�g���4�x� ����m~�Vk"�LZͽ˒��ϒ��Tͽ�E"���}��   �   ����i1�4�k�Q����յ�g�ԿF��L����	��B�
�lS��R��ֿ���yj����l���1��q��Qv��}�]����㫽-���M����J��0�Ґ����Ю��5)�P$Q���w�<Ԍ��9���ۢ�����4<��#䚿�����=y�.�R��I*�ll������	��g0���1����ń��������]��E���   �   �C"�"�`�-쓿�A��2:῔T�@�0�!�Z�*��.�Z5+��"�@�8-�|�⿛��Re���a��c"��I޾�ˏ�μ/���νԎ��,:]�j�����i/��&���j�����)h��0���I�P�]���j��]o��4k��^���J�H!1��X�iE�f��c���a�/�X��H�����\�����Ͻ>0����W޾�   �   �F�EY���M���R߿��@N�p&2�"C��AO��S���O�DqD�+3��(�~M�w�߿a����_���yF�~���y���Z�h����v���^&���#��Ox��̽�����d�.;��`ľ��쾫��yI��� ��$�T� �&���l	�cH7ž��� f�e�-�̽�w��"�%��n���-��^�Z��鲾�:	��   �   �i��G���*Ͽb��E�Lg7��LQ�fsg���v��Z|�Gw�R\h��5R�*8�p��{�WϿJ���M i���!��hԾ>2��"�����j��4w�������;��^��459�<�r�����-���4þ#9о��Ծ��о��þGɯ�~n��Ft��9�(�������%:�d��T���~��s�����t����7վp�"��   �   �@���j��a��.3�
0�|'P���o�֎���������B��j���Cp��mP�� 0�������%���>���m 8���t��Q�'�"l��Ȓ漠(���P;��ջh��n�o������|��6/�b�Q�Jem�&(�Y���|����m���R��/���������n�tl�P���@�;�<��4k㼎w���p(�4-������9��   �   ,]��C/ÿ�������V@�X#e�����������1���h"���$������B�d���?�
=�MM���¿E���/�I�Lz�J뤾\H9��?���׼ O�;䲬<�Y�<���;@�J����&�����܉��	�5~�V��j��SD	�`��ྺ�!����<� �?� �<�Ъ<l��<�<LvӼ�_�� :�pڥ��I���J��   �   g���@Ϳ���f,&�9K��ds�9��:����t��W����z��[v��������r��HJ��3%�����˿G	����T�>���4�D�鹽��Ѽ�"Q<�9 =�	=,�< ,g<��Ѽ��<�/׃��w���v��������}q��5���Fo;�ͼ�	���u<�b�<�T=J=�`^<(
μt��&�E��	���1��,V��   �   �����п���V)��O�vx�����8���z��,ʳ�8u�����ΐ���w���M�<�'����x/Ͽ���� �X����%n��B�H��[����мإm<��=x^$=Ԡ=�)�<`��;0"S�t� ���D��hz��[��$H���W���z��D�������I��>�;���<t�=�(=P=�C{<$�̼����r�I������Z��   �   ����?Ϳ,���+&�8K��cs�m��K����s��N����y��pu��㵍�ƨr��GJ��2%�,��.�˿�����T�Q=� ���D�~繽��Ѽ(Q<�: ="
=�,�<�,g<���Ѽ��<�7׃��w�� w��������{q��7���<o;�ͼP����u<�c�<,U=�J=Hf^<μ����E���� 1��+V��   �   �[���-ÿԑ��2��4U@�!e�i����������G���� ��#��d����d��?��;�@K��M¿���Q�I��x��餾F9��<�� ׼ c�;赬<�[�<��;8�J����&��������	�>~�]��t��XD	�a��ܾ�����n<���?�X�<�Ҫ<���<�<|nӼ�\���:��إ��H���J��   �   2?���h��s��X1��0��$P�ޭo�����!���}���@��C��R@p��jP�`�/�������⸲�����8�f��q���'��g���� �'� Q;��ջ���o������|��6/�j�Q�Sem�5(�^��������m���R��/���������n��j⼐�����; ���d`�Ws��~m(��*�����9��   �   ��i��D��9'Ͽ�_��B�d7�IQ��ng��v��U|��Aw��Wh�2R��8�Ξ��x��Ͽ�����h���!�udԾT/��F����� ��o������p�;��F��)59�<�r�����4���4þ,9о��Ծ��о��þJɯ�~n��<t���9���8���R$:�  �������q�����~����3վP�"��   �   H�F�>V���I���M߿ ���J��"2��zC��<O���S���O��lD�*'3�f%��J���߿�����\��&uF�'��u��>Z����q���W&�>�#�Mx�N�̽]����d�);��^ľ��쾭��}I��� ��$�Z� �'���l	�aH7ž����f��d�F�̽@�w�r�"���%�Si��,%���Z��䲾97	��   �   $?"���`�K蓿%=���4�RQ����!��*�.��0+��"����)��}����qa����`�_"�C޾Ǐ�|�/���νV���3]�2���$��/��&���j��|��)h��0���I�T�]���j��]o��4k��^���J�F!1��X�^E�f��C�����/�������b�\�����IϽ��/��Q޾�   �   H����c1���k������е�3�ԿW�ￄ����	��>�
��O��K��ֿ4����e��Q�l���1�i���o����]��}��۫�����H�F0�����k�̮��5)�Q$Q���w�?Ԍ��9���ۢ�����6<��%䚿�����=y�+�R��I*�dl�t����	���~0��}��񖽙����������]��?���   �   U[��H����3�Mf����jʥ�������̿r�׿G�ۿ�_ؿʵͿ^����ꦿ���h�g���4��t�H�)f~��e"�OQͽ!Ò��ǒ��Kͽ@"���}�V^��f��~�3��Pf��
�� ͥ�������̿��׿��ۿ�cؿb�Ϳ�¼�������*�g���4�x������l~�aj"�BWͽMƒ�BȒ�Jͽ�="���}��   �   ����￾V��m2)�r Q���w��ь��6���آ����8��ᚿ����{8y�f�R��E*�i�B������y0�v��얽5���������L�]��A������f1���k������ҵ���Կ���N����	��@�
��Q�EO�.ֿB ���h����l�j�1�jn���s���]�f���߫�<�����"E��0��   �   �/��#���f��J���d�-
0���I���]�{�j�lXo�X/k��^���J��1��T��>�<a�������/����������\������Ͻ2�/�D���IS޾�@"�O�`��铿?���6��R�:��!��*�X	.�03+��"����+��⿧���c��^a�b"�XG޾ʏ�k�/�:�νN���B2]�o���Ѝ��   �   ކ̽���j�d�7��Zľ���?���E�}� �l�#�� ���i	�wA1ž�����e�X^���̽�|w���"���%��g���%��@�Z�0沾A8	�ҤF�PW��`K���O߿F��VL�D$2��|C�D?O�b�S�>�O�.oD�T)3�J'�XL���߿􎲿v^��*xF�g��5x��vZ�9����s���X&���#�Ex��   �   �;��禽���0/9���r�7���%��-/þ&3о��Ծm�о��þ�ï�ni��kt���9���������:�,꼼����&��O����������4վ$�"��i��E��j(Ͽ�`��C�^e7��JQ��pg�P�v�VX|��Dw�6Zh�@4R��8�j��<z�(Ͽi���
�h��!��gԾy1�����㖓����<k�������   �   �ջ\��\�o������w��0/���Q��]m�������w���m��{R��/����x����n�8O⼠9���I�;���8X�(r��Zm(��*��{	���9��?��1i��M���1��0��%P�`�o�����A���~���A��w��vBp��lP���/������翏���֩���8�a��s����'��j���漠�'��JQ;�   �   �b�<���;�rJ��	�� ������z��Q	�7y�"��1��>?	����$���^���(/��?�<8�<X
�<��<,gӼb[��:�tإ��H���J�\���-ÿ:�������U@��!e��������� ��;����!���#��I�����d�\�?��<��L���¿&����I�Gz�S뤾kH9�|?��׼P]�;���<�   �   �
=T0�<�8g<P����Ѽ �<�jӃ��s��Rr��'���~���l�������f;�<�̼т��u<n�<�Y=�N=Pt^<<�ͼ ��ݺE����0�%+V����v?Ϳ���+&�*8K��cs��������Mt��ү��fz��v��|���ԩr��HJ��3%����5�˿z	����T�V>�w�����D�깽$�Ѽ8!Q<": =�   �   �k=l_�<P�j< �Y�Լ��:.��Uu���`���M���§�U��6dq���(�|����'���=�<�W�<\�=0B�<p��;���H'ٽZ�]�Q¾ b��h�t��C>ݿ|����3�M]�����������W������^T��T���*ޜ�n��|�\�\�2��f�[ܿZף���g���z���]L^���۽���@��;�b�<�   �   ��<�j�<�ݫ;p�m���Um��������ϯнN׽$н�Ż��%��hEh��� 3P� ��;���<�<d`�<@��;�:�	սn[Y�EY������d�L���F�ٿj���0�tY�O�����^�����<���	��?����g�������{X���/�6�n�ؿ�����c�J+��@��bZ�ؽ�6���w;Ӿ<�   �   ��9< YǺ����r�H�ힽumؽg��6��'��{+�:�&����v��Kֽ+��
B�P��� ��9�[<��n< HZ��!�FE˽vM�����{+�؎X�c���Ͽ�����'�t-M��v�D����y��N������S�����������f�u���L��:'�x��pοS����W���Ώ��(�M���ͽ�������H�M<�   �   5��� !��M��i���� �B��}g�L<��ϊ������e����!���g��2B�f����ݽW"�� �`_p�����8-����}���{:����Z<�l�E��݌�e����������o;���^������R���ۚ�������������-��6�^��j;�:���:��k)������zE�N����z(;�+���� ��4I�`�̻�   �   ,.m���ý@��z�M��o���_��o*���hӾ%�i���&ᾭ�Ӿ?7���N��5����L�������f��r�\)ܼ��-��
����#�=}��H�徏(.��Ly��l��^�ۿ�K	�"&���C�<4`���x����#�������oy���`��D�^U&��[	���ۿ�E�� �x�$�-�-�徫���2�$����r�2��K�����   �   '��|�1��|�%8��!�ԾR����Q���"��w,��/�`�,�3�"����l& ���Ծl(����{�5�0�kC�q�NN�|Q��P���D���o������z��|T��V��1���}%��FR'�f�=�*�P���]���b�:^��Q�`�>���'�*o�È�ｽ��Z��:hT��d������p���������U�-S�mo���   �   l�B�������¾����߬�$�<��W�D#m��z����,�z���m��iX��s=�*� .��þ�c��;B�m���s騽����<���7���B�����h��L.��p�k����ƿ�K￈���v�P,�x�5�H>9�(6�F�,���$
����ƿj睿@p��'.���ﾢ�����B����l�����]���=8 ��   �   �'���(о.����5��	`�RW��QE��4W��5[�����m����������,���Y�`��66�'��Fо�	���1C����u�!ѝ��aǽPD��Us�����B>�(|��z������}�� ���.�
�J.�����j�^+�n���v��0¿�ȓ|�	�>�������Cs�>E���ǽ8|��>籽&�����C��   �   G;�B�A�Vcv�z���d���B�ǿ�ٿt8�OS鿭���1ڿ_Dȿ�E���
���w��iA��q��Y;v늾�y4����߬�f��A�X�4�����B;j?���@�R^v����������ǿE�ٿ�4�qO��忁.ڿ9Aȿ�B��E���w��fA��o��V;S銾jw4���꽬߬������L�4�� ���   �   ����F>��|�p}��ɇ������N�
�|0�*���l�L-�۫��l�⿒2¿���|�|�>��������Fs��F��ǽ�y�� ⱽ�����C�~#��2#о���n�5��`�xT��2B���S���W������)�������K�������5�`��36�`$��Bо"��`.C����7�vҝ��eǽH�L[s�?����   �   j.��p�秝��ƿO�|���x��,���5��@9��6�b�,�����p���ƿ靿vBp�Z).�S�������B���Tj��	�������l3 ���B�'�����¾�������p�<���W��m�j�z����z�Z�m�eX��o=�� ��(����¾�`���B�����j樽���>���<���B����� ���   �   �T��X������{(���TT'���=���P���]�ȓb��<^�R�Q�J�>�n�'�fp����o���\���iT��e����p���<�����U��"S��g��ш뽪�1�.|��2����Ծ����M���"�#s,���/��,�#�"����8# ���Ծ$��Ā{�4�0�m<�ꓽ�JN��|Q��S��>G�L�o����L}��   �   �Oy��n����ۿ.M	��&�ТC��6`���x�6������3��ry���`��D�zV&�f\	���ۿuF��T�x��-�=��/���`�$���p�2��;�j���m�X�ý�����M�@k��PZ��w$��3bӾ�����} ᾩ{Ӿ�1���I��#1��7�L������b�f��l� %ܼt�-������#��������*.��   �   ,ߌ�2���'�����q;���^�(���T��=ݚ�U����������u.��r�^��k;����g;��*�������zE������^(;� ��ȳ ��I�pU̻���"!�yD��(^�P����B��ug��7��@���p����|�����H
g�X,B�����ݽ�����@Dp� ���x-���������}:�%���=���E��   �   �����Ͽ�����'��.M��v�J���{��l������A�������&���6�u�z�L�;'�Fx��pοu����W���������M�Q�ͽ���@X����M<�:<�$ƺ����d�H��䞽%dؽL����T'�v+���&�������Cֽa$��d�A��r�� ��9��[<��n< ]��$�oH˽	M������,���X��   �   7���d�ٿ����0�vY�������������ɑ��|�������g������{X���/�"�=�ؿy����c��*�/@��UZ�-ؽb3��x;,۾<P%�<�u�<��;��m����Lm�������]�н�H׽н����!��L>h�<��� P� ��;���<��<�_�<@�;>�߁ս�]Y��Z�����#�d��   �   �t���>ݿ����3��M]�仅�C��!��X������FT��%����ݜ��m���\���2��f�rZܿ�֣���g�>�_����J^�n�۽t�����;g�<�m=�b�<��j<��Y�HѼ��9.��Tu�����S`���M��ç�GU���dq���(������P��;�<hT�<��=�=�<0��;2���)ٽ�]�v¾�b���h��   �   ����z�ٿ~����0�fY�6��܈�����������h�������f��e����zX���/���X�ؿ���~�c�0*�0?��Z�~ؽ61� x;�ܾ<X&�<Dv�<��;`�m����Lm�������f�н�H׽н%����!��F>h�6��h P�@��;P��<�<�a�<`�;�;�-�սL\Y��Y��B���d��   �   C����Ͽ���>�'��,M�$v�����#y��a������9���ݑ��������u���L��9'�.w�2oο!����W��������'�M��ͽ�������M<x:<�ƺp���>�H��䞽+dؽQ����\'�v+���&�������CֽW$��6�A�8r�� @�9��[<8 o< �R�� �=E˽�M�����z+���X��   �   O݌�Ŋ�����&�o;�r�^�����Q���ښ�����=��9���l,��8�^�<i;����_8���'��'����wE���!���$;����� � ��I��C̻���V!�BD��^�J����B��ug��7��G���u���}�����O
g�Y,B������ݽI��<���>p�0|��@-����H���fz:����<���E��   �   TKy��k���ۿ�J	�&�:�C�X2`�|�x�[������Y���ly�,�`�nD��S&�"Z	�H�ۿ�C����x���-�������M�$�>����2�3����m���ý�����M�?k��SZ��|$��<bӾ����徇 ᾰ{Ӿ�1���I�� 1��*�L����1����f� j�|ܼ��-������#�m|���徨'.��   �   �zT��U�������#����P'���=���P� �]�6�b�@7^�d�Q��>���'�lm�ͅ�r����X��eT�,b����Wp������`�U�S�wf�����o�1�|��2����Ծ����M���"�)s,���/��,�&�"���8# ���Ծ	$����{���0��;齭蓽FN�BuQ��M���B���o�	����y��   �   �.�mp�ϣ���ƿI����t�8
,�&�5��;9��	6��,��
�2���ƿ�䝿�;p�q$.�7��#���K�B�,�콍d��T���n����2 �Z�B�	�����¾�������r�<���W��m�p�z����z�`�m�eX��o=�� ��(����¾�`��JB�<���䨽e���9���3�G�B�ݼ������   �   @���@>��|��x�������῿���H�
�:,�����h�B)�y�������,¿#쟿"�|�J�>����R�N=s�2@��ǽ9t���ޱ������C�O#��#о���k�5��`�yT��5B���S���W������,�������L�������5�`��36�[$�Bо����-C�ۍ���창͝�]]ǽ�A��Qs����   �   �>;#=���@��Zv�>���d�����ǿؚٿ�0忙K��忽*ڿ�=ȿ�?��Y���w��bA�=l�hQ;t劾�q4�B��^׬�d ��
�]�4������A;`?���@�R^v����� �����ǿI�ٿ�4�tO���必.ڿ;Aȿ�B��E���w��fA��o�]V;銾rv4���꽻ڬ��� ��4������   �   � ��8о���5�� `�R��u?���P���T��]���ɉ��d���-���㺄�-�`�I/6�� ��<о����'C������簽|ʝ�K]ǽ�B��Ts��ﺾ����B>�&|��z���������"���0�
�L.�����j�`+�p���w��0¿�Ɠ|� �>����v�
Cs��C�@�ǽ�u��eݱ�̜��V�C��   �   ��B�݉����¾"���Z��g�<�L�W��m���z�gy�	�z�݃m��_X��j=�����!���¾(\���B������ݨ�Q���&7��4콩�B�I���<��B.��p�k����ƿ�Kￊ���v�R,�z�5�H>9�*6�F�,���$
����ƿi睿�?p��'.����Q���x�B��콤f��ꈇ������/ ��   �   '�뽁�1�a|�v.��m�Ծ����J���"��n,�'�/���,���"�ց�� �0�Ծ����w{�$�0�B1�ᓽ�;N��nQ��L��C���o�]����z��|T��V��1���%��FR'�j�=�,�P���]���b�
:^��Q�`�>���'�,o�ň�ｽ��Z��3hT��d�w����p�b��)����U�.S�?b���   �   m���ý���7�M�Tg���U����G\Ӿ*�2����OuӾ�+��tD��v,��M�L������0�f��^�\ܼ��-�a����#��|���徆(.��Ly��l��`�ۿ�K	�$&���C�>4`���x����#�������oy���`��D�`U&��[	���ۿ�E����x��-���^���(�$�C��n�2��.�����   �   ���z!��=��dU����^�B�{ng��3��運�񵎾~x��9��*g��$B�~���ݽE������p��7��H�,�������Ez:����L<�h�E��݌�e����������o;���^������R���ۚ�������������-��8�^��j;�:���:��l)������zE�@�N���';�����Ұ ��I��'̻�   �   �+:<@ZźXp����H�Nޞ�j\ؽ�����	'��p+�K�&�C�����:ֽ:��J�A��Z�� �9��[<�o< P?�
��C˽�M�y���t+�ՎX�d���Ͽ�����'�v-M��v�E����y��N������U�����������h�u���L��:'�x��pοS����W� ��������M�3�ͽ�����H�M<�   �   �'�<8z�<@+�;؞m�����Em������q�н�C׽�н�����5h���XP��;,	�<H�<xi�<��;@8�C~ս4[Y�6Y�������d�K���E�ٿl���0�vY�P�����^�����=���	��>����g�������{X���/�4�m�ؿ�����c�F+��@��*Z�Fؽ�4���w;ܾ<�   �   ԣ�<�M�<�#<����@�d�H�5���9������p���Hʵ�����W���y@�\-ۼ �ϻTB<�a�<��<C�<@�@;�I%�݀��Dg���Ⱦ ��n������~�0\��8�d|c�����[��K(�������s��g����%���T�����hfc��8��S�������;o��r ���ɾ5�i�^��l�0� �%�(�<�   �   ���<(!t< ����3��"�/�b̈́�-ଽ�R̽7:ཞ��e߽b	ʽv���7�����%�0����5';8�<��<@ά< ƈ:��%�x��}�b�>�ľ����j�$�����޿X��:�4�t"_����r���Y����c��_���d�������������<_���4�F����޿`ԥ�:k�ց��ž�He��齂L1�@*��|�<�   �   `!�;/�l���d�M4����
���@#�\0�ٰ4�h�/�~$"������0]��<�Y�p�ռ ��(�< =$<p���&�(��hٽpV�:����J�^������ Կf	�8�+���R��}�Ub����A���|
��᧳�K���c��t�}���R���+��	��&Կߛ���^�y��6�����X��e޽p�3�0�����;�   �   3��RY<�x���l�y#�VM�ʸr�<!��(���c����K��n���k0q��aK�,!�>I콡�����0��X���i�`%��,�1���ʽ�{C�)���o���K�Š��%]ÿ�������H�@�Bue��,���=���5����<���F��4��F|e���@���������dÿ|�����K� ��6 ��
zE�Ͻ�;������)F��   �   <��9EԽta�܋X�`���J��X�ž�[۾}9�������<�ھF�ľ_c��ܐ���+V����`
Ͻ��T+��\�VE�D����,��0��ֳ�n3�l#���筿������p�*�,>I�$g��o���B��nj��J���z���/g��KI���*�l��|��t��0����3�9:����6.�6����N�|���K'��   �   ����@�;����?W����ܾ0��j��(�] 2�g5��1�i�'����<��۾H��4񂾜�9�j(��e����f�j�`ޭ�kk�Mez�Z�Ⱦ�:�`�Z�e����¿/h����<�+�*rC��0W���d��Ki�,�d�0DW�\�C��,�~��k�[�¿�d����Z��T��ɾlc{������Fcq���n��s���   �   �BM��󓾫�ʾ��B&$�y3C�&�^�Ut�����i������+t��y^�_�B�2�#�����ɾ�����UK��"�ũ�����bЧ�ݻ���vL�s���@����3��(w�����˿����S�&�!�~�0�~�:��?>�$�:���0��!�^[������˿q��!w���3��B���&���M�m�����/ܕ��鹽���   �   Ő��g5ؾ�����;��"g��]������ �����G=��k��������	@��H�f��w;�4���l׾�ϗ��L��3��������sKֽ�"�b~�!¾�z��RD�vҁ�e��C�ƿ�<�r���}���h���
���.���=迪�ƿ�������b&D�_T������0~�( "��׽w���k���,_���M��   �   ,վ-C�wBG���}�����󶵿,ͿɈ߿B뿸JￗB�J�߿�$Ϳ����c皿�}��F�O���Ծ����8�=��a��"M��b����6��h>����վ�?�8>G���}���������k(Ϳ�߿>��F��>뿽�߿�!Ϳ�����䚿��}��F����ǐԾY�����=��_���M������N=�� m>�{���   �   �}��VD��ԁ�>����ƿQ@�|������������������@�7�ƿ�	�������(D�+V�8����3~�|!"��׽����2����Z�o�M������/ؾ����;��g��Z��������������9������#����=���f�8t;�����h׾�̗�^�L��1�n��P����Oֽ"��g~��%¾�   �   Т3��,w������˿m���U�f�!���0��:�|B>���:�(�0���!��\�u�����˿���w�T�3�'E��u(�� M��m����ؕ��⹽��<M�E�ʾ6�	"$��.C�ײ^�lOt�����f�����|&t��t^�4�B���#���u�ɾ;����PK���������vҧ�����;{L�����E���   �   ��Z�%g��A�¿?k����\�+��tC�P3W���d��Ni��d��FW�Z�C�T,����m��¿f��J�Z��U�'ɾ�d{�P��V���\q�N�n�l��6���D�;�����Q��g�ܾo���e�8(���1�tb5��1�A�'���Z9���۾�C���킾z�9�G!���	��ƽf��j�᭽4n��iz�ѿȾ6=��   �   %���魿n��D��>�*�^@I��g�4q���D���k���K���{���1g�DMI���*�H��Ȑ�j�1��q�3�S;�0ᔾ7.�����N�H���?'�<����:Խ�Z�ɃX������D��8�ž�T۾�2���K���ھ��ľ�^��͌��%V�����Ͻ���(%�|Z��WE�_�����,�:3��Q��p3��   �   =����^ÿ��� ����@�\we��-��3?��f7��r��h=���G���4���}e���@�\������+eÿ�7�K�O��s ���yE��Ͻ֬;��{�� F����vJ<��n��Za��r#��NM�c�r����}�������G��5����(q��ZK�v&!�=@콟�N�0��J���Z�$��ֹ1�=�ʽp~C�@+��>q�;�K��   �   ����7"ԿT	�^�+�>�R���}�fc��:��g������ר����kd��P�}�F�R� �+��	�1'Կ���-�^�v�����(�X��d޽��3� ���@��;�`�; ��@�케�d��+�����͟�F;#�JV0��4���/�S"�4����kV��D�Y���ռ�Ў�p�<�C$<p���j�(�lٽ�rV�:�����;�^��   �   �����޿���4�|#_�\��&��� ���d�����Pe�����>�������L_���4�4����޿+ԥ��
k�v����ž�Ge���H1�@������<`�<x7t< R��`$����/��Ȅ��ڬ�M̽�4�$��/߽�ʽ3���������%��@l';��<�!�<�ͬ<���:�%�U�㽵�b���ľ�|�j��   �   A����⿔\�B8��|c�E���[��{(�������s��O���Z%���T��^���ec�B8�^S�o��t���;o��q ���ɾ��i������0� ����<���<HQ�<*<����=�,�H������������^���`ʵ����kW���z@��/ۼ@�ϻXNB<p^�<\�<�>�<�n@;HM%�J�罃Fg��Ⱦ� ��n��   �   ^�����޿l��D�4�f"_����<�������c�����3d������S������8_���4������޿tӥ��	k������ž�Fe�P齼F1� ���|��<\�<�8t< 9��8$��r�/��Ȅ��ڬ�*M̽�4�.��7߽�ʽ7���������%���n';,�<�"�<\Ϭ<���:��%����`�b���ľE�l�j��   �   a���q Կ0	���+�>�R�6�}��a��G��L���k	������&���b����}�H�R���+��	�m%Կ����%�^��������X�Ba޽t�3�����p�;�h�;����P�d��+�����ҟ�N;#�TV0�#�4���/�^"�>����`V��*�Y���ռ@̎�8�<�I$<p���>�(��hٽ$pV�J����4�^��   �   W����\ÿѸ����^�@��se��+���<���4������:��=E���2��.ze��@�\��l����bÿ���g�K�T������lvE�]Ͻ�;�\t����E����I<��n��:a��r#��NM�k�r������������G��=����(q� [K�v&!�)@�k񛽌�0�,H��XQ�����1�ʽ�zC��(��Bo�k�K��   �   �"���歿������L�*��<I�(g�n���A���h���H��%y�� -g��II�ʒ*������s뭿C/���3��6�ޔ��2.������N����='�l���R:Խ�Z���X������D��?�ž�T۾�2���V���ھ��ľ�^��̌��%V����bϽ��|"�,V�QE����ʇ,�0�����/m3��   �   ��Z��c��-�¿9f�����+�2pC�..W��d��Hi�D�d�rAW��C���+����h�Ш¿�b��R�Z�/R�ɾ�]{�α�z���NUq���n��j��X����;�z���Q��d�ܾp���e�<(���1�zb5��1�F�'���\9���۾�C���킾B�9�q ������f�j�Gۭ��i�cz���Ⱦ�9��   �   ʝ3�.&w�`��q�˿Y���tQ�H�!�T�0��:�\=>���:���0���!�`Y�a����˿���w�N�3��=��a#��F�L�zd��(��?ԕ��๽Z���;M�&дʾ2�"$��.C�ڲ^�pOt�����f������&t��t^�6�B���#�
��g�ɾ����PK���Z���`���̧�׷��btL����Z>���   �   y�3PD��Ё�Q����ƿ�9迶���{�b�,��~����(��5:�d�ƿ��������"D�hQ�V����)~�"�?�ֽU﬽�����Y���M�P����/ؾ���;��g��Z��������������9������&����=���f�6t;�|��vh׾�̗���L��0����Ŧ��Gֽ
"�^^~��¾�   �   �վz=�#;G���}�G���Ͱ��=%Ϳe�߿P:��B��:��߿Ϳ]���⚿޳}���F������Ծc�����=�BV��LE��D����3��g>�~���վ�?�2>G���}���������n(Ϳ�߿>��F��>���߿�!Ϳ����嚿��}��F������Ծ�����=��\���H�������1���d>�X���   �   �����+ؾY���;��g�iX����������6��f6�����-������:����f��o;����b׾zȗ���L��,����,���GֽM"�0a~�A!¾�z��RD�tҁ�d��C�ƿ�<�t���}���j���
���0���=迫�ƿ�������]&D�PT������/~��"�� ׽��\����W��M��   �   7M��듾k�ʾ^��$��*C��^�6Jt�	���c������� t�yo^�j�B�y�#�~����ɾ��IK�������5	���ʧ�2����uL����@����3��(w�����˿����S�&�!���0���:��?>�&�:���0��!�^[������˿r��w�z�3��B���&���M��i��I���ӕ��ݹ�v���   �   [�����;���NM����ܾ/��:b��'�]�1��]5�~�1���'����5��۾>��A邾H�9����� ����f��	j��٭��i�hdz��Ⱦ�:�Y�Z�e����¿0h����>�+�,rC��0W���d��Ki�0�d�0DW�^�C��,����k�]�¿�d����Z��T��ɾ�b{����8����Uq���n�=f���   �   T����2Խ�U�:}X������?����ž�N۾.,�Z���辗�ھ��ľY������V�����ν4|����M��KE�չ���,��0�����n3�k#���筿������p�*�.>I�$g��o���B��nj��J���z���/g��KI���*�l����u��0����3�:�Y����5.�̢���N����7'��   �   ����?<��g��XX�xm#��GM��r����������|B��Ñ��� q�zSK��!��4�;蛽��0�@1���.� ��¯1���ʽ�zC��(���o���K�Ġ��&]ÿ�������H�@�@ue��,���=���5����<���F��4��H|e���@���������dÿ}�����K����  ��LyE��Ͻ��;�Hs��@�E��   �   @��;P���켐�d�:%�����@��:6#��P0�v�4�6�/��"������N����Y�uռ�}����<�b$<�b��d�(�Cgٽ�oV�����H�^����� Կf	�8�+���R��}�Ub����A���}
��৳�K���c��t�}���R���+��	��&Կ�����^�q�����9�X�od޽��3�������;�   �   
�<�@t< ���<���|/�ń��֬��H̽�/�ҧ��߽L�ɽ(���勀�,�%��ߑ� �'; �<�+�<�׬<�2�:F�%����B�b�.�ľ����j�$�����޿X��:�4�t"_����s���Y����c��`���d�������������>_���4�F����޿aԥ�9k�Ձ�p�ž�He�(�4J1��������<�   �   �_�<�e�<��;0x6�8�����O�H���즧�.1��1���Ҁ��Nf������_D�8)��:���)+<���<L!�<�߽<@��:��(�ہ�r�e��Ǿ�v�sl��Ʀ���
��"�5���`����������U�����������4��D��
(a���6��J������?�m�8���Fɾj�}��f8���`&�<�   �   `�<`.O<��#��R��,�6���������Փν4⽴3�}Z�gF˽�窽�,��(z)�lI�� ݡ: �<���<Ĭ�< �o��K)�����a�Uþ����Uh����tܿ6h���2�<Y\�1��U~������IĽ��X���������E����b����\�tc3�D���YݿǤ�U�i�~���yž�e���뽶�8��,�� >�<�   �   ��p;X��D���6�k�W&��0L�Ƅ�!�#�(�0�L�4���/��"��$O��W��x�\� �ݼ�L���q�;x�<ɻPn,��ٽ_U�_����;��_\��웿+�ѿJ���)��eP��lz��n��UӤ�2��$����!��*����j��&�z�ЮP�2Y*�`�*�ҿ���Ƈ]�IH������Y�iὌ1;� � ��;�   �   �JɼD�C�����a�� U$�,�M�o�r�뇾�)���.�����$���p�͘J��� �lb��뜽�X4�8<��8@-����Q5��+˽[�B�Q����C�Y�I��;��B{��	L��q���>��b������]��x��Nܡ�f����1��os����b�"�>����M�����������.�J���b���� F�?�ѽ��B�p����~g��   �   NT����ֽ�W�Y����KžD`ھ��羾v� h羷Oپ��þ2�������U�>s�TsϽ$#��:!�`����H�q���~',��R�����M�1�s�}��X����߿Ԗ�Z)�\VG�"�d�X~�-���R���u���}��Cd���F���(�`��m�߿T����~�=x2�E�H���*�.��S���T��]� �.��   �   ���i�<�R����J%ܾ��r��L'���0�s4��t0��`&������ھ�򬾷 ��X�8�@��o4���5j�"�m�>!���n��Yy�PnǾ����X��)�����|�b���*�|�A�� U��b�j�f���a�L�T��3A�*�j��������$���'Y��Y�)1Ⱦ�#{�/u�Z�����w�pcu��`���   �   %�M�I̓��"ʾ+���U#�WB��V]�Ъr����W������q��T\�J�@��/"�8p�!Ⱦ%��B�J�/�ַ�ʹ���Z��b����L�y<��ר���S2��Ou�蠿Uʿ{���J��� ��\/�.	9�2S<���8�n�.�, �6���E��ɿ4���|�t��-2�����<���JM��������@���(y��u�	��   �   �G���h׾P8���:���e�����t���Ḩ�����jy���Q��?���ۆ��~d���9�z5�ٷվh喾<�K��l�f���^f����׽ G"���}�:7�����qC�����H�ſ�������i�����>���	��v������Ŀ�a�����MkB��>�z����t}��l"�2�ؽ�G��4ýA.	��4N��   �   �1Ծ,u�`F��i|�S��F�����˿u�ݿ�d鿣7���JNݿ�˿³��L���.{�ZE���(Ӿ���=��o��������������>������,Ծ�q�)F��d|�\���6�˿��ݿ�`鿶3�
��Jݿ�˿P���1J��+{�KE�����
Ӿx�����=�vm��! ��Q���������>��Ð��   �   h��9C�b�� ����ſO�����l�����@�:���
��x����p�Ŀ�c��,����mB�O@������w}��m"�8�ؽ{E���.ý*	��.N��C��Pc׾�4�9�:���e�т��K����ȧ�|�������v���N��s��*ن��zd�W�9��2�ܳվ�▾��K��j�����g��û׽�J"���}�q;���   �   W2��Su��꠿Pʿ����L�ȕ �
_/��9��U<�D�8���.� ����JH�%�ɿڐ����t�~/2�i��������M�n��ԛ��,���wr����	�b�M��Ǔ�-ʾ����Q#��B�SQ]�7�r� ���T��;����q�FP\�,�@�*,"�em��Ⱦ������J�$,��ҷ�K����\��S���(L��?��{����   �   Y��+��=��"�*��*�*���A��#U��"b�F�f�0�a���T�z5A��*�Dk���|���	&��U)Y�[��2Ⱦ$%{�}u�
���<�w��Xu� Y��'���|�<���������ܾ	�S����&�W�0��4��p0��\&������@ھ=L��B�8��8��0���1j���m��#��Nq��^y��qǾZ��   �   ��}��Z����߿L�� 	)��XG���d�>~�����ם��}v��X�}��Ed�J�F� �(�<����߿J���q�~�%y2�\�ў��\�.��R�� �T��U�d�.�^L��Q�ֽ�P��X�-���I詾9�ľ�Yھ���p쾚a羡IپA�þT-������[U�4n��kϽ���!���X�H�����a*,�FU���뾳�1��   �   9=��}��=N��rr�^�>��b�����a_������ݡ�����3��Nt����b��>����<���?��������J�-������ F��ѽz�B�ذ���[g��3ɼ��C�����<��N$���M��r��懾.%��*�����������p�@�J�;� ��Y��䜽�N4�t.��H1-������S5��.˽2�B������E���I��   �   *��ѿ4��"�)�dgP��nz��o��wԤ�23��3����"������uk�� �z�^�P��Y*���n�ҿ(����]�HH�a���jY��	��-;�hp ��;�gq;(��8u���k����B뽔���#�n�0���4��/��"�z�%G�(Q����\�D�ݼ��� ��; �<�ɻ~q,�8�ٽ�aU�X���-=��a\��   �   ����uܿ�h���2�>Z\��1����Z����Ľ�Y��A½�^���|����b����\�pc3�4��[Yݿ�Ƥ��i� ��yž��e���&�8����HF�<��<�DO< E#��C����6��󇽉���g�ν��H.�PU཮A˽J㪽:)��0t)�@���G�:<��<���<8��< �q�DO)����C�a��Vþ���DWh��   �   �Ǧ�/�l����5��`�X���������o�����s��⦴��3���C���'a���6�.J�5�r���I�m�w���Eɾgj��z�@c8�����*�<�c�<i�<0!�;`r6�p�����O�ű�������0�����ꀷ��f�����z`D�p+��D���#+<t��<��<�۽<���:�(�@���e��ǾJw�tl��   �   J���tܿJh���2�.Y\��0��#~��S����ý��W��'���T��������a����\��b3����oXݿ+Ƥ�ݪi�`��xž��e�[����8�0��H�<�< FO< B#��C����6��󇽎���q�ν��S.�ZUཱུA˽T㪽>)��6t)�@�� L�:���<���<ԭ�< ^p�M)�����a��Uþ���8Vh��   �   �웿��ѿ����)�reP�lz��m���Ҥ� 1����� ������i��b�z�f�P�X*�x���ҿ͐��݅]��F�s����Y��ὔ);��e �0$�; yq;p���t����k�����B뽗���#�x�0���4��/��"���3G�)Q����\���ݼ�����;H�<�ɻhm,��ٽ)_U�o����;��_\��   �   Y;���z��'K��zp�Ћ>���b�ݗ���\��1���ڡ������0��3r����b�x�>���������������J�4�����L�E���ѽ��B�`����Rg��0ɼ��C�C�����N$���M��r��懾6%��
*����������p�L�J�8� �yY콤䜽N4��+��x(-�����N5�i*˽��B������C�̨I��   �   �}��W��O�߿���>)��TG�2�d���}�Ǚ��Ϛ���s��
�}�DAd���F�:�(����߿U����~~��u2������2�.�qM���T�Q���.��K����ֽ�P��X�(���H詾<�ľ�Yھ���
p쾦a羬IپJ�þZ-������WU�n�ukϽ:���� �����H�8���F&,�#R��Z��c�1��   �   .�X��(��3��+z�&����*���A��U�.b���f���a���T�1A�
*�>h���n����"��f$Y�pW�~-ȾW{� q�1�����w�Tu��W��>���8�<���������ܾ	�T����&�[�0��4��p0��\&������Aھ8@���8�38���.��-j�V�m�.���l��Wy��lǾ���   �   R2�PMu�w栿Bʿ���fI��� �xZ/��9��P<�Z�8��.�� �>��GB��ɿ����n�t��*2�*��������M�m��핬�X���p����	��M��Ǔ�ʾ����Q#��B�TQ]�:�r�"���T��B����q�LP\�/�@�+,"�em��Ⱦ����H�J�t+��з�����0W��i}��dL��:��G����   �   ����C�d�������Ơſ���>��h����l<������t���忭�Ŀ�^��.}���gB��;����0n}�g"���ؽ�?��O+ý�(	�4.N��C��2c׾�4�4�:���e�т��K����ȧ��������� v���N��u��,ن��zd�Y�9��2�ǳվj▾��K�ni�����5b��H�׽VD"�/�}��4���   �   &)Ծ�o�F��`|� ��+����˿�ݿ/]��/���Fݿ ˿���@G��&{�E�;���Ӿ�쏾�z=��c�����遽�c�����>�����`,Ծ�q�#F��d|�[������7�˿��ݿ�`鿻3�
��Jݿ�˿T���3J��+{�JE�����
Ӿ4����=�Xj��(������u���>�>������   �   �@��C_׾2���:���e�]��������ŧ�5���1����r��FK��O��Lֆ��ud��9�?/�5�վ7ޖ���K�Ee�\���_��1�׽�E"���}��6��s��fC�����G�ſ�������i�����>���	��v������Ŀ�a�����JkB�x>�D���t}�Fk"���ؽJA��!*ý�&	��*N��   �   o�M�sē��ʾς�EN#�tB��L]��r�_���Q�����V�q�K\�p�@�("��i��ȾO�����J��&��ɷ�u���EU���}���L� <�������S2��Ou�蠿Qʿz���J��� ��\/�0	9�4S<���8�p�.�. �8���E��ɿ5���~�t��-2�ϱ���4M�m���������m����	��   �   U���7�<�n��?���^ܾ�������&���0�b4�l0�~X&�����ھ�謾���,�8��-��'���"j�֜m����m�Yy�nǾ����X��)�����|�b���*�|�A�� U��b�l�f���a�N�T��3A� *�j��������$���'Y��Y��0Ⱦ�"{��s�뤳�\�w�BPu�FS���   �   ~F��v�ֽ�K���X�,����㩾��ľ�Sھ}��Xi��Z�6CپD�þ�'��䦉�iU��g�4aϽa���� �Ɗ�z�H����g&,��R��d��B�1�p�}��X����߿Ԗ�\)�\VG�$�d�X~�-���S���u���}��Cd���F� �(�b��p�߿U����~�6x2�������.��P����T�O���.��   �   P#ɼ��C�q���G��I$�(�M���r�⇾� ��v%�������b
p�يJ��� �oN콏ۜ�j?4����-�葉��I5�))˽��B�����C�R�I��;��C{��
L��q���>��b������]��x��Oܡ�g����1��ps����b�"�>���Q�����������,�J���/���) F���ѽd�B�T���hDg��   �   `�q;��(d���k�]���:�{���#��0��4�x�/�<"�h��=��H��z�\��ݼ�ʶ����; �<��Ȼ�i,�}�ٽ�^U�=����;��_\��웿*�ѿJ�� �)��eP��lz��n��UӤ�2��$����!��*����j��&�z�ЮP�2Y*�b�+�ҿ���Ň]�AH�j���|Y��	��,;��h �P0�;�   �   ��<�MO<�#��:��ڸ6�<���w���׉ν��	)��O�m<˽Pު��$���k)�d1����:��<ȫ�<���< �l�|I)����٤a�Uþ����Uh����tܿ6h���2�:Y\�1��V~������IĽ��X���������E����b����\�tc3�F���YݿǤ�U�i�|���yžԬe�2��p�8� ��4G�<�   �   ���<܈�<0,�;H��d�뼎^C�O���_���O\��OW���*�������3|���4�p�ʼ�'���G<L��<���<�K�< �v;D ���ٽX�Y��N�����{�a��U��"Gֿ�_
�4�-��)U�)p��딖����ӗ�����q���Lީ�[ݖ�i��N?V�&�.��a�c�׿ڿ����c� �������_�4佔�,�����s�<�   �   �/�<ȸY<�����m���Y+��z���q��Ľ�ֽ�&ܽ�MԽ�Ŀ��l��p5r�n���L�� CX;<F�<���<t"�<��: ��rֽ��U������4���]������ҿJ-���*�NQ�ҹ{��R��#���v��6Զ��q��S���냓��o|��:R�Ο+�&	��pԿU��h�_��	�]㼾�q[�&\ཆY-�@!6����<�   �   �d�;��<�"8^�����ְ߽�&��>(�,��'�|��\x��ؽ�Y��8�K�X�ü`T���<X�*<`Ew�*��/v̽�8J�j���;C�.?R�y�����ȿj���a"��VF� 1m����������	���x����������rm�>�F��
#��z�	ʿ���F"T�t���Y���XO��ֽ��/��[�0h�;�   �   `�����7�+���A轕���qD���g�����삊�cJ��}Љ��p��4&d�j#@�f
��m޽�=��fq$��&��-���f�L�%�������8���������h@��݈��!�����P����5���W�4!y���8��W�� ���ݼ����x��mW�`�5����{f��A���Z�A�J9�]�� �<�h\ǽ�6��[��0�L��   �   ,ڀ�Hv̽���OO��j��-t��TS��+�о��ݾ׶ᾠ�ܾaϾ�3�������Ƃ���I������½zao�.F�������8�U���#�����X�)�̰r���{,ֿȽ��!��7>�4�Y��p��@����������o�j�X�d�=�P`!����jTֿ�H���s�,�*���񍾇�&�;x���.H���c#��   �   @��4���|�`����ҾB���~���J)�c,��z(�d����L���ȎϾ�m���w�/��齕�����X�Ҍ\��Y��˃�m�����&�%YO��Ǎ�f�����(��VN#��9�4K�PW�:[��{V�d/J� 8�rr"�: ����߸������n�O����n+��:�o�5<�N>��Fpi�>=g�׊���   �   wJD��@���T������X���9���S�,Rh�`.u��Zy��}t�6g�iJR�
8����gk��+h������x@�Sc�������1��,��(��BB�曚��g뾳e*�>�j��&��]���-0���������'���0��3�ZV0�<�&��������迯���ٍ��Nj��)*�Ww뾈��^XC��^�X���@������B��   �   Jv��&�;��
�G�2�= \��ၿFK���֠��Y��N���䨿���?��zĀ��Z�>�0��e	��x˾�����A�v$ ��u��EF����˽d,���q�<i���`�.�:���v�vB��٢��mݿ�_�����������-����N�����ۿ�D��5�� yu��9�b���ɷ��cq��b�dqͽ빥�~��u���D��   �   ��ʾD���=�|�q������3����ÿ��Կ��߿�T�?2߿g�ӿ#5¿׫�Rr��U�o��<����,ɾ4���4��+�砲�'�����Z�5��"���ʾ���=���q������0���ÿ��Կ��߿!Q㿥.߿�ӿ2¿_ԫ�p����o�	 <����
ɾ  ��J4��)�w���<*�����&�5�n&���   �   Ec�̑:�i�v�+E�������pݿ�c�����ҕ� ���/����������ۿG�� 7��'|u�Q�9���
̷��fq��c�nqͽ�����踽�q��D�@r����;��
��2�S\��ށ�9H��VӠ��V����`ᨿ����T<�����Y���0�Bc	�u˾���i�A�|" �jt���G����˽�/��q�Bm���   �   �h*�#�j�K)��;���3�ԅ����8�'�2�0�p�3��X0�@ '�������迱���m����j��+*��y�����YC�N_��V���<�������=��CD�a<��:O��M����T�D�9���S��Lh��(u�Uy�zxt�=
g��ER�.8�l��f���c������	@��]������f1��!�����LB�����l��   �   @\O��ɍ�������ڼ�PP#��9��K��W��[�~V��1J��8��s"�j!����X��������O�����,����o�~<�=��ji�3g�{���&��q�3�6~|��Z��G�Ҿ����������(�,��v(�u��e�������Ͼ�i��Xw�=
/�T��Z�����X�D�\�N\��l��jm����)��   �   ճr��錄�.ֿ,����!��9>���Y���p�B��6�� ��F�o�<�X�ΐ=�da!�j���UֿwI��2�s��*��⾆񍾸�&�(w���)H�<�@X#��Ҁ�Zl̽:�?HO�5f���n���M���о$�ݾd��e�ܾ�Ͼ�.�����Â���I����a�½�Wo�N@�����J�8�A���#�=��d�ྥ�)��   �   �ވ�Y#����ￔ���5���W�x#y�^�����QX��/���ཊ�2�x��nW�>�5����`g�񹿱�����A��9������<�K[ǽ��6��O���nL������7�L���6�F��RjD���g�����~~���E��:̉��l��d�+@�#�e޽7���g$������(�f�β%�������8���������j@��   �   �����ȿH���b"��WF��2m���������
���\���G�������sm���F�#��z�Lʿ���b"T�s���Y��nXO�?ֽ��/��H����; ��;�� �Z*^���� �߽ګ���<9(���+�C'�����s�ؽS��ލK�l�ü`�S���<�+< Nw�4��6y̽3;J�L����D�AR��   �   ����*�ҿ�-�X�*�OQ��{�VS�����cw���Զ�r��������� p|��:R�ʟ+�	��pԿ"���_�,	��⼾�p[�WZ�V-���5����<9�<h�Y< ܩ�$_��4Q+�Wv���l���
Ľ��ֽ�!ܽ�HԽr����h���.r�����C��`vX;TJ�<h��<�!�<���:h��,ֽ��U�;ù��5��]��   �   oV���GֿX`
���-�l*U�hp��&���O���헶����Y���ީ�!ݖ�,���>V���.�da���׿L�����c�G������+�_���$�,��h��hw�<P��<L��<�8�;x�����T]C���������\��=W���*��憚�44|�x�4���ʼ`1��@G<8��<(��<dG�< Wv;���ٽ��Y��O��q��j�a��   �   𰜿K�ҿ^-���*�
NQ���{��R�����Yv���Ӷ�q������H����n|��9R��+��	��oԿr����_�r��Ἶ]o[��X��S-���5�d��<(:�<��Y<�ԩ��^��Q+�Uv���l���
Ľ��ֽ�!ܽ�HԽ~����h���.r�Ș��C�� xX;�J�<d��<|#�<@
�:h���ֽw�U�E¹��4��]��   �   \���s�ȿ:���a"�VF�`0m�E��K��������i���~���'��@qm���F��	#��y��ʿr��p T����W���UO�ֽ��/� >����;P��;P��L�*^������߽ܫ���C9(���+�P'�����s�ؽ�S��K��ü�S� �<�
+<�'w�P��$v̽�8J�x���9C�?R��   �   ݈�!����￺����5�~�W��y���
���U����������P�x��kW���5����`d�Uﹿݤ��3�A��7�����<��VǽL�6�HH��8eL�D�����7����6�8��MjD���g������~���E��B̉��l��d�3@�&�e޽�6���f$�@��P���f�n�%�t���`�8�����>���h@��   �   ��r��I+ֿ���
�!��6>�h�Y���p�h?��n�����f�o��X�d�=��^!�2��Rֿ�F��Ԑs�֨*����z��&��q��6#H����U#��р��k̽�&HO�.f���n���M����о,�ݾo��o�ܾ�Ͼ�.��'���Â���I�����½,Vo��=�x�����8�7���#�>�����z�)��   �   �WO��ƍ����َ�����L#��9�
K��W��	[��xV��,J��8�zp"�����q�������L�O�#���'���o�)8�a7���bi�X.g�����8��(�3�~|��Z��>�Ҿ����������(�
,��v(�{��i��#�����Ͼ�i��Dw�
/�������d�X�F�\��V��+���m�/
���%��   �   �c*�۱j�S%��a����-�v�������'���0���3� T0���&�������O������q���hj��&*��r���;SC��V�6Q��9��>���#=��CD�<<��%O��<����T�A�9���S��Lh��(u�Uy��xt�D
g��ER�28�o��f���c��v����@�g\��s����-�����S����A�2���$e��   �   �^�ˋ:���v�z@��n���)jݿ�\�����������+����}���k�ۿ�A��Q2��tu�L�9�����ŷ��]q��]�!iͽ����丽�p�9�D�
r����;��
��2�N\��ށ�9H��WӠ��V����cᨿ����W<�� ���Y���0�@c	�u˾���НA�t! �q��BB����˽�)��q��f���   �   ��ʾ����=���q�l����-����ÿ��Կ8�߿eM��*߿e�ӿ�.¿7ѫ�<m��ƿo��;�W��ɾ_����4�� �a���#"�����X�5��"����ʾ���=���q������0���ÿ��Կ��߿$Q㿩.߿�ӿ2¿dԫ�p����o�	 <�����ɾ����^
4��&����"�����5�� ���   �   eo����;��
���2�Q\�z܁��E��`Р�iS�����ި�����R9��^�����Y���0��_	��o˾�{����A�u �l���?��}�˽+���q��h��n`�#�:���v�sB��ע��mݿ�_�����������-����S�����ۿ�D��5��yu��9�V���ɷ�$cq�Ua�Cmͽ~����㸽�n�͞D��   �   8?D�(9���J�����}Q�P�9�`�S��Gh��#u��Oy�st��g��@R��8�u��N_��^��2���H@�S������)��������!B�����dg뾤e*�6�j��&��[���+0���������'���0��3�^V0�<�&��������迳���ٍ��Nj��)*�1w�<��QWC�n[�NS���8��t���h:��   �   ���^�3��w|��V���Ҿ���� �ί���(���+�Ur(�J��������r�Ͼed����v�v/���齷���D�X��\�kU��_��1m�q���&�YO��Ǎ�c�����&��TN#��9�4K�RW�<[��{V�f/J�8�rr"�< ����ุ�����k�O�w��6+��k�o��:�:��jci��*g��}���   �   �̀��d̽F��AO�^b��bj��LH��)�о��ݾ��	�ܾnϾ)���🾓�����I����+�½Go��2�������8����#������N�)�ǰr���z,ֿȽ��!��7>�4�Y��p��@����������o�n�X�f�=�R`!����mTֿ�H���s�&�*��⾷�����&��t��%H����O#��   �   �����7�t��N.���dD���g�����Hz���A���ǉ�Wh��3d�@����uZ޽&.���X$�`����0kf�F�%�8���;�8�ȼ�������h@��݈��!�����P����5���W�4!y���7��W�� ���޼����x��mW�`�5� ��}f��B���W�A�>9�*��J�<�Zǽ��6�tG���WL��   �    Ƙ;������^��
��n�߽���	�4(�R�+���&�j��o�1�׽�K��F�K�,�ü�S��<�"+<��v�����t̽A8J�F���1C�+?R�x�����ȿj���a"��VF� 1m����������	���x����������rm�@�F��
#��z�
ʿ���E"T�m���Y���XO�&ֽ�/�pA����;�   �   �;�<��Y< s��PV���K+��r���h��uĽ΃ֽ�ܽ�CԽo���!d���%r�Đ��5�� �X;XU�<X��<L+�<�|�:د��ֽf�U������4���]������ҿJ-���*�NQ�ҹ{��R��"���v��7Զ��q��S���샓��o|��:R�̟+�&	��pԿV��h�_��	�O㼾vq[�j[�HW-� �5����<�   �   8��<��<`14<��������&���e�d���皽:���0���u���;W�T���� ]�9丈<ܣ�<Hg	=�y�<�B<l��O����D� ����I
��bO����|ƿX���> �&AC�@;i����/a�������ŧ��ƣ����]��Ej���D��[!��;��@ȿ����
IR����=�����K�9X̽�F��D;$%�<�   �   ���<��<�b1;�>z�����m_���	W��0I���*Ľ󀼽u������ M�  ��Pw ��
<�<���<��<�T�;�S�'���A��R������K�ق���¿#����s�r�?���d���j��U������/�����_!����e�Z�@�V��,9���Ŀ�-��K�N�3
�<��9�G���Ƚ����@�:��<�   �   0�<�<d��`��7?����OdȽB��6�i)��{����
'
�cG�G���fÉ�v(�TҊ��S;h�f< �w<���:�����U���N6��韾�t ��=A��^�������B�.�I6�|TX�Xz�����ﰕ��/��ƍ������z�y��X�T�6�
�����HB��]�����C�@{�5s����<��P�����@�z�`<�   �   L��<b�m����MнM��\�2��9S��l���|��ހ�O{���i��N�J@-���XĽp�z�Z�X�:�@��� �(���ɦ��	&�j��2�|�0��J|�6����ݿ��
���'�>�E���b���{��\��8G�����N{�t&b�*aE�<�'���
���޿���A~���2��t�rc���+�s���>W��W� v���   �   ~`�m�����<�R�s���&���_��	,˾T�ξ.!ʾ�k��i��������Gm��#6�v*�jH���SI����ຼ�S������X��~��;����_�[��3Hƿ����ʚ��F/�iG�ʥ[�,i��m��h��Z��\F�(|.��*�A����yƿ;̘���`��-�Ͼ ���U�������M*����:)��   �   �ٽ#d#��f��\��{V���8��b�&���v�7+����������ۊ侅���j���6�_��:���νb����u5�49�����`R���W�����A���>��ۂ��2����ֿ������*���:��2E���H��D���9�|�)����� ���տ�Ѫ��т��*?�������S;Z��
�G��VI�8$G��{���   �   j]2�8 ���V��e���E@+��lC�MV�n)b�M�e��La��T��_A�J�(���HB�����|�l-�A2�쯖���o�,u��ѧԽ�v/���C�׾���`X�0y���}���(ٿ�1�����9��J#���%��"�j5�<h����Em׿�G��������W��_�	�׾k���n 1��ؽ�����|�t ��_
��   �   �j＾%���+�$��K���o�d,��������!����Y����܆��(m�^qH�o"�����%׹�����e�.�Ő�Ta������ϡ����
���[�������Y�+���c�����z���<UͿ�N����4�P�6������%E�*V˿���L2��gb�y�*�MM������Js[���Ew��Q���֫��:L��2��   �   lչ����.�.��:_������\��R/���QſjgϿ��ҿa�ο��ÿ����U��������\�x�,�*��÷�7My���"�tUԽ�G���흽�Xֽ�U$�X|��й���n�.�N6_�����Y��,��xNſ�cϿA�ҿ�ο��ÿ����٥��� ���\�¯,� �����^Iy�h�"��SԽhH����\^ֽZ$��|��   �   ������+���c�?���i����XͿR翷���&�@!���K���3H��X˿X���'4��Vb���*�wP������u[���Hw�����;����D꽇�2�0섾u꼾҄��H�$��K�|�o��)������������&������چ�k$m��mH�l"�ͨ���ӹ����!�.���'`��ű��~���>�
���[������   �   ���NdX�n{�������+ٿ\5�����;�M#���%��"�<7��i�w���o׿_I��0����W�Ta�2�׾�����!1�d�ؽV���~|�v����hW2�>���Q���^�b��<+��gC�HV�E$b�,�e��Ga�s�T�S[A���(���N=�)����{�^-�-�,�����o��v��+�Խtz/��
��Z�׾�   �   ��>��݂��4��o�ֿ�������*���:�<5E�ܟH�.�D���9��)����� �W�տӪ��҂�,?�������<Z��
��E���I��G��t����ٽ�]#��f��W���P��O2�_�;���r�,'����ܱ�h��"�侸�������,�_�6���νq���:r5��9�����;W��� W�����C��   �   �_��\��\JƿT���N���H/�"kG��[�p.i�l�m�<�h��Z�v^F�l}.��+�Ǒ���zƿ͘�¨`���(�Ͼ����~��|���I*��⼪�>`��c�����<���s�����Ĝ��@Y��&˾^�ξmʾ]f������^����@m�86��%��A���JI����ܺ�DU������[��~��;����   �   GM|������ݿȁ
��'��E���b��{��]��XH�����{��'b�8bE��'�f�
���޿���kB~��2�u�c���+�e���^S�@�W� 7��x����T�(y���Cнr����2�2S�)�l���|�pڀ�l{�W~i�H�N��:-�<��tĽ(zz��P���:����h� �|���̦�&�l���4�t�0��   �   `�����}D�"�@J6��UX��z�����۱���0������=���t�y���X���6�X��a��B��}�����C�?{�s��&�<�sO��>���Sz�<��<�c��J��.*?������[Ƚ�8��G��U$��v�Ǣ��"
�:?�3���p����(�xÊ� �; �f<�w<���:\����X��/Q6�h럾�u ��?A��   �   �����¿N����t�D�?���d����������`����������!��&�e�j�@�R��9����ĿX-���N��
�;��F�G�5�Ƚj��@��:D#�<@��<��<��1;P#z� ��e_�Z.R��CD��&&ĽZ|��@���{���M�p���g ��
<Ĭ�<8��<8�<�H�;Z�G*���	A�
T�����d�K��   �   ����ƿ���� ��AC��;i�����Za�������ŧ��ƣ�����,���Dj�4�D�<[!�/;�@ȿ���/HR���:���H�K�V̽vC�@4D;D)�<ܟ�<0�<P74<�����&���e�����暽:���0��(v��n<W�8���� Ƚ9<��< ��<�e	=v�<89<���Q��(�D�"���NJ
��cO��   �   ���7�¿I����s�l�?���d����'�����k��������� ����e���@�����7���Ŀ�,����N�4
��:���G���Ƚh���ذ:�$�<P��<l�<��1;�"z�޿��d_�X3R��ID��/&Ľc|��E���{���M�t����f ��
<P��<$��<��<PR�;TV��(���A�'S����w�K��   �   �^�������B����H6��SX�lz����)���/��ٌ��������y���X�&�6���[���@��C����C��y�Xq��ޮ<�~L��X�� +z�X < �<��c� J���)?������[Ƚ�8��K��Z$��v�Т��"
�I?�?���r����(����;X�f<��w<��:,����U���N6��韾�t ��=A��   �   �I|����4�ݿ�
��'�<�E�t�b� �{��[��F�����{�|$b�|_E�ط'���
���޿d��?~���2��q�Ha��ۖ+�@���N�(�W��$������T��x���Cн\����2�2S�)�l���|�tڀ�x{�b~i�T�N��:-�<��lĽ�yz�RP��:� j��t �t���Ȧ�	&��i��m1� �0��   �   �_�9Z��GƿM���ؙ��E/��gG��[��)i���m���h�țZ��ZF�`z.�P)�����wwƿoʘ���`�����ϾĦ����������B*�������`�8c����ȸ<���s�����Ĝ��CY��&˾e�ξvʾgf������d����@m�:6��%�nA��8II�P��hԺ�DO�����W�|�~�Ғ;����   �   H�>��ڂ�,1���ֿ
������*���:��0E�B�H���D���9�z�)���
� ��տvϪ��ς��'?�z���
��w6Z����@���I�4G�s����ٽ�]#��f��W���P��I2�_�=���r�0'������l��*�侼��������_��5���ν9���n5�9���XO���W������@��   �   G��z^X��w��|���&ٿ%/�����8��H#���%���"�^3�Vf�H��5j׿�D��y���
�W��\���׾>����1�;�ؽ����f|�)��3 ��V2����Q���^�[���;+��gC�HV�J$b�0�e��Ga�z�T�X[A���(����Q=�"�����{�-��+�����o��q��2�Խtt/�l����׾�   �   G���!�+���c�݁��8����RͿsK�~���Z�d�F��!����A��R˿1����/��6b��*�H��
�\m[���o��򲑽գ���B�؈2��넾R꼾����@�$��K�x�o��)������������)������چ�r$m��mH�l"�ʨ���ӹ�怂���.�)���\��ج��㝴���
���[������   �   �͹��}���.��2_�����W��7)��UKſ�`Ͽʏҿ��οx�ÿ|��袞�������\��,�(�V���eBy��"�KԽ�@���蝽�Uֽ�T$��|��й���f�.�F6_�����Y��,��xNſ�cϿE�ҿ	�ο��ÿ����ޥ��� ���\�ï,�������Hy���"��PԽ�C���靽	Tֽ�R$�|��   �   �鄾�漾
���?�$�:K��o�
'��=����������
������<׆�Qm�(iH�@h"������ι�.}��,�.����FX��u���������
���[�����]���L�+���c�����x���:UͿ�N����4�R�8������)E�.V˿���O2��ib�v�*�7M�������r[�L
�_s��L���ۢ��.?꽯�2��   �   �R2�?���M���Y�I��W8+��cC�oCV�Xb��e��Ba���T��VA�r�(�G��7������{�-�#����fo�
p��i�Խ�u/�����׾թ��`X�,y���}���(ٿ�1�����9��J#���%��"�n5�>h����Hm׿�G��������W��_���׾!���o1���ؽ겏��
|����+���   �   ��ٽ<Y#��f��S���K���,��[�����n�*#���� ��ϼ��~����¨��X�_��/���νZ����d5�9�p񎽪O���W�Ȧ���A���>��ۂ��2����ֿ������*���:��2E���H��D�§9�~�)����� ���տ�Ѫ��т��*?��������:Z�<	�C��HI��G��o���   �   ��_��\��|���<���s�{�����S��] ˾z�ξ�ʾ�`��J�������D8m�16�, �F8�� ;I�L�弜ź��J��~���W�M�~���;����_�[��0Hƿ����ʚ��F/�iG�ʥ[�,i��m��h��Z��\F�(|.��*�C����yƿ<̘���`���Ͼب��^��j���tD*�@�����   �   �(K��r���;н�����2��+S�ڷl�Ǿ|�hր�b{��vi��N��3-�y���	Ľ�iz�2C��:�@���] ����qǦ��&��i���1�u�0��J|�3����ݿ��
���'�<�E���b���{��\��8G�����N{�v&b�,aE�>�'���
���޿���A~���2��t�Bc��k�+�?����P���W�����   �   ��<�Pc��;��^ ?������TȽ�0��������q�ҝ��
�76�����&���.(�ĭ��`=;X�f<��w< ��: ���IT��uN6��韾�t ��=A��^�������B�,�I6�|TX�Xz�����ﰕ��/��ƍ������|�y��X�T�6�
�����JB��^�����C�:{�s��8�<�YO��Z���7z��%<�   �   ���<���<��1;(z�غ��^_��뒽N���?��{!Ľ�w������Sw��<M�����XL �8+
< ��<���<(�<0m�;�O�'���A��R������K�؂���¿"����s�r�?���d���j��U������/�����`!����e�\�@�T��-9���Ŀ�-��J�N�0
�<���G�7�Ƚ������: $�<�   �   ���<���<x)�< ��:��m������o5���a��i|�K�����u���T��/#� ˼����}<���<�;=��=��=���<8����l���z(�N���o��7�����k���&,�:��W-��L�0l�0|������7	��i�����0�l���M���.�4O�����5�����:�2���E���1�ʗ��X�Ӽ8�<���<�   �   �|�<�ѫ<pU<p���$�мT�/�,o�����V碽����v���\����P䛼 A� ��<�F�<޷=���<�%v<��������)%�8�����]4������#�����J��\�*�fXI��g��̀�����4��ع�� ؀�,�g��J���+������A2��T��c7�����8���z-�z��|KԼ &�;(��<�   �   �N`<@nF;`�k��f��r�~ا���н¾�R3����.c �����%ǽ�᛽��W�(&켠��P-<��<H��<�:%<{��ᐽ��T��]����*��Et��̥�^׿v=��W"��?���Z��~r��S���&���3��5r�.�Z��V?���"�>��ؿ�n���8w���-����+q��kT#�u�����׼ �5;03q<�   �   ����%��_��3�����K�9i7��!N��F\�gt`��AZ�-LJ��2�^�������-@��⨼@P��Б�;@7�:���ۅ��9���|���;^D��`�����#�ƿ_��J�� �/�
�G��2\���i���n�$ti�D�[�
,G�`4/�������˂ǿ����8b��@��tѾ8����1��xA�`��� X=��   �   L�0��ܗ�t齜�#��T�Y��$���E��{���`⵾@���&
��g���!�}�1�L�����ٽ���~
��c�� zL�\�ϼP�t�a���q�\�7S��(�	��RF�ￇ�L���޿���f�� 1�$�A�M���P��mL���@��0�x��N��I�ݿ��s7����G���
�4����@b��>�⥅�y�����؇¼�   �   ���~��r�H�0���v5����̾������	�(��m��r� �t�e�Ⱦ?ե�5��$�@��6�/
�J��`�t��tb���ҽ��9����!�9)�E�h�ؘ� ���&� R�����I&�6!/���1�z~.�:%�T[��I���D;��s��ߵh��d)�.h�Č���[=�۽ґt�^.����r�c��   �   L����a�@䛾N2̾����3���k-��Q>���H��9L���G�ʛ<�-+��F�ݟ��zǾ����-Z���3���8Op�B"9�NH[�˛���k���u����}
��@���}��h���~¿*��=���b�
�� ��9��k���	�p4�����Զ���$���E|��8?�l+
�mɽ��w�f�:޵�<Hh���H��^��ǽ�   �   =+h�d)��p�ᾟ���W4��wU���r��������n���0��������o��qR��n1�u_�WXݾ@���<{b�jw�\������V�c�pG����C�>��֓���پ#��J��Ҁ�� ���շ��IϿ�v�����Z�v��B�߿5Ϳ�ĵ�5����~��H����5�׾�󒾬�=��)�����RQk�����_�Ž����   �   �C��}����fF��Us��*������t���8����y���ܸ�R*���?���\��bp�@�C���?6�T䠾7QX���
�M���"�~��F���2��Z����[��?���w�����bF�Qs��'������U������pv���ٸ�}'���<���Z���p�&�C�z���2㾼ᠾ�MX�}�
������~��I��8��T��W�[��   �   ��پ$���J��Ԁ�]���ط��LϿz�q��A^����T�߿�7Ϳcǵ��7����~���H����	�׾������=��+�����PMk��􅽶�Ž����$h��$��ǰ�&���S4�%sU�~�r�]��������퍿������i�o��mR�bk1��\�Tݾ����vb�~t����k���j�c��J����ܗ>��ٓ��   �   �
��@���}�Ak��u�¿L�⿬���4�
����;�Nm���	�I7�������`&���H|��:?��,
�]˽�2w�Cg��޵�BEh�X�H�4Y���ǽ���ׄa��ߛ��,̾���b��g-�7M>��H�R5L�r�G���<�_)+��C�^����uǾ�����(Z�B������>Jp�f!9��K[������n���u������   �   �	)���h�ژ��"��y)迶S����xK&�,#/���1�L�.��;%��\��J����<��Vt����h�,f)��i�܍���\=�u۽��t�)����c��������f�H��~��S0����̾V��n��7|	�������0� ���H�Ⱦ�Х��1����@�|2��詽��J�<]���yb�G�ҽF�9����%��   �   _UF�����N���޿r��~h��1��A��	M�z�P�joL�8�@��0����.����ݿ+���<8���G�m�
�����Ab��>������p��L���t¼f�0�|ԗ��i�8}#�r�T��T��S����?��(���ݵ���\������x}���L�q���ٽ���D��Y��sL��ϼ$�t�����\��U���	��   �   �`�-����ƿn��~����/���G��4\���i�l�n��ui���[�0-G�F5/����������ǿ)����8b�A�RuѾh����0��t:㼀u�� �;�]�����^��*��J��E��b7�oN�l?\�m`��:Z��EJ��2�/���w�����!@�8Ҩ� �����;�I�:�����ޅ��;�E�|��;!F��   �   |Gt��ͥ��׿N>��X"�?���Z�8�r�xT��R'���4��&6r���Z�fW?�`�"���w�ؿ,o�� 9w��-����q���S#�G�����׼��5;�Gq<�h`<`�F;(�k� [���r��Ч�n�н���.�$���^ ���齎ǽLۛ��W���0h㻨�-<���<�<�8%<0����㐽���U�����Y�*��   �   �����$��������
�*�0YI���g�R΀�#������)���Z؀�v�g��J���+�������2���S���b7�S��R8���y-��x���EԼ@?�;��<���<�ګ<�j<�`���м��/��#o�Y���Sꞽ�⢽퀛�5s��:�\����ڛ� V�x��<J�<��=��< v<D������+%�|���`���^4��   �   ��������,忎��W-�j�L��l�Q|������7	��W�y���ޕl�T�M�:�.��N�_��l5��v�����:�����.D���1�ʕ��d�Ӽ��<܊�<���<���<X,�<@�:0�m�d����n5���a�Ri|�:���&�u��T�D0#��˼0���y<d��<::=|�=��=h��<����n��&|(�7���@p��7��   �   '����#�����P��T�*�HXI��g��̀�c������g����׀�J�g��J� �+������X1��LS���a7����7���x-�w���AԼPI�;��<��<�۫<l< _����мx�/��#o�\���Sꞽ�⢽����4s��>�\����ڛ� S����<�J�<�=`��<p$v<��������*%�����8��^4��   �   WEt��̥�׿:=�.W"�d?���Z��}r�S���%��63���3r�֭Z��U?���"�b���ؿ�m���6w�l�-�H��zo���Q#�����h�׼@6; Nq<(m`<��F;@�k��Z�D�r��Ч�a�н���.�&���^ ���齙ǽXۛ��W���@f�H�-<(��<t��<�@%<�y��	ᐽ"��'T��\����*��   �   �`�;���p�ƿm�����H�/���G��1\�X�i�Θn�Hri�z�[�l*G��2/���������ǿ'����5b��>�'rѾB쁾���5-���0�[�� ;�0W���(�^�M*����
E��b7�lN�p?\�!m`��:Z��EJ��2�6���w�����!@��Ш��{��@��;���:�물�څ�9��|��;�C��   �   �QF�0���K��@ ޿F���e�~�0���A�2M���P��kL���@���/��������ݿ%}���5��g�G���
�R����<b�j;�q����d��d��to¼��0��ӗ�/i�}#�X�T��T��P����?��+���ݵ�"��c������x}���L�n����ٽ̱����U��eL� �ϼ��t�d����\�>R��n�	��   �   �)�q�h��֘�����$��P�����G&�d/���1��|.�08%��Y�&H�R���8��q����h�2b)�6d�҉��eW=�۽̅t��"����:�c��������-�H��~��B0����̾O��m��9|	�������5� ���M�Ⱦ�Х��1����@�P2��穽��J�hY����ob� �ҽ�9��& ��   �   �{
��@���}�*g���|¿���g�����
�&���7��i��	�1��������G"���A|�T5?��(
��Ž�
w��a�׵�T;h���H�W��|�ǽn����a��ߛ��,̾���]��~g-�7M>��H�V5L�v�G���<�c)+��C�c����uǾ����j(Z���^���vFp�N9�"B[�|����i���u�����   �   �پ%�u�J�р������ӷ��FϿ�sῤ��\W����߿�1Ϳµ��2���~�A�H�����׾�P�=�@!��}���Ck��񅽞�Ž7�� $h��$��������S4�sU�{�r�]��������퍿������o�o��mR�gk1��\�Tݾ���~vb��s�C�������b�c��C�����S�>��ԓ��   �   �<��t�O���_F�:Ms��%��k����������Ms���ָ�k$��:���W����o��C�#��I-㾡ݠ��GX���
�Ʊ���~��B��0��i����[�c?���w澸���bF�Qs��'������V������sv���ٸ��'��=���Z���p�*�C�{���2㾞ᠾSMX���
������~�KC���.�������[��   �   �h��!�����k��AP4�,oU���r�ޟ������ꍿ���i���^�o�]iR�Yg1�SY��Nݾ�����ob�o�����9�����c��C�����s�>�c֓�˘پ��J��Ҁ�� ���շ��IϿ�v�����Z�z��H�߿ 5Ϳ�ĵ��5����~�
�H�����׾p� �=�d'�a���JFk�������Ži���   �   ���sa�(ܛ�/(̾v������c-�I>���H��0L���G�4�<�8%+��?�ѓ��pǾ���S!Z���������;p�b9��>[������j�0�u�ٱ���|
��@�x�}��h���~¿)��>���b�
�� ��9��k���	�t4�����ֶ���$���E|��8?�e+
�Lɽ�Lw�,e�>۵��>h�L�H��T��~ǽ�   �   $~�������H�T{���+����̾o��,���x	����[���� �&	�}�Ⱦ�˥�M-����@��,�uߩ�2�J��P�Z�.mb�`�ҽ�9����!�,)�=�h�ؘ� ���&� R�����I&�8!/���1�|~.�:%�V[��I�!��F;��s���h��d)�h꾑���[=��۽b�t�P#�ҋ��yc��   �   ��0�Η�?a��w#��T��P�� ���";��
����׵��y��L ��_���p}�n�L� |�d�ٽ����6���B��JL�`�ϼl�t�t�����\�S���	��RF�쿇�L���޿���f�� 1�$�A�M���P��mL���@��0�z��P��M�ݿ!��t7����G���
����G@b��=����h��p��8f¼�   �   B����8�^�G#��u���?��\7��N�p8\��e`��3Z��>J�p
2�L��xm� ���@�0����R�����; O�:p䬼�م��8�`�|�l�;VD��`�����"�ƿ^��H�� �/��G��2\���i���n�&ti�F�[�
,G�b4/�������΂ǿ����8b��@��tѾ
%���/��45��X�� Q:��   �   �x`< EG;��k�<R���r��ʧ�*�нܭ�z*����dZ ����tǽ�ӛ��W����P� �-<��<Ġ�<PQ%<,s���ߐ�����S��I����*��Et��̥�]׿v=��W"��?���Z��~r��S���&���3��5r�.�Z��V?���"�>��ؿ�n���8w���-����q��T#�*�����׼�6;�Rq<�   �   8��<�ޫ<v<pC��Ȭм��/�o�����S枽�ޢ��|���n��6�\����P͛� ��0��<xS�<�=��<�0v<�������)%�*�����]4������#�����H��Z�*�fXI��g��̀�����4��ٹ�� ؀�,�g��J���+������B2��T��c7�����8��iz-�uy���GԼ�<�;��<�   �   d�=(��<��<��<@q��H�������\"���8�Dw=��&0����H�ɼ�6� �z;�<2�=�}+=�;=F}*=<��<�@��D2b�����z��y;YK� `�u���Idƿ�������[/�x�G��\���j���o���j���\��;H��0�j��D���ȿ(���6�c����-FӾ����w�L��x�u��?{<��<�   �   ���<d��<`w<@1�:P�l�T��v?/�n�X���q��kw��+i�~.H��A�I�� ��/<p��<�$=,=P�=���<@꛻
�]����ݖu��ɾ���K\����p?ÿ���7��w,��ID�zhX�
	f��j�4�e��vX���D� -��������Eſ����_����K5Ͼ���:���8��pv���f<��<�   �   ��<��&<�ˤ�4�¼h4� ��Vi��á��;)ѽXս2�̽V���+��d�e��T�xh�@��;8ĩ<���<�<�<�y�<`���"gP�X���Kg��~��yf��"Q�Ɏ����M��_�P)$�R:�d�L��6Y���]�Y���L�(B:��a$������̖���N���T�h�wpþ��p����v�@.z�pc%<�ܧ<�   �    ������z�#�G(���ý�b��Y9���*�ܠ6�1�9��E4�� &����ߎ�͑��6k��9���.߻�Y<d�<0aH<�H����=�+�ཉAQ�5+��<����?��H��j����ֿb��Pb�d7+��v;�T/F���I�z�E��:�n�*�P"���\�׿�o��fG����A�����0��4HY���N=`��ⅼ�=;�S�;�   �   <H����i�&ʻ��o���0��8Z���~�У���������3��%����w� �Q���'�W��k���0�A�X���𣂻  k��!;�,�*��½��5�U���I��C)��i��혿~*��M,�ZZ�0���{&��q/��c2���.���%�b��r��Pl��^����i�&u*���D��'<�Mн��G��������S��   �   7揽}�!�&���a������k����Ǿ��ܾ��龖���'�پ��þKΨ����U|W����)Zҽ��|���莼������dy��ܒ���}��ž{��jRG���������;ɿ���j����^��r���B�������=�ǿ�'��#���=G��J� rƾ��\��嚭�v+3��>˼�}ɼ��%��   �   ������;��-���׬�YؾeE����`�"���+�ۆ.��*��� �`��N��K�Ҿ�����|��3����惏���'�P�����b>��c��8L�����q$���#�R�Y�	*����� �Ŀ�xݿ���\����f �����M￙mۿ�¿Fq��2����9X��!#�y��՟��oM��K���Ō�,�'��~���?�-4���   �   ,DA��닾R��1}�������6��P�q�c��p�h�s�y�n�ïa�QM���3�� ���T���O䇾%�:���ｋ��x�8����L\��o����� �w�d��@m�&-��]��3��κ���M���:ÿ�'Ϳ�?п�J̿Y����k��{Ҝ�!����fZ�� +� �96��~~u�����+����a�#)�X2F�TК������   �   �B��^Nþ����)��P��6v�"����W���L���Ƣ�ݖ�����������r��pM�+�&����Ŀ�_���B-2��L޽3↽B�8�x�:�3���ך��6�?���Iþ#���)��P��1v������T��!J��Ģ�2��� ���ؽr��mM�y�&��������"���C*2�JI޽�����8��:��������6��   �   T���o�b)-��#]�(6��i����P���=ÿ�*Ϳ�Bп�M̿���n���Ԝ�샅��iZ�(#+�� ��8��āu�����-����a��)�+F��ʚ�1���g>A��狾3M��0w��j��|�6�jP���c�	p���s���n�g�a�MM�1�3���D󾮊���ᇾL�:���ｦ	����8���PR\��t�������w��   �   �(뾴�#���Y�',�� ����Ŀ�{ݿ�� ��kh ����"�pۿ0�¿s������ <X�R##��{�zן��qM��M��ƌ��'�
y�N�?�X-��9�����;��)���Ҭ�KSؾB����x�"�}�+�ڂ.�9�*�=� �"��hH����ҾA�����|�3�������,�'�ȵ����A��2��L������   �   ���PUG�l�������ɿC����P�����t�v������������ǿ)��$��)?G�
L��sƾ�À�N��H����)3��5˼�nɼ��%��ޏ��	��&�"�a�I����f����Ǿ}�ܾ{��V��辉�پ��þ�ɨ�h���XvW���'Sҽ��|�Ȏ�H⎼������.}�������}��ž�   �    F)��i�D�,���.迨[����R}&�Vs/�4e2��.��%����^���m�F�I���i�v*�H쾣E���<�]Mн�G�(򜼀��P�R��1����i�����i�e�0�B1Z�w�~�^���'~��h��Y/��� ��d�w���Q��'�n��j�����A�Ț�����  ��&;�h�*��½��5�TW���L��   �   ��?��I��������ֿj��zc��8+�`x;��0F���I���E� �:�Z�*�#�|��@�׿pp���G��/�A���.1���HY���;`��܅�@f=;Ѕ�; ���㊼p�#�p ����ýFX���3�w�*���6���9��?4�&������3�����j�\&�� �޻`m<��<cH<0W��.�=��ཊDQ�c-������   �   O$Q�)ʎ���«��_�@*$�S:���L�8Y���]�Y�t�L��B:�Tb$���i����O���T�|�tpþR�p���d�v�P#z��q%<�<T�<�&<������¼��3�]��b�����J!ѽ;Pս��̽J	��+%��H~e�PK�8�g�p��;�̩<���<D?�<�x�<����kP��[���Ng������g��   �   _L\�W��Z@ÿ���7�6x,��JD�.iX��	f���j���e�DwX���D�>-��������Eſ������_�����4Ͼ;��w���7���v�0�f<8��<���<���<Psw<@��:��l����8/���X��q�Zdw�^$i��'H�&<�?���ϼ��!/< ��<&=�,=�=���<@����]�j���u���ɾ����   �   � `���dƿ7�����Z[/���G��\���j���o�ޙj�b�\�f;H�n0�$�������ȿ����d�c��� EӾ⧂�I������u�H{<T�<�=���<���<0�<ph��d���p���R\"�8�8�"w=��&0�4��P�ɼ�6���z;(�<�=r|+=��;=�{*=(��<�U���5b�ݦ���z��z;L��   �   dK\�����?ÿ���7�zw,��ID�(hX��f�p�j���e�4vX��D�z-�������Dſ@�����_����3Ͼ������C6���
v��f<س�<���<l��<�tw< �:��l�t��8/���X��q�^dw�\$i��'H�<�?���ϼ��!/<\��<J&=,=��=���< ���]������u���ɾ́��   �   p"Q��Ȏ�����迾^��($�zQ:���L�6Y���]��Y���L�A:��`$����s꿂����M��� T��unþ��p���~�v�(z��z%<�<x�<@�&<`�����¼6�3�@���a�� ���D!ѽ9Pս��̽P	��5%��X~e�FK���g� ��;�ͩ<@��<�A�<�|�<P���gP�)X���Kg��~��jf��   �   �?�JH��Ε��3�ֿر��a��6+��u;�.F�,�I��E���:��*�$!�޺��~׿5n��F����A���m.���DY�~��4`��Ӆ� �=;���; ���ኼ��#�" ��|�ýX���3�p�*���6���9��?4�&������4�����j��%����޻Xq< �<�mH<�6����=�A���@Q��*��۹��   �   �B)��i��옿W)���*�vY����z&�Pp/�b2���.�0�%����"���i�𿿠����i��r*����`B��l
<�SGн�G�4眼���@�R� .����i������i�@�0�,1Z�h�~�[���'~��j��]/��� ��n�w���Q��'�e��K����A������q��  �5�;�ޞ*�?�½��5�)T��TH��   �   T���PG����������ɿ}��6�Z����bq�T�����(����˸ǿ�%��9!���:G��H��nƾ>���|������� 3��)˼tfɼ�%��ݏ�-	�ƿ&��a�3����f����Ǿy�ܾz��W��辏�پ��þ�ɨ�i���SvW����Rҽx�|����hێ�\���t���v��J����}��ž�   �   �!�(�#��Y��(�����ڈĿ5vݿ,��[���De �����1￧jۿP�¿�n�����#6X��#��t�wҟ��jM�#D��d����v'��r�*�?��+��B���6�;�y)���Ҭ�7SؾB����v�"�|�+�ۂ.�<�*�B� �&��nH����Ҿ@����|��3�����~����'�ܪ�@��k;�����L�˼���   �   �����k��#-��]�2������qK��8ÿ�$Ϳ�<п�G̿e����h���Ϝ�����bZ��+�k �+2��Sxu����:$���a��)�4%F��Ț������=A��狾M��w��`��v�6�fP���c�
p���s���n�l�a�MM�5�3���F󾫊���ᇾ�:������j�8����F\��k����h�w��   �   �<���Fþ��M�)���P��-v�K���wR��xG��M���n���n��쉿,�r�tiM���&����A��������$2��@޽�ن��w8���:�������h6��>���Iþ����)��P��1v������T��"J��Ģ�4���$���ݽr��mM�|�&������������)2��G޽^ކ��|8��:�`���ٕ㽕
6��   �   ;:A��䋾|I��rr������6�vP�R�c�^p���s���n���a��HM�2�3����R��Ѕ���݇�9�:�/������8�ޔ��E\�~m������w�9��1m�&-��]��3��˺���M���:ÿ�'Ϳ�?п�J̿]����k��}Ҝ�$����fZ�� +� �$6��&~u�����)��b�a�H)��#F��Ś�����   �   2�����;��&���ά�|Nؾ=?����݈"���+��~.�?�*�e� �����A����Ҿw����|��3�����w���'�|��,��t;��r��L�]���M$���#�H�Y�*�������Ŀ�xݿ���]����f �����Pￜmۿ�¿Hq��3����9X��!#�y꾭՟�oM�'J��Ì��y'��r�T�?�(���   �   ,ُ�Z�+�&���a�����b����Ǿژܾw��!~��辒�پ=�þ�Ĩ�	����nW����;Iҽ��|�����ˎ�|�����w����h�}�ižn��`RG���������8ɿ���h����^��r���D�������?�ǿ�'��#���=G��J�
rƾ����������$3�+˼�aɼ4�%��   �   p ���|i�����fe���0��*Z���~�;����y������*�����<�w�?�Q���'�g��:�����A�􁨼�-��  �6;�֜*�F�½9�5��T��zI��C)��i��혿{*��J,�ZZ�.���{&��q/��c2���.���%�d��t��Rl��_����i�$u*����D���<��Kн��G�XꜼ��x�R��   �    �� Ԋ�<�#�����ý3O��q.�ɜ*�y�6���9�Y94��&�����{�+���8�j������޻��<�&�<`�H<����=���#AQ�+��2����?��H��h����ֿb��Pb�d7+��v;�V/F���I�z�E��:�n�*�R"���^�׿�o��hG����A�����0���GY���9`��ׅ�@�=;���;�   �   T�<8'<�T���¼�3�����[������ѽ~Hսޫ̽�����Rqe��?���g�P��;�۩<���<�J�<䃥<�ܵ��dP�DW���Kg��~��rf��"Q�Ɏ����M��_�P)$�R:�d�L��6Y���]�Y���L�(B:��a$������̖���N���T�f�ipþZ�p���"�v� z��w%<��<�   �   ���<���< }w<�H�:H�l����b2/�\�X���q�]w��i�� H�5��1�� ���7/<���<R*=�,=��=x��< ܛ�ր]������u�
�ɾ|��K\����o?ÿ���7��w,��ID�|hX�
	f��j�4�e��vX���D�-��������Eſ����_����E5Ͼ�����W8��pv� �f<��<�   �   �7=�	=D��<0i|<p�; V�쏇��a¼�㼄"缈A̼ t�����ur;� �<$��<č*=X}M=��[=�L=6�= J'<�����ɽ%|E��Υ��`��д8�b}�g���Y�Ͽ����^�r�%��A5�ֵ?�FbC���?�_5���%����#J��Q~ѿ����x��&<���X-��VxR�S#���A�0����ئ<n�=�   �   �^	=`��<4��<H�<����$�����ܼF��"��$��v���𼰝��������<���<-=�;=�N=�QC=d�=��#<���q!Ž&fA��������C|5�"y����zz̿�����N�"��.2��Z<���?�6S<�t72�R	#�v}��)���οڶ���s|���8�Rw �~Ũ���M�8�߽L�<�PR��H��<�%�<�   �   0�<�@�<�TW;��I�����58�.�q�����������������I���`P�tu���� u�:8��<2�=��#=:a&=�U =�><LT򼃹���5�ll���@�,���l��8����¿Gt��T	�2	�0`)���2�"6�4�2��5)�����}	��3�_�ÿ#{���ko���.�c��螾�A�)fнν.�0`��(��<H��<�   �    ��;�#ܻ�RռG�c���½���d��&E�����_�j �k]۽�˭���v���`�=��w</�<�t�<	�<���;H�Լ�p��Df#����O1ؾ�q��HY�rᎿ)ֳ���ٿ׳��~�����F$��'��$���v��UR��Y�ٿ�F��S����[�ai��gܾ&����5-����U��.��X�+<�[b<�   �   D���R�$����}�ѽi3�2Q.��jL�f�c�I(r��v��+o�u�]�&D���#��% �?b��¼d�4ټ�v���(<x^< vm;t߶�L슽����	r�m|���
�@_@��~�Ti�� t¿���W���j.�Ng�(����r�
�{���������d:���W~��-A�����T��~�x�$l�s������������:`�/��   �   �aP�y
�������4���g�F���c���z����O��*n��l���y����?��,d��g\��;(����򻖽ڲ���k�@�ں��0����zkb�Te��I��t���?뾕$�F�Y�W�������sĿOpݿ���4��6� �j��
����ۿOÿU⦿*i��lY���#����\䠾P�M��3�N7}��2Ἠ�@��B��RѼ�   �   y�����@S�"J��m��MwӾ;���f�T��"K�`�8��,���;Tx���=��GvG�p�	�""���>����L�8뛼<�2�A��~V �Ty��Si���{�~�3��	e�䋿���~U����ɿVԿMX׿�Pӿpnȿ&������\���e�b�#.2����P���"�����!��%��H�C�pjɼ�������jd��   �   }���da�<����˾Q���iR���+��<��vF���I��lE�)):�}�(�J`�����Hž>*���W�a��;���vlE�\�ּE��ƚ�Ȇ����AE������gӾ�<�E~6��`�x����s��J��q|��$��yȪ�����=ޓ��P��y]��3�t@��{о������B�E��!���<��TȼĞ���]��⿽�   �   �e\�Y���c�׾~X�N,�l�K�}vg��}��M���h��ݱ����z���d��~H��)������Ҿ˲���V�3
���75��ܼ���h�=�ު�Q��`\�������׾�U��,�m�K�rg�%}�LK��|f��������z��d��{H�%�(�����Ҿ)���V��
��죽N55�T ܼD��О=��㪽~���   �   0����kӾB?���6��`����� v�����
���&���ʪ��¡�N����R���
]���3�_B��~о������B���ｵ���N��lȼ�����]�yۿ����'^a�,����˾b���O�ć+��<�orF�ޥI��hE�~%:�-�(�i]�Ė��1Dž3'��y�W�!��񉱽�gE�$�ּH�����X̆�T��^FE��   �   �l���}�v�3��e�拿!��X��i�ɿ
Կ�Z׿Sӿ�pȿB���Á��肊���b�02���f�������u�!�{'����C�$fɼ�������d���������9S�F��<h���qӾ#��c�����G�$�2�����_�;_t���:��FqG���	������>�`���X L����2��E��*Z ��{���   �   TC�$�M�Y�&�����vĿ�rݿQ��37���� �m��V����ۿ
ÿ�㦿[j��IY���#���뾩堾��M��5�8}��/ἐ�@��kB�d@Ѽ�UP�k��n��L�4�Q�g��������n���uJ���h��d���ɒ���;���`��6\��6(�������~��8�k� Xں �0����qb��j�ͮI�Hw���   �   ��
��a@��
~�k���u¿��⿵����/��h�f������
��|��b��"���j;��nY~��.A�g���U��·x��l�����P������?�: H/�H����$�C��3�ѽ�-��J.��cL���c�� r��v�P$o���]��D�L�#��  ��Z���d�hټ��u���(<^<�fm;�涼�J���r�&���   �   hs�KY��⎿�׳�Y�ٿõ������� H$��'��$�Ά�4���S��Q�ٿjG��䘏��[��i�ihܾ����:6-�����S�P����+<�pb<0�;��ۻ�<ռ��F�����X�½��=���?�B���Z�� ��T۽�í��wv����`�=�X�<x7�<4y�<�	�<@��;��Լ;t���h#�f���3ؾ�   �   �,���l��9����¿�u뿖U	�
�a)���2��6��2�66)�$���}	��4���ÿh{���ko��.����螾�A��eн �.��M��8��< ��<��<�L�< �W;�mI���켰*8���q�����x�����X��� D��0VP�l��� C�:@��<¬=��#=2b&=RU =�6<�[򼈼��T�5�n���B��   �   \}5�e#y�o��[{̿���.���"�/2�b[<�B�?��S<��72��	#��}��)���οǶ���s|�e�8�w �Ũ���M���߽��<�p@����<�*�<�a	=h��<\��<�<p{���t��<�ܼ�?�"���$��p����ē���n����<D��</=�;=PN=~QC=H�=�#<(��$Ž hA�M���=����   �   ��8��b}�ۻ����Ͽr���N^���%��A5��?�HbC�t�?��^5�p�%�n���I���}ѿ�����w��s<����x,��wR�P!���A��~��<ܦ<��=�8=�	=���<Xm|<p�; O仈���|`¼�~�P"��A̼�t��h�@kr; �<X��<Ȍ*=<|M=��[=��L=j�=�@'<�����ɽ{}E��ϥ��a���   �   �|5�P"y�����z̿�����(�"�Z.2��Z<�d�?��R<��62��#��|��(��ο���fr|���8�rv �,Ĩ���M�A�߽��<��3��`��<�,�<6b	=T��<��<H�<0y��$t����ܼt?�"���$��p���𼰓���n����<d��<8/=;=�N=RC=&�=X�#<��"Ž�fA�t���	����   �   �,�p�l�I8��+�¿�s�zT	����_)�2�2�V6�X�2��4)�����|	��2��ÿz���io�l�.� ���枾aA�Ybн��.��5�����<��<@"�<tN�<��W;xkI����X*8���q������x��	���T���D��,VP�l��� H�:���<*�=n�#=>c&=�V =�@<T򼕹��$�5�gl���@��   �   7q�,HY�����tճ���ٿ����������E$��'��$�Ԅ�j��eP����ٿE�������[��g�eܾ.���
3-�^���M�������+<xyb<��;p�ۻ�:ռ�F�O����½���,���?�:���Z�� ��T۽�í��wv�z��0�=�H�<L9�<|�<x�<p�;�Լ#p���e#�*���0ؾ�   �   D�
�"^@�V~�Zh���r¿I�⿍���b-�&f������4�
��x����������8���T~�+A�����Q��?�x��h�l�����������:�/�x�����$������ѽ�-��J.��cL��c�� r��v�R$o���]��D�P�#��  ��Z����d�Hټ �u���(<*^<��m;�ٶ��ꊽ���tr�\{���   �   �=�>
$�w�Y�.������rĿMnݿg��2��� ��g��i��O�ۿ�ÿ>িYg��_Y�"�#���tᠾ��M�?-�,}���`�@�\B��:ѼnSP���� ��
�4��g�󪌾����e���qJ���h��e���˒���;��`��5\��6(�������V����k�@�ٺ�I0����gb��b��I�-s���   �   6g��,z���3�~e�{⋿���bS��g�ɿ�Կ�U׿�Mӿ�kȿ�����}��I����b�'+2�7������R���x�!���,�C� Vɼ������ d�����Q��49S��E��!h���qӾ��c�����G�%�5�����b�;`t���:��3qG���	�<���>�P���(�K�p᛼�2��=��WT ��w���   �   �����dӾ�:��{6��`��􃿥q������y��|!���Ū�����ۓ��N���]���3��=�wо;󒾔�B�3�ｪ������ȼ����"�\�"ڿ�,���]a����x˾H����N���+��<�mrF�ߥI��hE��%:�0�(�l]�ǖ��1Dž.'��V�W�ޓ�
����dE���ּ:�����Ć�3��>E��   �   \\�ۛ����׾>S��,��K�Jng��}�I��$d��=����z���d��wH���(����:�ҾI���V�
�1壽)5�L
ܼ(��p�=�Cܪ�����_\�d���n�׾xU��,�f�K�rg�#}�LK��}f��������z��d��{H�)�(�����Ҿ����V�I
�@룽 15�\ܼذἦ�=��٪�g���   �   ��eYa�����˾}���L�p�+�<�nF�ˡI��dE��!:�z�(�Z����5?ž#����W����ˁ��\ZE���ּ�2��r���ņ�'��AE�����qgӾv<�:~6��`�u����s��I��r|��$��{Ȫ�����@ޓ��P��|]� �3�s@��{о����{�B�%��N������@ȼ؅����\�4ֿ��   �   �������S4S��B��3d��mӾ�{�`����pD�����������;�o���6���jG�T�	�@��(�>��㴼P�K��ۛ��2�0?���U �y��,i���{�u�3��	e� 䋿���|U����ɿWԿPX׿�Pӿsnȿ(������^���g�b�$.2����@������K�!�F$����C�\ɼ�������d��   �   �KP����P���4� �g�L���k�������nE���c��7���̍���6��K\����[�v0(�^��������؜k� ٺ�0�p��(gb��c�l�I�^t��y?뾋$�>�Y�S�������sĿOpݿ���4��8� ��j������ۿRÿW⦿+i��oY���#����D䠾��M��2�3}� 'Ἠ�@��TB�|1Ѽ�   �   0u��@�$�����i�ѽ5)�fE.�n]L�
�c�8r�\v��o�3�]�D��#�z �dQ��6�d�`�ؼ@�t�P)<x?^<��m;�ն��ꊽ���	r�N|�� �
�6_@��~�Ri���s¿���X���j.�Ng�*����t�
�{���������f:���W~��-A�����T��A�x��k����*��0����˸:`�.��   �   `7�;@�ۻP+ռ��F������½]��t���:���bU�� �?K۽M���Jhv�L��ȭ=���<�G�<8��<��<p �;P�Լ�o���e#�p��61ؾ�q��HY�oᎿ(ֳ���ٿ׳��|�����F$��'��$���x��WR��Y�ٿ�F��U����[�`i��gܾ����5-�����Q����X�+<��b<�   �   &�<�T�<�X;�RI�d��6!8� �q�%����r����Į���=��&JP��`�����@Z�:H��<V�=n�#=Lg&=BZ =`K<�O�ɸ��ՙ5�Wl���@�,���l��8����¿Gt��T	�4	�2`)���2�$6�4�2��5)�����}	� 4�^�ÿ&{���ko���.�^��螾�A��eн».��G�����<D��<�   �   zb	=T��<���<@�<�_��l����ܼ:�. "�R�$�hj��𼨇��PA��8<t��<<3=�;=�N=�TC=��=�#<���!Ž	fA���������@|5�"y����zz̿�����N�"��.2��Z<���?�6S<�t72�T	#�v}��)���ο۶���s|���8�Pw �xŨ���M���߽N�<�0F�����<�+�<�   �   x�=�=�C�<p��<(W"<@p�:���0����?��5�P{󻀈���� <�Z�<���<dC)=b`R=�Wp=D�|=��o=xTA=dG�<��4�&X�����xu~�˧Ǿ��Z!J�k8��G��Ƀ˿)����)�2�*����B;�7�Z�̿aL�������0M�H� �ξ�ᆾ��"�k]�������:,ڰ<8�=�   �   �=���<8��<P*Q<�Z; ����3Y�h5��$��T%���r����(� �K��/<���<�m=��>=8�`=��p=�g=�<=�I�<�A)�!����h�{iy���þmr���F�� ��:J���Hȿ�����������4����������u�T2ɿ/s���S���I�.���ʾ���u&�ﻧ��V ����:�s�< E�<�   �   ���<�U�<X�<�酻�Չ��7�1!�P�@��NQ�.�Q�T�@��#� }߼�(X�@J;�[�<��=~!1=H�L=��N=:�.=�@�<�~	�B$n�����j�d&������<��y��[��mܾ�}�޿Di�����jA����)�v��\V��Z*߿�e��Y+��?{���>�
�b��&x�vm��|����`-;��<���<�   �   ��<< �f8�C}�lu��rT��~��*��Ž~8ӽ>ս�2˽�����a��*�_���
���R���;d�<8d=��#=X=�<࠼��GN��0���S��N������,�1�d��ݐ����
�Ϳ,��������45�~��%<�����Ϳ���4���e��C.��������P_�����Y���_����;8mr< �<�   �   `I����ټ2ZM��Μ�7�Խz?����V�.���9���;�S�5��%'������N�����l�������P�V<h��<9�<�j�<@�P�@�'��ɽ� 7������ھ�v���J� р�휿ʷ��gϿ ��ȏ�g�;�k�8�οv���w������5K�%4�"hܾr5���?��B޽ԁ[�l;�� ��:X�<�`�;�   �   ��� ����ǽ>7�h�3�p[��}��=��sw��ܭ��H���\���,s���M��9$�����B��^�7�|b�� 5t;0oe<�lR<��Ǻ�����r��P����u�+����T*-��\�|	��]���I0��{BÿS`Ϳ>�п��̿K¿���dx��^,����[���,�	|�'鸾�Sy��G��g����&���Y�@���jۺ8cZ��   �   "T��2&⽘L#�j�Z�fJ��5���뾾u3Ҿ�0޾�ᾱSܾ9�ξ�Ĺ�%ڟ����sK��z�U�½�n^������a� �;��Ժ�W����s�T�'�D�O��M�ӾFH��m6�l�_��ڃ��Z������u����;����񡿕���ʐ]���4������ѾD>����D���k������:#��V˻���l��   �   :n�I�-��r������CǾa��
��08����� �I���^��W���Q����Ř��|e�m1!��	Ͻ��h�p\ѼpY �P5����w� h*�[b����֍f������oྨ��Nm2�(�R�Жo�����)��f����K�l��P���/�B�Eܾ�?��j�a�ж��y���,��l��X����n����R*���   �   �(�w�cV��Iܾa��!�Ws8�NJ��U� �X��T�P!H���5�����T�0#־�㣾lSm��z ��ƽXNV��\�����--�4�ؼ^�j�3�ӽ��(�w��R���ܾF^���!��o8��J��U�C�X��T��H���5�.���R��־�ࣾ&Om��w ��ƽTIV��X��`��9-��ؼ��j��ӽ�   �   �f�����s�]���p2���R�ǚo��������2+��h���󁿲�l��P�	�/�D�9HܾB����a���T|����,�@m��8��8�n�4���$���f�5�-���r������>Ǿ�����4�L��Y ����[�0U�;��h������we��-!�mϽ��h�TѼ�S �`>��x��n*��g�����   �   /"���Ӿ�J�xp6���_��܃�]���������>����~�V��t���V�]�э4�J��1�Ѿ�?���D�� ��������3#��8˻���b��M����WG#���Z��F���0���澾5.Ҿr+޾���xNܾ[�ξD���X֟����jnK��v�+�½�e^�, ���a�`�;��Ժ8a��d�s�?�\�D��   �    .��ۖ��,-��\�5��I���\2���Dÿ�bͿg�п��̿dM¿{���y���-����[��,�(}��긾�Uy�	I��h��|�&� �Y� ���@�ں FZ���x���w�ǽ@2�x�3��[���}�}9��@s������9�������Xs���M��4$����^<���|7��T�� }t;�we<0lR< NȺ�����v��q��h�u��   �   �ھ�x�$�J�lҀ���˷��iϿ'��ԑ�i�� Ὸ�ο����x��n���~K�5�qiܾO6���?��C޽T�[��9��@-�:��<���;���8�ټ�MM�}ǜ�Z�Խj:���V�.���9���;�U�5�) '�����¨����l�\r��G����V<���<�;�<Di�<��P���'��#ɽ$7������   �   ���^�,�W�d��ސ�4����Ϳ�迕������6�F���=��6���Ϳ����4���e��D.�a��q����_�4���Y���]�� �;@yr<`�<(�<< ��8@ }��j�lfT�gw��N孽��Ž�/ӽw5սW*˽񥵽tZ��Ŀ_�v�
�H�R�0?�;��<�g=��#=|X=|�<�����LN��4���S��P���   �   �����<�Jy��\���ݾ���޿�j��8��B����*����$W���*߿f���+���{���>�5
���%x�Om�9|�� ��I;x�<Ԍ�<���<�_�< �<P����ŉ�|%�'!��x@��CQ�V{Q��|@��Pk߼�	X� �;�f�<��=�$1=,�L=��N=�.=P=�<p�	�0)n���%�j�'(���   �   Rs���F�����J��[Iȿ���p��$��p��@5�ƃ���� ��u�d2ɿ-s���S��߅I������ʾ����%�㺧�U � �:�w�<LI�<@=\��<���<�9Q<`�Z;�ظ��Y��*��<�����hh��(�(���J��/<X��<6p= �>=@�`=�p=�g="�<=DF�< M)�<���mj��ky�,�þ�   �   z�"J��8�����+�˿�����*)�B�,����(;��6��Y�$�̿ L��'���0M��G��ξᆾ��"��[��^��<�:Pݰ<��=��=.�=�E�<H��<�Z"<���:���P����?�5��{������ <�Y�<\��<�B)=�_R=�Vp=(�|=d�o=�RA=\C�<��4��Y��Ħ��v~���Ǿ�   �   �r�ϧF���CJ���Hȿ���������Έ��4�"��$�����t꿉1ɿsr��RS���I�F����ʾ����$�t����R � 5�:�y�<K�<�=p��<���<�;Q<��Z; ָ��Y�\*�������Lh���(���J�/<l��<Np=D�>=j�`=`�p=X�g=�<=�H�<XF)�����|i�,jy�2�þ�   �   ����<�"y��[��ܾ���޿�h�����@�p���(����U��)߿ud��Q*��r{�&�>��}
����dx�`k��y��L���w;��<��<l��<�a�<��<𪅻0ĉ�P$�&!�Vx@�|CQ�${Q��|@���$k߼�	X� �;g�<�=�$1=��L=l�N=P�.=�A�<p~	�L$n�����j�K&���   �   B���,�S�d�ݐ����Ϳ�}������^4����e:��S���Ϳ^���2����e�&B.���������_�����U���R�� �;`�r<�<��<< Є8}��i�peT�w�� 孽N�Ž�/ӽY5սF*˽䥵�iZ����_�P�
���R�pA�;��<�h=!�#=tZ=��<����FN��/�9�S�"N���   �   �ھ�u���J�0Ѐ��뜿�ȷ�-fϿs����e�3�e�G�ο���)v��(���� K�02�eܾ3��b�?�y=޽>y[��,�����:0 < ��;������ټBLM��Ɯ���Խ0:�޵�9�.�u�9�{�;�N�5�' '���������j�l��q��`B����V<���<H@�<tp�<�bP�t�'��ɽ�7������   �   �)��̓��(-�&�\�L����.���@ÿH^Ϳ�пs�̿VI¿���zv���*����[��,�z�渾�Ny�D��a����&�`�Y���� Nں :Z�~��|�����ǽ�1�,�3�b[�Z�}�l9��3s������5�������Ss���M��4$����+<���{7��R��`�t;��e<H|R< �Ǻ����6p�������u��   �   ����Ӿ�F��k6���_�]ك�>Y������[����9��S쪿\������_�]�ӈ4�C����Ѿ>;���D�������輠#��˻����_��L�����F#���Z�hF���0���澾'.Ҿi+޾���sNܾ\�ξE���W֟����_nK��v���½�d^�������a�P4�;��Ӻ�N��~s��콨�D��   �   W�f�1���blྦ���j2�4�R�g�o������&���c���Z�l�P�^�/�c?��@ܾ<���a�~���r���,��Y���r�`�n�R��6#��Ze潽�-�*�r�h����>Ǿ̳�����4�H��W ����[�1U�=��h������we��-!��Ͻ0�h��NѼ�C ����x�w�b*��^��!��   �   6�(�� w��O����۾�[�&�!��l8�	J�6U�h�X�
T�H��5�����O��־�ܣ��Hm��r ��ƽ�<V��C��H���-��}ؼؑj��ӽ�(��w�ZR��]ܾ8^���!��o8�J��U�C�X��T��H���5�2���R��־�ࣾOm�fw ��ƽGV�TQ��X� -�d{ؼ�j�I�ӽ�   �   �`�E�-�p�r�X����:Ǿ0��N���1���	 �Ď�~X�-R�Ȗ羥�������>qe�V(!���ν�h��=Ѽ�, ���h�w��c*��`���f�f�c���boྙ��Bm2� �R�̖o�����)��f����O�l��P���/�B�Eܾ�?��?�a�����x��ȗ,�@c��`{���n�@��- ���   �   �H��C�C#���Z�HC���,��D⾾O)Ҿ8&޾1��Iܾ#�ξf����џ����gK�Hq�O�½dW^��込`a�0Z�;@�Ӻ$N��
�s�콰�D���(�Ӿ7H��m6�c�_��ڃ��Z������v����;����񡿗������ː]�4������Ѿ4>��k�D����������!#� ˻h��[��   �   �{������ǽ�-�M�3��[���}��5��.o��w���	�������� s��M��.$�����3��nn7�H=���u;��e<��R< LǺ����!q�������u��*��ؔ�I*-��\�y	��\���I0��{BÿT`Ϳ@�п��̿�K¿���fx��_,����[���,�|�鸾oSy�jG��f����&���Y�@6�� (ں,Z��   �   ����p�ټ8CM�������Խ�5�����.��|9�W�;�)�5�4'�v��ػ�ß���l� X��ﹻ�W<\�<�I�<�v�<�FP�$�'�|ɽ 7������ھ�v���J��Ѐ�휿ʷ��gϿ"��̏�g�?�m�9�οw���w������7K�$4�hܾe5����?�B޽`[��3�����:�<0��;�   �   ��<< ��8@}��a�p[T�q��!ޭ���Ž�'ӽ�,ս�!˽�����R��b�_���
���R�Ћ�;�+�<�n=� $=^=���<Ї��^EN��/��S��N������,�+�d��ݐ����	�Ϳ-��������65�~��&<���翀�Ϳ���4�� �e��C.��������)_�����X��HZ��`�;�r<p�<�   �   4��<�f�<��<����췉���!��n@�N9Q��pQ��q@���XW߼��W��8;`u�<>�=*1=�L=��N=0�.=PF�<�v	��"n���c�j�Q&������<��y��[��nܾ�}�޿Di�����lA����)�v��]V��Z*߿�e��[+��@{���>�
�_��x�Nm�.|��d�� V;(�<Ȑ�<�   �   =��<���<HCQ<��Z;�����Y��!�����`���]��hk(� �I��&/<��<,t=��>=v�`=��p=��g=��<=�L�<�=)�Ƣ���h�diy���þjr���F�� ��9J���Hȿ�����������4����������u�U2ɿ/s���S���I�.���ʾ���b&�����V � ��:lw�<�I�<�   �   �%�<�6�<0ݠ<�s<� #<��;@�;��7:�r: DU; ��;`0j<� �<܊=R�,=��T=@�w=���=Rč=�q�=(Vj=?�=Ȓ<���R�ý�7�*����ݾ���M������	���]����ҿ����^��l��f���ҿdܺ�ǟ�၃� �O��r����H)���L�����K-����ļ@�:�<��<�   �   ��<`+�<0�<��.<�f�; Ŕ� 鋻 ֻ�Lܻ���� �B�S�;��<l{�<H=�hA=�g=��=(׈=���=�Jf=�=P�$<~�#���3��ӑ���ؾ�����I�{[���o�� \��5'ϿF�ῂ��>�������uSϿ·�V���;�� 2L�4��p�߾� ���H�c��0z��J���;�:���<�C�<�   �   �w�<�]<���; }
��-�\����ʼt���\������¼���������"�;�k�<d=��6=D�\=�s=T�t=(�Y=��=�9<����Ȱ���(�Ή���@;���L�?��t��ڔ�0���]Rſx-׿ڔ⿁u��u�p׿'DſI���<���Au��wA��-��Ӿ(ِ��;���ݽ��b�@A��@]9;(*u<x<�<�   �   �=< ��9�.9��EǼ����8L��v�T���������V��Z�c���-�X�ڼH���j<��<��=�~@=�P=N�C=n�=��T<�꽼K皽�`��9y�������T�/��`��툿�Р��ߵ�`ƿP�пbԿ]�пjƿ-���ٝ��8󈿍�`�l�0�i��h��Օ��0�&��*½��>��q� �;��U<8�f<�   �   �ݐ�`������,vj�����v�ŽБ�qM ��=�a��7��M���ƽ뚽�U�x�����ؚa<P��<K�=ߚ"=�=�.l< ��6h��o�.�X�ϣ�V��x?�(�F�VKs��!��.��o߰��>���W���鹿@Q��^r��j�����r�'OF��x�+�ޕ���a�5e�c��N��`����; �<p��;�   �   ����=�����ѽ_��=%�p�>�
3R�/�]��`�"�X�8,H���/���v���8����;�LՓ�`�;8��<ȱ�<�5�<x�t<�<��D��ҽ��3�+щ��Dľ�)���)��zP�G�u�Jn��tQ��t�����������������0t��O�?�(�j����þT����k8�vn��aq�l�Ƽ�Vs��ڟ;��\;P�ػ�   �   x�I�w���|���z�%� �Q�/|������#�������@��c���Q���
'���_k��>����[5ǽ�2p��ؼ@�����]<T��<��b<��X�<	�`j��?c��^�l�G~ؾ���,��xK��:g�i�|��L�����݄��Y{�+3e�EI���)�V�	�T\վ�v��2�[�3R�/���"�0RT��Q$:@/(;���� <���   �   =3��
��!I7��"r�L������pϾPt�5�`��j� i߾/Nɾ\ƭ��8��Z`�t�$��*޽Ɵ��`��P�����	<0�.<@]�: V���0c�0�Խ�*��%y��A����ܾI����!�&p8�uJ��U�`�X��-T��PH� 6�I�����:׾,��S2p�@^#��ʽ��Y�$n����@� �N;�Q�l#����9��   �   &���!9�� ���R���о����=����~#�%&�j�"���Ԧ
�Z?�"ɾ���E�q��{+�z߽�]~��S�0����;@O];pJ%�ڬ�~"�����]9�����N��|о�{���:����{#�&�z�"�*�b�
�;�ɾ�����q�gx+��߽�V~�K�@������;�-];�[%�ڳ��'���   �   ��*��*y��D��*�ܾƓ���!�Gs8��
J�BU�X��0T��SH��"6�ZK�����=׾�.���5p��`#���ʽ(�Y� s��@�@� �N;�����R�9�Y-��)��&D7��r���������ϾIo��.��h�wd߾ Jɾ�­��5��e`���$��$޽v����������
<��.< �:�`���8c��Խ�   �   �^�Vş���ؾK��|,��{K�>g���|��N��ɀ��D߄��\{��5e�kGI���)���	��^վ�x��ޏ[�T�l1����"�`UT���$:`X(; f��L.���{I�/���s�����%�9�Q�a|�ԭ�������g<��R��������#���Yk���=����.ǽ�(p��	ؼ@����]<���<��b<��X�4�	��n��}f��   �   {Ӊ��Gľ�+���)��}P�V�u��o��3S���u�����2��C���
����2t��	O�ʕ(����q�þ����Cm8��p�>dq�0�Ƽ`Ns�P�;�-];��ػ���8�=������ѽή��
%���>��,R���]�x`�ΫX�M&H�B�/�p�����V2��p�;�lœ��:�;���<���<�5�<(�t<XL�0D�[ҽ'�3��   �   dѣ�R��WA�i�F��Ms�#�����᰿v@���Y��~빿�R���s��r���8�r�~PF��y��,�喦�Xa�f��c�� ����� �;��<���;0���|���l���jj�"�����Ž���H ��8�������3D꽽�ƽ䚽��U�����Q����a<Ċ�<��=��"=��=�%l<X���n�<r���X��   �    ���@���/��`��Ҡ�)ᵿhaƿ��пYcԿ��п�ƿ"��������󈿍�`�(�0���{i��F�����&�Y+½��>��q���;�U<(�f<HN< Q�9H9�D5Ǽ���-L���v�vM��@�������O���c���-���ڼp��x�<���<��=��@=ĭP=��C=~�=`�T<��yꚽ*c��<y��   �   �B;����?��t��۔�/���gSſ�.׿��xv濲v�1׿�Dſǽ��u<��jBu��wA�.�5Ӿ?ِ��;�j�ݽJ�b�d?�� q9; 1u<�@�<\}�<H]<#�;`&
�8�-������ʼ��뼜K�����(�¼�Ђ� L���T�;\v�<�=�6=��\=p�s=�t=��Y=e�=�9<l���˰���(�-����   �   R�ؾf����I�\���p���\���'Ͽ������M��N�ΎSϿ5·�c���;��2L��� �߾� ��0H�p�ｂ.z��G�� g�: ��<,G�<���<�/�<`�<��.<p��; ے��ȋ��\ֻ�)ܻ�p��  �5�p�;0�<��<�=�jA=<�g=l �=T׈=���=�If=f�=|$<��������3��ԑ��   �   �ݾ���p�M����O
���]��ćҿ��7��a��V��;����ҿ ܺ��Ɵ�������O�r���㾒(��āL������+����ļ�L�:���<��<�'�<�8�<�ޠ<�s<#<@�; �;��7: .r:�EU;���;�/j<D �<d�=��,=�T=��w=(��=�Í=q�=�Tj=��=`�<p���ý$�7�䮔��   �   D�ؾ�����I��[���o���[��'Ͽ������O��]���RϿl������f;��1L�T���߾����H����,z��C�����:T��<4I�<l��<h1�<��<(�.< ��; ���0ŋ��Zֻ�'ܻPo��  �5`q�;d�<4��<�=�jA=f�g=� �=|׈=���=fJf=S�=��$<��󾽄�3�ԑ��   �   �@;�����?�tt�[ڔ������Qſ�,׿�⿏t��t�d׿CſH���(;��:@u�vA��,�Ӿ�א�V;�.�ݽ��b�(8����9;`:u<�D�<܀�<X$]<�-�;�
� �-�$���Pʼ��뼨J����鼬�¼�Ђ��J���U�;�v�<�=,�6=�\=�s=��t=�Y=3�=П9<t���Ȱ���(������   �   7���e����/��`�-툿�Ϡ��޵��^ƿ�п�`Կ��пƿԅ������򈿃�`���0� ��f��"�����&��&½N�>���p��;�;	V<X�f<�W< ^�9�9��1Ǽ����,L���v�M����������O����c�P�-�$�ڼ���`�<���<+�=d�@=ܮP=f�C=�=@�T<�罼v暽K`��8y��   �   Σ���}>�ޒF��Is�� �����ް�X=��WV��^蹿�O���p�������r��LF�w��'�s���C
a�\b��^�����pi��C�;h�<`��;P���t���6���hj�C�����Ž��罌H ��8�j��o��D꽣�ƽ�㚽��U�0���N���a<���<O�=��"=��=�7l< ��4e��n���X��   �   �ω�Cľ�(��)��xP���u��l���O��wr��%������������-t��O���(�r����þܪ���g8��h�bXq���Ƽ �r���; s];0�ػ�����=�[����ѽW���
%�I�>��,R�}�]�V`���X�@&H�6�/�c��k��.2���;�<ē��B�;���<��<�<�<(�t<�.��D��	ҽ��3��   �   �^������{ؾg���,�%vK��7g�O�|�K��C}���ۄ�:V{��/e��AI��)��	��Xվ�s��d�[�{N�5)��zw"�@1T� ?&:@�(;C��'���xI�Ϡ��A�����%�«Q�|����������X<��I��������#���Yk���=�Ҹ��.ǽ (p��ؼ������]<���<c<@RX�nz	�Eg��0a��   �   �*��!y�?��ˮܾS��f�!�tm8�tJ��U��X�D*T�RMH��6�*F�J��>6׾�(���,p��Y#��ʽP�Y�t[���L@��O; ��l��д9��+������C7�Ir�m���Z���Ͼ0o���$��d�td߾�Iɾ�­��5��V`�z�$��$޽������`u���
<h�.< �:�K���)c���Խ�   �   �����9�����K���о�w��\8����x#�&�m�"�5���
�6�ɾ����q�_s+��߽J~�06��:��P�;��];07%����� �������9�����N��Nо�{���:����{#�&�{�"�,�b�
�;�ɾ�����q�Jx+�.߽�U~�G��i��@ť;@�];�5%�T��Q���   �   [(����	@7��r��������~Ͼ�j������2��k_߾EEɾs���,2��
`�B�$�M޽������;��p$
<P�.<@�:�M��-c���Խ]�*�%y�^A��ʱܾ6����!�p8�nJ��U�a�X��-T��PH� 6�I�����:׾
,��;2p�^#���ʽƵY��h��`�@�@�N;��������9��   �   .sI�����q���3�%��Q�C|�X�������)8�����p������
Sk���=����,&ǽXp��׼@��� ^<���<�c< HX��{	��h���b�^�9�~ؾ���,��xK��:g�f�|��L�����݄��Y{�-3e�EI���)�U�	�P\վ�v���[��Q�Z.���~"��DT� �%:@�(;�9��� ���   �   �����=�ݶ���ѽ��� %��>��&R�C�]�� `�:�X��H�N�/������*��z�;�(���p��;��<���<|C�<�t<(-��D�aҽK�3��Љ��Dľ�)���)��zP�@�u�In��uQ��t�����������������0t��O�?�(�i����þH���hk8��m�`q� �Ƽ�s��	�;�x];0�ػ�   �   `����������_j�ĭ��K�Ž܀�ED ��3��������:��|ƽ�ۚ���U�|������0�a<,��<��=�"=t�=x>l<���e�`o�֋X��Σ�9��o?�!�F�PKs��!��.��p߰��>���W���鹿BQ��_r��l�����r�(OF��x�
+�Օ���a�e�ab��F���v��5�;p�<pƹ;�   �   �^< �9��8��%Ǽ��n#L�vv�G��������I����c���-�Tmڼ����<���<}�=x�@=�P=��C=T�=��T< 潼y暽�`�`9y�����؈�J�/��`��툿�Р��ߵ�`ƿS�пbԿ_�пlƿ/���ٝ��9󈿎�`�k�0�h��h��̕���&�k*½Z�>��q�@,�;0V<X�f<�   �   `��< +]<�B�;��	���-��u�� �ɼ��뼰:���鼬�¼Ŀ��P��А�;��<�%=<�6=t�\=��s=��t=��Y=6�=x�9<���\Ȱ���(������@;���G�?��t��ڔ�1���]Rſx-׿۔⿂u��u�r׿(DſJ���<���Au��wA��-��Ӿ ِ�t;�N�ݽ �b�T>��`~9;@6u<�D�<�   �   4��<$2�<|�<��.<�; o�������?ֻ 
ܻ0O��  �6���;\$�<Ј�<5=�mA=<�g=�!�=�؈=���=FLf=4�=�$<������3��ӑ���ؾ�����I�z[���o�� \��4'ϿG�῅��?���� ��wSϿ·�V���;��2L�2��n�߾� ���H�<�ｪ/z�$I���[�:�<�G�<�   �   pƪ;Б�;�;C;�k�: ~u: ݅:@�
;���;��<��P<썚<���<-�=,v2=Z�W=�wz= �=l��=��=v��=���=@�Q=�Q�< D��a�`���"Q�	W���K���GB�(Jn��\��g(��7򭿇g�������g��F���=T�������mo��C��"���?��@�h��������U��Ѽp� �F9`��;�   �   � �;`�D; wg:�,���+� �T��d6� v��`�
;��;�gS<p��<���<�)= �E=��j=h��=T}�=Z��= ��=p �=D7P=^�<��ûl,Z������L��Y����ݾ
��>�6Bj�����&���b������0]��H��ң���M���Ak��w@��E��.�f뤾G�c��z��ط�^;N��NƼ��� ��9`\�;�   �   ���:@���p߷��6!�H,^�,����!���ې�`��X=��\�� E8;(�N<��<K�=�;=n�c=N��=@��=�ӊ=�=��K=�c�<��a��2F��V߽2�@������Ҿ*M�!65���^��4���ݔ�S���B������L���&����Ҕ�N��["_��T6����j׾�A���U���
�0���018��ꧼ0Qû�ޠ:@U;�   �   �;�`���*�� �ͼx���� �j{4��?�a>�dU1�l}�@㼸���@(!��C<���<�_ =D�L=#k=,w=k=��B=�w�< ��9И'�Pƽ��-��;��خ���9�B&�Q,L��q�<؈�U����ԝ�ݓ��{���+i��������p�1L��&�1U�Y�þv1���+?��6�������8���t��D:� Q�: 	�:�   �   X6-�tñ��i���D���z�3���"��ҥ��1���n�����\Km�8�%�T����8�|<x��<�].=P�J=�,N=�R4=���< ��;�)�����W�Йj��u����㾨��O�4���U���r�Y�x<��~���5�������X r�g�T��4��o�rY�SY���3r�]�"��˽�#e�|�׼X�� ��9���: ���   �   `����5!���q�t���wν{���9�8��3��������	����W:���&���&�����p�;���<�=+�%==�#�<��<HѴ��ф��:��>�D�턎�ů��;%��tl���6�zP���c�tvp�L�t�
�o���b�r�N�[N5�������B���, ��|$G���l����!�8�v�����@�M; c�9���   �   Tz�5���������l��l�:�"�T���h�zt� �u�+�m�8�[��B��P"�*����|��Pg��ܼ ��$τ<(��<��<���<��<<@S��WE�	ý2^�\�g�*����o;f6������+�*;<�עF�?�I���E���:��)�K|�f��y�Ⱦ$D��B*a�pU�k½X�V���� i{��^�;p͐;�ci�(��   �   l�u�������4�M�`�⭅��x������*ȯ��뱾B�����"����Vw��H�<t�%�ؽQK����@�Ի�u<<@j�<D��<�OS<�㧻������ĉ��05��y��q��3zɾ"L�ln�-�����\] ����R��6��
(�m�¾�.��KAk���'���ܽ ΀�(o� y˻@��; �<@vp;�K(�D���   �   4$��q����<��w����������Qо�\�9��V��R��߾�ʾܧ��&R��r�b��'��p�pf��^g�`����O
<0:u<��H<�:t���"'J�-����?�<�!�v�\���њ���Mо3X侞��&R����߾#�ɾ����uO���b�|�'��k彉b���a� t���W
< <u<��H< h:졤�@.J��   �   ���45�ޱy�u���}ɾbP��p��������_ �������B���+�c�¾1��Ek�}�'���ܽ�Ѐ�w�Ћ˻���;��<@�p;0=(�~��0�u�6��\��x4��`�ê��?u������Eį��籾�����������Qw�x�H�sp�&zؽ�F���x�@\Ի�<<4m�<0��<�HS<�������(���   �   la���g�艞�Os;j:��[��.�+��=<���F���I�/�E�T�:�(�)�#~�#i���ȾF��-a��W�n½h�V����@|{�_�;pא;�7i�@蔼�s�ѭ��P��������k�:���T���h�4t���u��m���[���A�0L"�z���gv���Eg�@�ۼ���4ׄ<���<���<���<��<<�S�|^E��ý�   �   ��D�*��������(���n�9�6�	P�2�c�1yp���t���o���b���N�%P5���G���������l&G�~���m���!�h�v�������M; ^�9P��}��,/!��q�ꔣ�ypνHs��@5����T���.���	����.3��h ��ҕ&�l焼�=�;���<�=�%=^=�!�<�<�ڴ�WՄ��?���   �   5�j��w�����\��N�4�3�U�,�r������=������` ������6r���T��4��p��Z�uZ���5r�|�"���˽�%e���׼��� �9 ��:@���'-�h���"c���D���z�l��9��՞������ㄫ�`蔽?m�T�%��� ��8�|<��<(a.=��J=�-N=�R4=���<�;�.�`��@Z��   �   a=��䰿�;��&�.L��
q�Hو�j����՝�锠�q���j��X����p�2L���&��U�#�þ�1��S,?��7��E���L9� �t��>:��q�:@?�:��:���(!��T�ͼ^��ȝ �Dr4��>��V>�K1�Vs�0��@���`� �"C<��<d =��L=x%k=�w=*�k=`�B=Tt�< &�9��'�vSƽX�-��   �   ���PҾ<N�d75��^��5���ޔ�$������@�����������#Ӕ�sN���"_��T6�
�k׾
B��J�U��
�(��� 18�(ꧼ@Mû���:�U; ��:@Q��pƷ�x'!��^������ΐ�`�� �<� )�� �8;H�N<���<|�=|�;=�c=I��=䞊=�ӊ=x=��K=�_�< �a�@7F��Y߽>�@��   �   [����ݾ���>�2Cj�6��u������#c��\����]���������N���Ak��w@��E�R.�.뤾��c��z� ط�D:N��LƼ@��  :�d�;�
�;��D; �g:�啺��+�@�T� 26�����; ��;xtS<8��<��<�+=ԌE=B�j==�}�=���=껓=$ �=6P=dZ�<��û0Z�j�ｃ�L��   �   �W���⾿��XHB��Jn�4]���(��X򭿛g�������g��&���T��a���mo���C���[��D?��1�h��������U���мP� �G9���;�̪;��; GC;���: �u:��:@;�;�< �P<썚<H��<�=�u2=�W=dwz=��=��=b�=��=��=ڐQ=lN�<PUỺa�$���#Q��   �   :Z����ݾ#�(�>�+Bj����ˆ�����_b�������\�����O���vM���@k�w@�E�4-�Tꤾ��c��y��ַ��7N�4IƼ����o :@o�;��;��D;�0h:�ƕ�`�+��|T��(6�@����;���;xuS<���<�<�+=��E=j�j= ��=�}�=���=��=f �=�6P=�\�<p�û�-Z����X�L��   �   ����HҾ�L��55��^��4��kݔ�þ������Ĝ������U����є�JM��� _�:S6����h׾k@��܂U�1�
�g����,8��⧼@4û@S�: EU; �:�
������H !�(^��논���͐�X����<��%��`�8;P�N<��<��=��;=d�c=q��="��=DԊ=t=�K=d�<@~a��2F��V߽�@��   �   D;�����B9��&�^+L�bq��׈�����ӝ�ڒ��i���h��������p�P/L�V�&��S�3�þ�/���(?��2��b���$3�ثt���9����:���:��:������T�ͼ(��� ��p4���>��U>�DJ1��r�D�⼀����� �@#C<8�<[d =�L= &k=~w=��k=p�B=\z�< \�98�'�Oƽ>�-��   �   +�j�wt��Z�㾧���4�i�U���r�M�R;��D�������G�����q�&�T��4��m��V��V��,0r�r�"��˽re���׼8�� ��9@M�:�?�`-�4����_���D�4�z�L��I�����S𼽩������!蔽�>m��%�󯼀����|<4��<�a.=��J=�/N=8U4=��<�ɔ;'����V��   �   /�D���������"���j��6�iP�-�c��sp���t�R�o���b��N��K5�p��P���B�������� G���>g���!���v��ὺ 0N; �9����t��@+!�D�q�N���oνr���4�*������ ����	�Q���2��; ��b�&��愼�B�;�ú<U�=Ԡ%=-!=�)�<��<�ɴ�}τ��7���   �   �[�Y�g�5���om;N3��6����+��8<�=�F���I���E�=�:�y�)��y��a����Ⱦ7A���%a��Q�#e½��V�����@�z�`��;��;��h��ޔ��o�ԫ���������f����:��T�T�h��t�}�u��m�d�[���A�L"�K���3v���Eg��ۼ����ل<܌�<���<� �<��<<��R��RE��ý�   �   ���-5���y��o��,wɾ�H�[l���y���Z �����������#龜�¾n+���;k�D�'�u�ܽWȀ�t\� 9˻� �;�<@�p;�((�����u�O��~���4�B�`�}���u������$į��籾n������𩐾Qw�e�H�^p��yؽiF���w��RԻ��<<�r�<H��<(`S<p�����H����   �   ���)����<���v��������� JоT�%��M��>��
�߾��ɾΠ��L��P�b���'��c�*\��fW�@.��hv
<�Xu<��H< k:����"J�L��>��z�<�t�v���������MоX侅��R��ٌ�߾�ɾ����qO���b�f�'�Lk�)b���`�`f�� b
< Ku<�H< P:�����J��   �   ��u��	����_ 4��`�秅��q��N���r����㱾���š��d����Jw���H��k��qؽ�?���m�Ի��<<�{�<�<�eS<н�����& ����05�<�y��q���yɾ�K�Yn������X] �{��P��3��(�j�¾�.��9Ak���'�2�ܽ�̀�,l� g˻� �; < �p;p&(�����   �   &l����������������:�(�T�Ѡh��t�>�u���m�B�[���A��F"����Dn��,8g�4�ۼ@�X�< ��< ��<��<��<<�R�tTE�}ý�]���g�熞��o;66�������+�$;<�ҢF�>�I���E���:��)�K|�f��u�ȾD��**a�MU��j½ �V�(���={� �;��;��h��۔��   �   Tp��0'!�J�q�-����iν�k���0���d����}�;|	�V���*�����Ĉ&� ф�0��;�Ѻ<ص=�%=0$=�-�<��<�ʴ�iЄ��9����D���������%��cl���6�sP�~�c�tvp�L�t��o���b�t�N�\N5�������>���# ��_$G�����k���!�`�v� H���N; ��9����   �   �-������[���D�v�z�����������s鼽y���F}������&1m���%��ܯ�@����|<��<�g.=&�J=�2N=�W4=L��<�ϔ;D'����HW�j�j�nu����㾙��F�4���U���r�Y�z<�����7�������Z r�i�T��4��o�qY�MY���3r�@�"���˽�"e�0�׼h�� ��9 .�:�=��   �   �:�X����H�ͼ���R� ��h4��>�8L>�6@1�vh���L���  �PCC<x�<~j =0�L=P*k=�!w=B�k=��B=l}�< ї9�'�EOƽ��-��;�������9�8&�J,L��q�<؈�V����ԝ�ߓ��~���-i��������p�1L��&�1U�U�þo1���+?�~6��V����7���t��:� ��:���:�   �   ��:�� ����!��^��ㅼ$
��(�p��0�<�`�@9;�N<���<��=t�;=��c=<��=���=~Պ=�=ܽK=(g�<�ja��1F�_V߽��@������Ҿ#M�65���^��4���ݔ�U���C�������M���(����Ҕ�N��["_��T6����j׾�A���U���
�쐨�x08��觼pDû�(�: ;U;�   �   0�;`�D;�Gh: ����o+��aT� 6� ���@A;���;�S<���<P
�<�.=E=��j=(��=�~�=���=���=,!�=\8P=�_�<��û�+Z������L��Y��w�ݾ��>�4Bj��������&���b������3]��I��ԣ���M���Ak��w@��E��.�e뤾A�c��z��ط�;N��MƼ����! :i�;�   �   ����^���W�(�м�o��Hf{�^�@ꔺ�K�; �|<��<p		=�	/=�nT=��w=짋=��=���="#�=@��=�Δ=��y=d�-=�<����bo���7Y��a����վ6.
�j�*��/J�KDf��n|��P�������P��|���f���J�N�+�K�B�۾�j��I#s�� ,�:��,¢�B�b���'�zr	�X�������   �   L���dj����āܼ�I��p�����B��ß���9;�B6<$9�<���<fK=x�D=��i={��=Pt�=KX�=tơ=��=�=d�w=F�-=LR�<@���:��֦��U�W���Ҿ���"�'���F�pTb�S"x�A��%q�����$x�9�b��2G��(�ā	���׾�"�� n��7(�����읽B�Z��F!�X��\�0���   �   $`�N�����l� �����׼���%��`�� ���Y�;�t�<��<6�=X�?=|qf=�߃=\��=���=�_�=��=�:r=x-=䍍<�㍼���������I�i,���Ǿ�� �e�ƚ<���V���k�l�x�6m}�`�x�jxk���V�~�<�������˾����R_�I���ֽ@ڏ���C�jL��2��ۼ@"��   �   `��R�����t"��(�#(��"��f�l���ͼ�7����׻0"�;���< c�<��'=��R=x�u=�V�=]L�='̄=��g=Ȧ*=��< ?T��Hc�'��Z�6��R��J�f�� ��.�,��E�{X�lGd��`h��d���W���D��,�	��R��M޸�;Ɗ�HKH��4W����s��9 � �⼘9��ԫ���*ϼ�   �   \�����n�:�@�W���p�H����N���"��ds����q�~P�Z#���ټ�@�`�v;�R�<��=b 7=��Z=~~n=tTn=��V=+�$=8��<0��z<�M�½���j��~��,о[� �����_.��I?��J��M���I��>��c-���������/Ͼ� ��&�o��+�l���㖽
p;���漸������\�����   �   �w	���;�L!q������������ҽ#4ݽNJ߽3ؽm�ǽk)��4��f�M��R��8�)���<���<C�=�l;=�H=�>=��=�٭<��E�4��8�����%G�<�������k�۾���4��3R#��u,��d/��+��!"�E�]� �R�׾�ﭾ ���VE���	� ���]���������H��X���i����   �   "H$�l�n������Aɽ/@�������X�&��,���*�0"�2��X��za̽*����B�����  d��q�<x��<��=��=Sm=�V�<��f:�2ۼ�E��^۽4�#��7a��W���I���%׾I:���h����U�������f�3Ѿ	���]u��8LT�7��Pν��}�X��0�g��_g� X���e���A��nǼ�   �   wO�vA���;ԽxC���&�v(C�D�[��.n�V|x�rfy�1�p��\^��nD��$�RO��i��ڝw���P����2<�z�<� �<<��<�e�<�>J;@	���XF�T+���A�A�3���i��p��w ��k�¾�վ's�ܑ㾅޾�mо��������x��$�S�ܮ��ڽs������� U�@ �:xM<�-�;��e:��=�؄��   �   !4���ʽқ�p�4�g�^�3w��v��ǐ��"���eg��酧�~c��k���£o��"C�p��H�սda���5��7� ��;�"�<p[�<��e<��M;�le�H��1��ʽ����4���^��t���
������ԣ��d�������`�������o��C�0���սO]��h/�s7�P��;�'�<^�<��e< �M;Xve�d���   �   /��D���3��i�\s��y#��ǻ¾�վ�v྘��޾9qо��������Hz����S����e�ڽ��������U����:�F<�'�; �e:��=��~�JrO�>��E7Խx@��&�#$C�b�[�:)n��vx��`y��|p�W^��iD���$��K�?d����w�^� ���x�2<���<�<���<�d�<`$J;����]F��   �   �۽!�#�h;a��Y���L��H)׾�=���j����R����˶�%j�j6ѾI���-w��OT�f���ν��}�$��@�g��~g� 鼹�e���A��jǼ�D$�:�n�����<ɽ\:�_������&��	,�&�*��+"��-�(Q���Z̽X$��F�B�H��� wb�0{�<���<?�=�=�m=�T�< kf:�:ۼ�H���   �   I���(G�:�������_�۾n����-T#��w,��f/���+��#"��F��� ��׾?�Y��YE�2�	�Q���]������������8����i���ju	��;�q��	��a��������ҽ�-ݽZC߽,ؽ��ǽ�"���-����M�x@��P�)��<���<�=�o;=��H=��>=h�=�֭<��E��������   �   v��<�j������о�� �h��^a.��K?�oJ�ޞM�b�I���>�e-��������[1Ͼ�����o�$+�T��>喽Br;���<��LÄ�������x��������:�*�W��p�^���tJ�����.n���q�P�f#�dvټ(�?� Ew;�^�<��=,$7=��Z=|�n=�Un=�V=t�$=���<����<���½�   �   ��6��S�� ������J����,�.	E�X�
Id��bh��d��W���D�΃,�Ƶ�q��"߸��Ɗ�"LH���"X�� �s��: �Љ��:��X���`*ϼ��Ｎ��>���p"�`(��(��"��_�����̼)���׻�V�;���<m�<��'=P�R= �u=�W�=�L�=h̄=X�g=��*=��<�KT��Mc�x���   �   zI��-��UǾ� �p��<���V���k���x�Un}�e�x�Jyk�s�V��<�S��J�#�˾Y���/S_����/ֽvڏ�"�C��L�D3�ۼ�!��^��K������ ������׼������P�� ����;�}�<h��<��=��?=$tf=���=%��=!��=`�=��=@:r=4
-=Љ�<�鍼���������   �   'U�I����Ҿ>��۰'��F�5Ub�#x����qq����w$x�x�b��2G��(�	���׾�"���n��7(����r읽��Z�|F!��<\�t�� ����h������~ܼpF��������B�����@:;�L6<�=�<���<dM="�D=:�i=��=�t�=�X�=�ơ=��=��=x�w=��-=tN�<�$���<�����   �   �8Y�7b��G�վ�.
�Ƨ*�0J��Df��n|��P�������P����|�c�f�b�J���+�����۾@j��X"s��,����,�����b���'��q	��������H����\���V���мDn��d{� \� ޔ��M�;��|<��<_		=t	/=FnT=|�w=���=ԗ�=`��=�"�=ԅ�=Δ=܆y=�-=
<P�������C���   �   �U�����Ҿ����'���F�6Tb��!x����p�����]#x�tb��1G�N�(��	���׾�!���n��6(����락h�Z�`D!� �dX�ı𼠙��pe�����|ܼ�C��T����B�����`:;�N6<�>�<h��<�M=P�D=T�i=��=�t�=�X�=�ơ=��=�=�w=-= Q�<!��Q;��$���   �   :I�*,��hǾ�� ���9�<���V��k�p�x�l}�2�x�3wk���V�V�<�ִ���˾�����P_����ֽ�׏���C��H��+��ۼ��4X�dE�����P� ���񼠴׼@��������������;�~�<X��<7�=ظ?=htf=���=P��=X��=e`�=�=l;r=�-=���< ㍼N��������   �   r�6��Q��v�J��H��G�,��E�7X�Fd�s_h��d��W��D�j�,������Zܸ��Ċ��HH����S����s��4 ��~⼐0��D���� ϼ0��,�����l"��(��(�"��]�j��<�̼'����׻`[�;���<�m�<L�'=��R=��u=�W�=jM�=̈́=��g="�*=��<p8T��Fc�ک��   �   ���P�j��}���оd� ����7^.�H?��J�.�M�ÞI�>�>��a-�������F-Ͼ������o��*�Ҵ�����i;� �漼 ���������H��4�������:���W��p������H�����8m����q��P��#�uټ�?�`Lw;�_�<�=�$7=8�Z=~�n=�Vn= �V=Y�$=ܐ�<�t��w<�/�½�   �   9���#G�ε������4�۾i�����uP#��s,��b/��+��"�C��� �9�׾�쭾���SSE���	�/���]�����$|��ؾ�X����i��㹼6o	�2�;�~q�
��&������L�ҽD,ݽSB߽E+ؽ��ǽf"���-�� �M�d?��8�)�(�<���<��=�p;=L�H=�>=��=�߭< RE�֠�����   �   r۽��#��4a��U��bG��;#׾7��5g����R������>c�H0Ѿ ����r���GT����rνR�}�Fz���g�`�f� �� �d�x�A��]Ǽp>$�N�n�C���h:ɽ 8�n��Ԭ�p�&�	,�ĕ*�V+"��-��P��}Z̽$����B�H����Ob��|�<���<��=>�=�p=(^�<�h:P(ۼ�B���   �   5'���>��3�̃i�zn�����U�¾�վ{o��㾯޾'jоl�ƌ��Lu��H�S�Ȫ�H�ڽ�|��J��0�T����: h<�c�;�hg:`�=�Hr�6lO�(;���4ԽE?�ސ&�@#C���[��(n�Uvx��`y��|p�NW^��iD���$��K�d��0�w��� ������2<��<��<0��< n�<��J;,����QF��   �   �,��ƃʽ�� �4���^�r��������������`��E��-]������a�o��C������ս1W��6%��P7� �;$5�< k�<�f<��M;@Te�v��?.��.�ʽ���4���^�3t��5
��]��������c������l`��������o��C�����ս
]���.�0o7����;�+�<�c�<�f< �M;�Ue�t���   �   ZjO�K9���1Խ(=��&��C�p�[��#n�qx��Zy��vp��Q^��dD��$��G��\���w��� �pc�p�2<���<��<\��<4r�<`�J;l���~SF��(��b@�>�3���i�ap��# ��(�¾�վ s����r޾�mо�����x���S�Ů���ڽ"��������T��9�:�W<PK�;��f:@�=��q��   �   l=$���n����7ɽ�3���s����&��,�M�*��&"�?)�ZH���R̽)����B��y���)`�Ԋ�<��<S�=��=|s=ta�< ;h:4)ۼ�C��R۽F�#��6a�(W��fI���%׾:���h����L�������f�3Ѿ���Vu��$LT���ν:�}�V��@�g� =g� Ǻ� �d�X�A�,^Ǽ�   �   �n	���;�|q�����������$�ҽR&ݽ�;߽W$ؽ˕ǽq���&����M�l)����)�p<���<��=Vu;= I=؝>=��=t�<@JE�j��v��"��$%G�消�;���.�۾���!��(R#��u,��d/��+��!"�E�[� �M�׾~ﭾ����VE���	�����]�,���@���0��8��p�i��幼�   �   ����p����:�T�W�Z�p�����6E��Z��bh��B{q�P�O�
#��`ټh�?�`�w;dn�<��=.*7=��Z=<�n= Zn=��V=-�$=8��<xr�x<��½}����j�y~���оE� �����_.��I?��J��M���I� �>��c-���������/Ͼ� ���o��+�6��㖽,o;�������4����������   �   ��������j"��	(��(��"��W������̼��@S׻���; ��<Hz�<��'=��R=��u=�Y�=�N�=+΄=�g=��*=�!�<�5T��Fc�4���6�OR�� �D����$�,��E�wX�lGd��`h��d���W���D��,�	��P��J޸�6Ɗ�6KH����V��
�s��8 �@�⼼5��\����#ϼ�   �   �Y��E�����`� �����׼,������v�@A����;D��<���<��=�?= xf=t�=ć�=���=oa�=��==r=d-=(��<����䥁�]���BI�K,���Ǿ� �]���<���V���k�l�x�6m}�b�x�lxk���V�~�<�������˾����R_�<���ֽ
ڏ�$�C�|K�00�xۼ���   �   0���xf��(���{ܼ�B�������B����� ::;�V6<$C�<(��<�O=��D=|�i=$��=�u�=zY�=pǡ=��=��=|�w=*�-=�S�<���q:������U�K���Ҿ����'���F�nTb�S"x�B��%q�����$x�9�b��2G�	�(�Á	���׾�"��n��7(���罷읽��Z�rF!���([����   �   
@���ﯽ{P��sѓ�Ѐy��C�v	�pW��P���<D�<=PC<=� f={O�=���=�z�=3L�=,C�=p>�=`�=�ڊ=huZ=��=@�;Й��I����	��9O�������@T龈�
�����.�_�8��l<�x�8�O�.��;�����U�O����q��̈j��v1��x���ѽ����c��hl���ӟ�a�������   �   �!��T������K����~{�$�G�P������� ��;L��<C�=�B0=��Z=�#�=��=Hy�=��=.u�=^�=�?�=���=�(Y=E�=� �;`�������,=���K�V���;���?����",�:�+���5��9�U�5�6�+��[��(	����h:���j��Ģe�l-��3�J2̽�!���������������e���]���   �   [V��,��kt��a{��8L���wV�4Q%����s��a
�`�)<D@�<�=pI8=��`=��=�[�=��=v��=�3�=3��=K�=��T=�Z= u�;D��k�������m�@����Į�xپ҇�����"��F,��{/�',���"���\��	!۾��������wjW�y�!��[�&����F��a��������*ӡ��   �   U����K��^q���������@r��oL�:�"�h�뼈ٍ� �����;l��<���<O+=��T=&�w=�C�=&��={w�=꿍=:~=fUL=��=P��;L�ȼ0�����V�0��;u�3���FǾ�L�V��u� ��^| �X�"��L��X�r1Ǿ�͡���}�h2A����sս/^��mۃ��Zl��j�J!x������!���   �   �L�������s���욽?=���ȏ��ꄽ��m���K��#������=p���<���<v=�<=Χ`=lsy=`[�=��=Pi=�B>=�7�<С<����
&i�b
Ͻ���ϼY���������Ҿo��®��#������
�����.��Ͼ��������[���$���d*�������oM�¿6���7��#I��-c��g��   �   ~�~��Џ��z��������wg�������G���㡽�-��8Tz���F�^�D����m���W<P��<U�=�>B=� W=��Z=L=�')=LL�< R<X?���gI��g��@���;���t�ʃ���ɳ���̾b�ྎ����53�JIݾgBȾ5�����ʂi���3������h��C8�r���� & �� ��6���Z��   �   J+m��ꏽ�^��W&��(\ӽ��㽆c�Fw��G����ALӽ����]p��vx]�N2�H'q���T;Tv�<I�<�=�r+=��%=��=�I�<0��;t���@/�G"���%����M��|��&��#I���鸾�y¾��ľ￾R󳾦"���1��
?h���7�Ď
��ƽ�����E*�8LҼ�&����o�v��<�Ǽ"��r�:��   �   Xh�s��wV��l���8�E�E> �E�(��,�*)����Sq�W����ȽE�����F� �м�����	*<P�<���<���<tP�<���<@p	;0��������=Ľ^h���(�!�M���p�,�������㙾�
���S��.��8�z��hV���.�}4��!Ľ�8�����.���ջ ��� �J80ϖ� �[�XqѼ�$��   �   @(r�x����ݽ��	���$� �=���R�qzb���j��Nj�|a�u�O�"7����N��q�H�p��v�8WQ� =;�K=<�Bx<�[<0Q�;`���|��<��%r��u����ݽn�	��$���=��R�1vb��j�ZJj�a�H�O�U7�������볽n�p�jp�HBQ���;Z=<pNx<8[<�_�;����d|��:��   �   ����@Ľaj�z�(�r�M���p�k���� ���晾f���U�����h�z�mlV���.�7��%Ľ�;�����8��P:ջ 9�� �?8�ᖻH�[�hsѼ�$�h���T���⽎6�KB�; ���(�,�W)�ɽ��m��P���ȽB��F��м ʴ��*<�<���<Ї�<$T�<���<@v	;�������   �   �$��T)�J���M�Ӥ|��(���K���츾d|¾��ľ�������$��x3��ABh���7��
�4ƽF���lJ*��SҼ`-����o�`{����Ǽ���L�:�+m��鏽4]���#���Xӽ��㽌^ｱq��C�����"Fӽ䤷��j���n]��)��
q�@U;8��<Q�<��=fu+=��%=�=�J�<`��;����C/��   �   �j��/����;��t����˳�8�̾��^�����5뾾Kݾ�DȾ�6������N�i���3��������j���F8�������( �T#��6��Z� �~��Џ��y������	��gd��報��C��^ߡ�)���Jz�\�F���Ą��` ���W<	�<M�=BB=pW=��Z=HL=�()=L�<N<�C���kI��   �   UϽ���l�Y��������
Ҿ������$�J���
�����0�Ͼ-���Ң���[�%�$� ��,,��#����rM�z�6�@�7�*&I�0c��i�?M�� ���'s���뚽�;���Ə�脽@�m���K���#� ������o���< �<�z=��<=�`=�uy=R\�=D�=�Pi=�B>=�6�<��<����$*i��   �   ҫ�B�0�:>u��4���HǾ�N�l����D��z} �	Y����Z�2Ǿ�Ρ���}�`3A����0uսE_��p܃�]l�j�`#x�� ���"��捚�/L��Bq��������fr��kL�ܖ"����`ύ�Z��0��;���<B��<�R+=ԭT=Ĳw=�D�=���=x�=?��=L:~=$UL=��=0��;�ȼC����   �   �����@�ą��Ů��yپ�������"��G,�`|/��',���"�u�ü��!۾���⢌��jW���!�6\�����nG�����q�������ӡ��V��M,��bt��{���K��vV��N%���⼠ss��,
��*<�F�<�=(L8=��`=��=�\�=���=���=4�=L��=+�=L�T=\Y=�e�;Ȭ�[����   �   9>��K�!	���<���@很���,�¶+�.�5�9���5�x�+��[��(	����h:���j����e�E-�e3�2̽�!�����������"f���]���!��X�����������}{���G���� ��� ��Ф�;���<��=dD0=��Z=K$�=�=�y�=��=Du�=V�=�?�=���=�'Y=��=��;T���L����   �   ��	��:O���������T���
����)�.�t�8��l<�g�8�-�.�};�}��uU�����rq���j��u1��w��ѽ���c���k��8ӟ����o���?���ﯽ7P��,ѓ�<�y�^�C��	��V������<|�<=,C<=� f=YO�=���=�z�=�K�=�B�=#>�=�=rڊ=LtZ=k�=��;қ��J���   �   ^=��K�j���;���?����+���+�Z�5�:9�ڦ5���+�[�(	����x9���i��\�e�?~-��2��0̽l ����������p����d���\��� �������땓��{{�N�G��������������;Լ�<<�=�D0=�Z=j$�=2�=�y�=��=eu�=w�=�?�=���=l(Y=��= ��;��������   �   H�����@���*Į�vwپl��t�	�"�F,��z/�;&,��"������۾<���j����hW���!��X��뻽����D��������!���/ѡ�@T���)��r���x���I���rV�L%�l��8ls��
�*<hH�<��=�L8=Z�`=��=�\�=أ�=��=V4�=���=��=��T==[=�z�;���휒��   �   P��O�0�s:u�(2���EǾ�K�������D{ ��V����-��V쾍/Ǿ̡���}�0A����pսL[���؃�"Vl�2j�zx�2������e����H��
n��"��4����r�hL���"����dˍ��M�����;���<���<ZS+=T�T=@�w=�D�=F��=rx�=���=�;~=�VL=?�=0��; �ȼ㹄��   �   �Ͻf���Y����#���Ҿk�ﾞ��\"����P�
�G��E,�|Ͼ��ޟ���[�*�$�t��&��S����iM��6���7��I��'c�*a�I�����[o��[蚽�8���Ï��儽��m���K�|�#�t��� �o���<t�<&{=N�<=x�`=�vy=�\�=��=fRi=�D>=(=�<`�<�屮 "i��   �   �d��]����;��t�����ǳ�h�̾ݑ����>��K0�oFݾ�?Ⱦ�2��Ύ���~i�O�3�Q��_���d��<8�������� �&��6��yZ���~�̏��u��:���J��ra��h����A���ݡ��'���Hz�܍F������������W<L
�<��=�BB=\W=�Z= L=+)= S�<Xa<x6���bI��   �   ����!�_���M���|��$���F��S績�v¾��ľ(쿾|����/���:h��7���
�Oƽޑ���=*��=Ҽ@����o��h�� �ǼN����:��!m�M叽 Y�� ��dUӽ���\ｪo�������%Eӽ'���cj���m]�")� q��U;���<�R�<��=�v+=��%=��=4R�<���;�	���:/��   �   ��:9Ľ�e���(���M�z�p�ℇ���Iᙾ���P����*�z�&dV���.��0��ĽT3��*��d��p�Ի G�� e8P�����[� aѼ�$� h����P��\���4��@��9 ���(�D,��)�T��lm��O����Ƚ���F�Ԑм0Ŵ��*<��<l��<h��<Y�<ܴ�< �	;x���H���   �   �r�Hq��0�ݽb�	�s�$��=���R��qb�2�j�ZEj�a�s�O��7�|��2��,峽<xp��f�!Q���;�t=<�gx<�/[<Е�;Pđ��k���
��r��q��ևݽ��	�l�$���=��R�[ub�k�j��Ij��a���O� 7�x��P��j볽�p��o��?Q���;�^=<�Tx<`[<`y�;0ܑ�Hp��,��   �   h����	O��Z��`3��>�F7 ���(��,��)�v���i��H����Ƚ�镽F�H~м����`:*<H$�<4��<Г�<T`�<���<��	;$������f��[:Ľ�f�`�(�ݝM���p�����.���㙾�
��XS����	�z��hV���.�_4��!ĽM8��z��p-��pջ 㪹 �R8������[��fѼ��$��   �   |#m��叽�X�����*Sӽ����Wｸj��
�����>ӽ蝷�ed���b]��8�p� �U;��<*^�<و=�z+=O�%=��=0W�< ��;���r:/�=�� #罝��dM��|�*&���H���鸾jy¾��ľ�?󳾗"���1���>h���7���
��ƽA���8E*�tJҼD$���o�Xq����Ǽ���x�:��   �   6�~��̏��u�������4_��j���>��x١�##���>z��F�&� q���r�h�W<�<u�=�GB=hW=��Z=L=�-)=(W�<8g<�4���bI��e������;�Ғt�c���Mɳ�g�̾1��i����#3�=Iݾ]BȾ	5��������i���3�������jh��fB8���x���$ �*�&6��|Z��   �   HJ��煕��o��.蚽�7��^��ㄽ@�m�v�K���#����,戼 Qo�� <�<̀=L�<=ԯ`=Lzy=^^�=>
�=�Ti=�F>=�@�<��<\ "i��Ͻ��	�Y����I����ҾA�ﾰ���#�����
�����.��Ͼ���������[���$����1*��R���6oM�Ⱦ6�@�7��!I�+c�Bd��   �   �����I���n��C������0r��eL�B�"�L�������$��P��;ଙ<���<�W+=��T= �w=~F�=���=�y�=���=�=~=�XL=��=��;d�ȼ˹����齻�0�;;u��2���FǾ�L�G��k���Z| ��W�!��K��X�n1Ǿ�͡���}�[2A� ���sս�]��&ۃ�JZl��j��x�����o ���   �   >U���*���r��2y���I��rV��J%�x��@bs���	��*<O�<�=�O8=d�`=/�=>^�=���=��=>5�=z �=o�=�T=�\=���;��漄�������@���xĮ��wپƇ�����"��F,��{/�',���"���[��!۾��������pjW�n�!��[�ꠚ��F����R��h���Uҡ��   �   I!������#���9���|{�<�G��� ���`��@��;���<��=hF0=��Z=8%�=��=gz�=��=v�=�=U@�=���=�)Y=G�=0�;����?����<���K�C���;���?����,�6�+���5��9�T�5�5�+��[��(	����f:���j����e�h-�~3�72̽�!����������R����e��Y]���   �   E�3�#0�	�%�8(��  ���Ͻ�'����U�4J� n�B<|��<��1= pd=� �=�L�=��=6_�=��=�T�=e͡=o�=�Lv=d5=�о< �f���ܲ���\��B6�k�q�����0��1ѾH��=`��W���^��,��xҾ�b�������>���XQ�P)��q��l��㽮t�Ԡ���V
��O���&��.0��   �   �R0�/%-��'#��4��g��ܖν8��R0X�9��@8�ح%<�C�<�)=��\=�N�=���=X�=%��=��=�1�=��=���=�\s=�"3=\K�<��d�����n�������13���m�Us��A��:�;?��w�m��������fξ�޴�͂��zB}��L��;%�J ��`�w�ݽ|��(��:%�5���M#���,��   �   ��&��$����K��jL��v~˽+ ���`����`�\����;$Ь<��=��D=P'p=��=m��=pL�=!�=6��=���=,r�=�>j= ,=8ĳ< �g�~[���n���+��b��!�����þ��־�a�
�� �>:־P�¾����z����n��@��5������ڽ��̽ŬнB��O���u4�9G�Ǽ"��   �   �i����^I�l��ô�HaȽ�#��:r�`�#��[�������$4<�t�<4=�I=��o=NІ=��=|r�=E2�=K��=�-�=�Z=a�=P_�<����B	��I��n�߽Ӽ���Q���J���ֲ�ۚľ��Ͼ|rӾ5Ͼ�þ�����͚��ł�,UV���+����J�޽�
��X�����kƽk�޽,3��>�	�B~��   �   ����N�����L��k��Ƚ�-�� ����EO����/�� ����(<X��<�R=�1==N�_=Jey=��=M��='��=��h=DyA=�*
=T�< ������M����ͽLA���<�@�j��A������)𭾈h���"���ε��䪾@���M���Zib�k*8��!����[���;|���F�������H��M+��HԽfN��� ��   �   ��轝�𽏰�d�߽��ͽ�?��)����&��T�Y�:� ���ʼH'�p��;\C�<��<ݎ#=V^C=��W=�^=PjX=|GC=�>=:G�<(�'<��������y�9޼�4���,'��:M�>�q�¯��a�<R��r��������ݏ����k9`���:� ���齚C���:��hqe�N�R��1Z��v��	���%���"ý��ؽ�   �   �ŽMԽL޽¢��H�Muݽ�hԽ�>ǽ���T����0��H�T��Y� /��`���@�<x��<���<P�=��'=&%=?=j��<t��<@i�:dU��.�V(w�Bǰ�l.�w��1�),M�jie���w��ۀ��M��S�y�,4h�<O�?h1��~���I8��<�{�>�7�N������vT���#�AM�Ђ~�yᘽ۰��   �   3Ħ�����9ҽ�
�7&�&��d	���D�������(ͽ�Y������xES��[���� 4�X><���<dE�<h��<�z�<�sj<@mm;H�"���Ӽ*53����)���Uؽh���i�LV,���<�҄H���M��L�J�B�.�2��3�?���5ҽ����e^��{�<���@a�X6� ~]�Hz��D���A-��lc������   �   v܏��J��н�r��'���c*�[e����PB�*:�FH���޽)ȳ�q����7��Dּ��1� F9`�;(\<�Ϥ; t���E�4ʼ�����^�&ݏ��J��Rн3q&���$(��b����a?�@7�zE�U�޽�ó�W����7�h8ּ��1� �90A�;�l<��;���`�D��ʼ����^��   �   ������`Wؽ����k��X,�J�<�ۇH��M�L���B�Q�2��6����:ҽ���4l^�&����� a��!6���]�(��� ���E-��pc�B����Ŧ�t���9ҽ
�p$�~������@��h��%��$ͽ�T�����`=S�TT����� �2�H><$��<M�<���<���<�j<`�m;��"���Ӽ�33��   �   n)w��Ȱ��0���1��.M�{le���w�Z݀��O����y�7h�!?O��j1�����佑;����{�88�������� Y�(�#��EM���~��㘽/ݰ�cŽZNԽ�޽����G⽈sݽXfԽ�;ǽ��r���-��x�T�fR�t!�� z����<���<���<��=Χ'=+"%=�A=���<���<@��:0S�� ��   �   ��y�༽����.'�:=M��q�`���'���T��J���O���Rߏ����� <`�-�:������<F��:=���ue���R�H6Z���v�!��9(��E%ý��ؽ���>�𽜱��d��߽��ͽ$>���3$��x�Y�~ ���ʼ��&����;0M�<���<��#=�aC=��W=��^=�lX=�IC=P@=0J�< �'<�������   �   �N����ͽ�B���<���j��B��E�����Lj��@$��Jе�Q檾����t���Kkb�,8��"����]·�~���H�������J���-��yJԽ�P�� ����oO�;���M����㽚Ƚ�,������"BO�����&��`�X�(<���<�V=5==H`=�gy=��=K��=��=<�h=dzA=�+
=��<@�������   �   aK����߽K����Q���LK��ز�\�ľ\�Ͼ�sӾ�Ͼ;þ� ���Κ��Ƃ�\VV���+�u����޽V���Y��"���lƽF�޽,5��@�	�?��j�n���I������ aȽ#��8r���#��U��0暻24<B{�<7=��I=D�o=Yц=� �=>s�=�2�=ѫ�=F.�=xZ=��=�^�<���8	��   �   � ��u��K+���b��"�����2þ�־c�"����;־�¾1���점��n�@�W6�M�����ڽ_�̽��нa�ὑ���(5��G���"���&���$�������L��j~˽����ܵ`�L��З\�0��;TԬ<��=��D=
)p=ɇ�=��=�L�=!�=���=!��=Or�=�>j=� ,=�³< �g��]��   �   'p��^����23���m� t�������;���!����
��\�⾨ξ�޴�ₙ��B}��L��;%�F ��`콤�ݽ��ὒ��}%����N#���,��R0�p%-��'#��4��g����ν:8���/X�7��(4��%<
F�<�)=��\= O�=N�=��=Z��=*��=�1�=��=���=8\s=4"3=0I�<��d�����   �   ���]���6� �q�����a0��f1Ѿ}��[`��\���^�����:Ҿ?b��l����>��LXQ��)�vq��k򽈖�8t�}���cV
��O�s�&��.0�*�3��"0��%�(��  ���Ͻc'��2�U�tI� l��B<���<��1=pd=� �=dL�=|�=_�=��=vT�=͡=�n�=�Kv=c5=tξ<��f�ι��   �   �n��΄���13��m�Cs������;��� �ܛ�����F�⾦ξ�ݴ����+A}���L��:%�h�0_��ݽ7�����$����M#���,��Q0�t$-��&#��3�f��h�ν7���-X�@4���/���%<TG�<��)=�\=JO�=j�=��=l��=H��=
2�=��=й�=�\s=�"3=,K�<��d����   �   @��|��g+�b�b�s!�����Sþ��־�`�����9־�¾~���n����n��@�v4�����оڽs�̽ĪнF��D���d3�F���"���&���$�R������I���{˽����j�`�����\����;�֬<��=��D=�)p=��=H��=$M�=�!�=ɜ�=h��=�r�=�?j=,=tƳ<@�g� Z��   �   -H��{�߽���B�Q���I��|ղ���ľc�Ͼ�pӾ��ξ_þ����~̚��Ă��RV���+���� �޽���U����|hƽ��޽J0����	��|�h�ӱ��G�����콧]Ƚ5 ��P3r���#��O���Ӛ�94<~�<8=��I=��o=�ц=!�=�s�=<3�=9��=�.�=�Z=��=�c�<0熻`	��   �   K����ͽ�?���<� �j�?@��8�����f��� ���̵��⪾w�������`fb��'8�=����ü���x���C�������E��
(���DԽ�J�� ����VL�Q��*H��Ƹ�tȽ;)��ĝ���=O�>��(!��p჻��(<$��<�W=�5==�`=thy=�=���=~��=x�h=|A=.
=0�<0����{��   �   h�y��ڼ�,��u*'�18M�>�q������IP��k���y����ۏ�8���5`���:�7�����S?��7��pje���R�H+Z�4�v����!���ý�ؽ�~轊��H��_뽠߽�ͽ[:��ٹ���!����Y�
{ �4�ʼ��&�pȆ;8O�<F��<a�#=dbC=J�W=��^=�mX=�JC=,B=lO�<�'<x��J���   �   � w�ð��)����1��(M��ee�Ƌw��ـ��K��0�y�*0h�T8O��d1��{�0z�e3����{���7�&������M�X�#�z9M��z~��ܘ�3ְ�hŽ�GԽ�޽��⽔B�oݽ�bԽb8ǽ��}���z+��*�T��P����pq���<,¯<��<� =��'=E#%=BC=Z��<T��<��:PI��~��   �   �{�������Pؽ����f�S,�
�<��H���M��L�T�B�\�2�30�����/ҽ���V\^�4s�(ﲼ`�`�(�5��b]�l�����N9-�vcc�����ξ��� ���3ҽg�l�*��Q���=��	��I�㽟"ͽ�S���~�� <S�XS�쩂���2� ><���<�N�<���<l��<��j<��m;h�"��Ӽ�-3��   �   �؏��E��!н�k#����$�7_����;��3��A���޽s��������7��&ּ��1� 9v�;��< $�;���D��ʼ���2�^�
׏��D���нl�K$����&�sa�����>��6�E���޽�³������7�7ּ�1� �9�G�;�p<���;�����D��ʼ:��X�^��   �   ��������4ҽ�㽰�p������=:����򽖌㽝ͽ�N���y���2S��J�,��� �0�H4><���<<Y�<��<ȍ�<Țj<�n;�r"�@�ӼR*3��z������Qؽ0���g��T,�,�<���H���M��L���B���2��3���85ҽ���"e^��z����pa��6��y]�Xw�� ���>-��hc�����   �   �Ž�IԽ�޽t��}B�nݽ�`Խ�5ǽ��˃���'����T�~H�<���7���<<ί<���<�=(�'=t'%=EG=(��<���<���:$C���Pw��°�d*꽡�1��*M�Dhe���w�2ۀ��M����y��3h��;O�h1��~���8����{���7����H����S�D�#�b?M�|�~��ߘ��ذ��   �   P�������>`�߽��ͽR9��!���k���Y��t �d�ʼP�&����;�Z�< ��<O�#=�fC=^�W=:_=@qX=TNC=kE=rU�<H�'<Б�x��z�y��ڼ����U+'��9M�(�q�P�����Q��>���]����ݏ����J9`���:����^��gC���:���pe���R�,1Z��v�	���$���!ý��ؽ�   �   ��M�F���I����㽧Ƚ�(�������:O�p��p��ໃ�е(<���<\=:==�`= ly=��=(��=숀=:�h=�~A=q0
=��<����Lz��J����ͽ@���<�I�j�%A��]����ﭾXh��["���ε��䪾0���B���Fib�X*8�z!����3���|��yF��E����H���*��hGԽrM�R� ��   �   (i���mH�B����^Ƚ) ��F2r�,�#��J��л��(F4<Ƅ�<v;=��I=��o=ӆ=t"�=�t�=_4�=R��=�/�=�Z=��=�g�<�چ�*	��G����߽����Q�o󂾼I��hֲ���ľ��ϾerӾ&Ͼ�þv����͚��ł�UV���+����)�޽�
��SX��d���jƽ�޽�2����	��}��   �   ��&�u�$�������J��l|˽�����`������\��̛;�ڬ<��=��D=�+p=��=8��=N�=�"�=���=:��={s�=�Aj=�,=�ɳ<�g��X����:��r+���b��!��e���þ��־�a������9:־J�¾����v����n�}@��5�l�����ڽf�̽��н�����O4�G���"��   �   dR0��$-�P'#�D4��f��ٕν]7���-X��3���-���%<@I�<��)=�\=�O�=�=<�=���=Ȅ�=�2�=&�=h��=�]s=2$3=�M�<��d�j��2n�����|13�L�m�;s��,��,�;3��n�h���������cξ�޴�˂��tB}��L��;%�F ��`�i�ݽf����-%�"���M#���,��   �   �n��5l��?����݂���b�v�;��E�!}׽$�����hR�p�o<p�=�M=�9�=��=u�=��=L��=̉�=��=�=-9�=ܧM=h�=�o<(T��������}׽�E���;�U�b�l܂�͛���j��#m���l��9��5��]�i���I��~,�f�����1� �������,��I�2�i�7������Gn���   �   ���ز���#��ͺ��~u_��09�x{��pս�=������(aa<�0=H�H=L}{=>��=
��=t:�=ᱧ=-:�=���=���=�{{=��H=Y/=]a<�����>���qսx{��/9�t_�����'"��:���m�������D-��8����e��E��(�ϊ���.���p��x��(�(�|�E��e�^����.��K����   �   +W��Q܎����l2u���U�ڼ1�>y��ϽD��� ��x�>�а3<�0�<�:=8dl=P,�=�d�=�%�=ү�=l%�= d�=\+�=bl=�:=�,�<��3<��>���U����ϽYy�<�1���U�+0u�<���ڎ��U���C���%��d2t��WW�T9������T��"����򽶘����U9��YW��4t�N'��IE���   �   ����zւ�(Lx�ȑb�ȒF�`�&��P���ȽҊ���#���|�0�;�<ax =<fR=T�x=��=@�=���=��=��=��x=cR=�t =�
�<P��;��|���#������Ƚ�P��&�b�F���b�KIx��Ԃ�����v��kes��\���A��&��z� ���ս(p̽��ս|�ｴ{�h&���A�x�\�Qhs��w���   �   Q�i�}�g��]�� L�3�4��	�Q��۝½�d���J4�l���@B��.x<���<�C,=yS=�o=�F�=�=�E�=h�o=^uS=?,=|��<(x<���@���,P4�(g���½R���	���4���K��]�=�g���i�N�b�& T��B?���&����*�콻�ǽ�,��$���r-��7�ǽ{��T����&�E?� #T���b��   �   Y&G���G���@��?4���"�V�������|R�����_���-;D:�<6k�<��!=�r?=d�Q=��W=ıQ=�o?=~!=�_�< -�<��-; `�0��6R���*������&��_�"�p=4���@�T�G��"G��|?�3S1�Q3��?�ͼ��躽zP���U���3|�kV��"R��g뺽@���A��5�>V1�J�?��   �   �i$�,�'�L>%�������2��!��ƽ�ң������><�<���c� :�>[<ʭ�<��=#2=�==0=�=���<�"[< :pd��'��G<� ����֣�<�ƽ�/���������;%��'�nf$������D`���'ѽѩ�ID��0T��/�.#���/��
T�G���ԩ�~,ѽ�e�����W���   �   H��u
����6\����Z:����콠�ֽ ��ᢽ����rM����Ј���ͻ���;Xnj<��<L˲<��<�]j<�r�;��ͻ���,��V}M�^���9梽�$��T�ֽ�콮:�����MZ�?���r
��`��k�׽�ݶ�5�����a��R$�Ā��J���ܓ� O��Ԉ缔X$��b����㶽��׽Ћ��   �   �<н���Ko�����@ �@@ �W����l�(��4:нs����Ú��Zv��5�� z���:û f: �4;��
:�]ûІ���,�Ա5��ev��ɚ�R����?н8���p�����@ ��? �����vj�*���6н𒷽M����Sv���5�x�To�� û��:@,5;�:P4û�{��p �^�5��^v�Aƚ�����   �   䢽#��|�ֽ�콁;��j���[�����t
��r��d�׽Hᶽ����$ b�JX$�H���T���擼dY���缮^$�jb������涽q�׽���!�Hw
���]����D:��̹���ֽ���nޢ�&����lM�B���}�� zͻ@ɰ;�j<`'�<�Ӳ<@#�<�oj<���; �ͻ<�������wM�⌅��   �   Ƽ��֣�*�ƽ�����̴�.��u=%�!�'��h$�@�����;d��v+ѽKԩ�0G���T�.�/�3#�N�/��T�FJ��Tة�X0ѽ�i�����x���k$���'��?%����j��~�����ƽKѣ�����N:<��� �c��>:�O[<Ե�<��=�5=D=�3=��=��<�3[<�-:d���xD<��   �   �R��򓽾������8��ϵ"�8?4���@���G�=%G�??�XU1�G5�{A��㽤뺽�R���W���8|��X���T�������C�8�nX1�~�?�y(G�|�G�7 A��@4���"����h��$����^R�z����_��8.;lA�<,r�<ۅ!=�u?=`�Q=��W=��Q=�r?=/�!=Tf�<�3�<�-;�`� ���   �   �O4��g����½�S���
�l�4�l L��]�f�g��i�o�b�""T�ND?�*�&��������ǽ�.��>����/��� ȽT����~�&�G?�3%T���b�\�i�_�g���]�L�6�4��
��Q����½,d��,I4�ܡ�����9x<��<0F,=�{S=J�o=�G�=6�=�F�=��o=�wS=pA,=��<P!x<@~�,����   �   *�#�J���V�Ƚ�Q��&�֒F�>�b�Kx��Ղ�䩄��v��gs�s�\���A��&��{���ｂ�ս�q̽b�ս����|��&�$�A�$�\�js��x�����Jׂ��Mx���b���F���&�Q�ĵȽ������#���|���;��<Sz =hR= �x=��=��=h��=��=��=.�x=�dR=+v =��<���;�|��   �   @��A���g�Ͻ8z�M�1���U��1u����nێ�5V��[D��u&��V3t��XW��T9�������L��"��$��i��ڷ�sV9��ZW��5t��'���E���W���܎�0��H3u���U�M�1�~y�J�Ͻ)���z����>�P�3<t3�<:=lel=�,�=We�=F&�=<��=�%�=�d�=�+�=�bl=:=2-�<x�3< ?��   �   Z���?���rս.|��09��t_� ����"������Α������-��d���
e�2�E�4�(�ފ�3��p���������(���E�5e������.������c���!����#�������u_��09��{��pս�=�����p��ca<91=��H=�}{=t��=;��=�:�=��=J:�=���=���=�{{=��H=�.=�Za<���   �   �n����~׽F�D�;���b��܂�󛐾�j��&m���l����5����i�>�I�$~,���C��� �������r,���I�%�i�7������?n���n��%l��-���}݂���b�M�;�|E��|׽������8Q��o<��=�M=�9�=��=X�=牧=&��=���=��=��=�8�=�M=��=��o<PY��   �   ���n>��rqսX{��/9��s_�y����!��簖�	���J����,�������e��E�9�(����`������ҝ�ߊ���(�ؤE��e� ���<.��ێ������^���#��V����t_��/9��z��oս�<�����p�xga<�1=\�H=D~{=���=\��=�:�="��=e:�=���=���= |{=&�H=�/=�^a<���   �   ��5�����Ͻ�x�h�1���U�/u���� ڎ��T���B��%���0t�`VW��R9����Ֆ���
����򽴗����YT9��XW�`3t��&��|D��UV��xێ�����0u�f�U�f�1��w���Ͻ���L����>���3<,6�<  :=4fl=&-�=�e�=y&�=t��=&�=�d�=,�=�cl= :=�/�<د3<8�>��   �   ��#�q���ƴȽ�O�s�&�ϏF�эb�_Gx��ӂ�ৄ��t��7cs���\���A�&��x�
���սvm̽��ս���@z��&���A���\�;fs��v��y���OՂ��Ix���b���F�`�&��N�8�Ƚć����#�(�|�`0�;��<�{ =*iR=��x=��=Z��=���=��=��=��x=�eR=�w =��< �;p�|��   �   �J4�*d����½�N������4�Z�K���]���g�S�i���b��T�@?�H�&����D��*�ǽo)�����W*����ǽ��p����&��B?�� T���b���i���g��]��K���4����L����½�`���C4���������Bx<p��<tG,=||S=�o=�G�=��=SG�=|�o=�xS=�B,=p��<�*x<�L�𦲼�   �   R�����8������"��:4��@�v�G� G�z?�fP1��0�@=�<�㽷亽�L��R��-|�S���N���纽�㽞?�s3�zS1�Y}?�E#G�g�G�h�@�q<4���"����������ꓽ�R���h�_��`.;,E�<u�<��!=�v?=�Q=~�W=|�Q=�s?=K�!=2i�<`7�<��-;H`�����   �   ̹��Gң�r�ƽ�轋��ذ�����8%��'�gc$�������Z���"ѽu̩�@��n�S��/�'#��/��T�-C��~Щ��'ѽz`�����I���f$��'��:%�O��v����*��e�ƽ�ͣ�Ĵ���5<� ���c� �:�U[<��<��=�6= =�4=��=B��<�9[< �:� d����?<��   �   Gᢽx����ֽ����4�����WW�=���o
����к׽Hض�\�����a�jJ$��q��<��4ϓ�8A��`z��P$�6�a�Q����ݶ���׽��pr
�r���X�)���3��V�콂�ֽ3���ۢ������iM�ʽ�Hz�� oͻ�Ѱ;��j<�(�<,ղ<�$�<xsj< ��; �ͻ����&���tM������   �   e:н���<k�&����= ��< ������d�X��&1нm������Jv���5����`����» >: �5; �:��»�l��X�v�5�
Uv�����K����6нg�㽬h�W���0= ��< �����jf����P4н����Ծ���Qv��5��xm���û �:�65;�=: .û�y���𼮩5��\v��Ě�����   �   ,�Ut
���Z����r4����d�ֽZ��1٢�!���TcM�p���m��P>ͻP �;��j<�3�<�߲<</�<�j<�ϰ;�|ͻ�������mM�|���Vޢ�����ֽf���4����'X����Wq
������&�׽�ܶ�������a��Q$�X缬I���ۓ��M��\�缺W$�� b�M���ⶽ6�׽���   �   �h$��'��<%���������������ƽṃ����z1<�D��x�c��:�i[<���<F=%;=|=79=��=���<PN[<��:��c���:<�����iУ�:�ƽ��轸��x�����%:%��'��e$�]��)���_��O'ѽ�Щ��C���T���/��-#�v�/�D
T��F��Vԩ��+ѽ�d��4������   �   �%G���G�h�@�>4��"�b�������YꓽnR����_� �.;8M�<}�<�!=�z?=�Q=6�W=8�Q=xw?=[�!=�q�<@�<`,.;��_�v���R��퓽W���#��0����"�<4���@�l�G�C"G�v|?��R1�3��?�u�㽚躽>P��^U���3|�3V���Q��!뺽�㽲A��5��U1��?��   �   ��i���g��]���K���4�}��M��(�½�`���B4�𕲼`��(Nx<���<�J,=�S=�o=|I�=�=�H�=��o=�{S=F,=l��<�8x<������H4�8c��=�½�N��!���4���K�2�]���g�n�i���b��T�RB?�o�&������콊�ǽ�,������H-�� �ǽC��3����&��D?��"T�.�b��   �   r���>ւ��Kx��b�ߑF�P�&�vO��Ƚ����(�#���|� =�;x�<�} =`kR=*�x=��=x��=ƙ�=���=�=~�x=$hR=Hz =@�<� �;��|���#�����j�Ƚ�O�д&�y�F�Ўb��Hx��Ԃ�Ǩ���u��<es���\���A��&��z� ��ˋս
p̽p�սZ�～{�S&���A�P�\�hs��w���   �   W��-܎�|���1u�`�U�,�1�xx�m�Ͻq���V����>�@�3<�8�<t!:=�gl=�-�=Uf�=@'�=2��=�&�=�e�=�,�=fel=:=4�<�3<x�>�N������h�Ͻ�x���1��U��/u����ڎ�gU���C���%��O2t��WW��S9�����D��
���򽪘����oU9��YW��4t�>'��4E���   �   ���ǲ���#������6u_�S09�{�+pս=��0�� ��ha<w2=�H=�~{=��=ȩ�=&;�=���=�:�=:��=X��=d}{=|�H=*1=�da<�	����=���pս{��/9��s_�����"��)���`�������=-��2����e��E��(�ʊ���"���k��q��!�(�r�E��e�X����.��@����   �   ��������0�3�Ӿ�ĸ����w�C@;�8c�K$���+���<��<�J =�(a=�؇=�3�=+��=YS�=Fß=i��=i��=@�x=`UO=��=N��<�|�;��L���
��wj������)ڽ�'�yL���*��D5���8��P5���+�t�T|�������J��g����P1.���V�%ԃ��'�������Ծa龧����   �   .0��1���Zо襵����
's��b8��v��ߥ���)�@"�3�<�
=H:^=<$�=�K�=���=D�=��=�h�=lJ�=�xq=��G=��=�D�<0ԣ;h�d��o��l�a�����ؽ����X�GJ(��F2�Bt5���1�q(���VK�J���6��f�8����K�
g*�PR��6�����hs��ʭо!�o��   �   /�����WپL�ž@���^���T�g�V20�X��g����H$�(��䳉<�=� U=�ހ=e�=/�=��=Ȳ�=j�=��}=@[=P�/=R"�<�Ԃ< ������z��*{u��Z��Q�ս$M �����!�2�)�%�+���'�4k��Y�%�LL콎 ۽�=׽��#��eb��0E��<s�6���B��-Lž��ؾF���   �   ־>pҾ-/Ǿk���ޞ����b�V�h�#�P
꽵������R�x�p<��	=(�D=P;o=��=b��=ۋ='��=�ux=r�Z=��4=b =�d�<0r�;�4!��ܼ|�8��~��4~��2�ҽ��l�
��l������6��m��W@�:�3�н�e�����Hfɽ������1�Ƃ[�f\��d��%���<�ž�Ѿ�   �   ͷ��}���䄰�YM��Y֍���o��B��o���׽���V`�`�4�8�3<>L�<Rj,=�S=��k=Pv=\s=`?d=��J=$(=�v�<��<���;���Ƽ~�"��d����Ї���fҽ7��K��
��r�M�Z�����,�޽�Ľ����U��ä��;ܥ�l!½#�R�eZ=���g�wM���2���z��Vd���   �   �����瞾�����D���v�eR�:X,����>>ǽE��h���=r�P��;�R�<:
=V:.=@VC=��I=��B=B.=yt=�s�<pHL<@�����z�����Zi5���n�ь�����\�ýmSؽ�e�Ȱ��O���R7��}���utͽ${��c���ԅ��n�&Pg�p<z�����Ī��[*���2� �?�fje����t��4K���   �   �䃾�q���|��j�VR��.6�;�Ԇ���#��������+�L��@�`�P�9<Xߺ<�{�<�=3�=��=*��<��<��~;��+��+ռ�N+���i��������[���ѽ��޽��֘�~��Ng�Ԛ޽HeϽ�-���7��雉���a�(�8�T!�H��ƹ#���L�<Y������������2�6��nT�:em����   �   �CQ��S�X�M��B�^�1�`��:�����4]��4݋���G�D{����u�@p��h�<D��< ��<�D�< Ew<��;P��������V��9h������ʺ��׽���X�����������v��>Z�q�ܽ�WȽ����Q���#x��B��T��ϼ(r��(Ȅ��P����ܼnd&��Ms�����^�ܽL	�Bi"��8�H��   �   2q �f%�`�$��S�C��O
� ���Thڽ�����5���s�<�4�`��(-���� ��`�:; �:G���ނ�� ���L�����<��M.齋~�&n��s ��!%���$��U�XD��P
�����@hڽ.���|4����s�d�4�H���$��@�� �����:; ��:P���҂�
 ���L������7���(齸{�Mk��   �   H��T�����M����
v��4Z�,�ܽ$YȽ����S��$(x�RB�\Y�'ϼH{���ф��Z����ܼ�j&�VUs�����L�ܽ	�Ml"�8�WH��FQ��S��M��B��1�������&�� ]��m܋�Z�G�8u��x�u�������<���<��<M�<�Ww<p�; o��<���O�J1h�b���&ƺ�T�׽�   �   ��X����ѽ��޽6�罼��*�콢h轮�޽�gϽ"0��M:��h���xb��8�&�$���#�D�L��\��o���c���#�6��qT��hm�c��惾�s���|�}�j�(XR�"06�#<����0$��d���v�+���� b`���9<V�<��<[=њ=��=0��<0��<�;8�+��ռ�G+�`�i�朑��   �   ��n�ʊ��j����ýJSؽf��������9������wͽ�}��}e���օ���n��Tg�`Az�s�������%.��5���?�\me�����v��M��Y����鞾!���F��;�v��fR�hY,�e���>ǽ4E������7r����; W�<g<
=�<.=�XC=��I=�B=�E.=�x=�|�<�\L<�ꅺ��z�d����c5��   �   J�"�nd�0������hgҽ.L��
��s������v���x�޽&�Ľ����W��Ц��kޥ��#½��S�v\=� �g��N��x4���|��f��|������]����N��h׍�^�o��B��p���׽n���`���4�x�3<fO�<l,=��S=��k=�	v=�s=(Bd=��J=�(=^~�< ��<��;����ż�   �   pܼZ�8�e~��w~���ҽ:��3�
��m�������F��s��IA�����н1g������hɽ���' �"1���[�n]��/e��t�����ž��Ѿ�־�qҾl0Ǿ#l���ߞ�ԉ��k�V��#�%������`P��p<�	=d�D=�<o=n�=4��=e܋=&��=xx=�Z=�4=#=jj�<���;�+!��   �   ���R���{u�n[��*�ս�M ����m!��)���+�v�'��k��Z���SM콄۽�>׽��Ҥ�Ac��1E�>s��6���C��$Mž��ؾS��(0�����Xپ�žᩬ�޷���g��20���������H$�����<��=b!U=߀=�e�=��=���=]��=�=>�}=�[=��/=R%�<,ׂ< 9���   �   ��d�vp���l�	���n�ؽ
��tY��J(�{G2��t5�D�1�Xq(���K�����~�뽸轮����K�tg*��R��6��L���s��P�о�!���0�����徸о2���	��V's��b8�w��ߥ�p�)�0!��3�<I=�:^=h$�=�K�=&��=z�=��=�h�=�J�=\yq=0�G=��=0E�<`ԣ;�   �   ��L���
��xj�=���J*ڽ�'��L���*��D5���8��P5�}�+��s�|�n��<�����������A1.���V�&ԃ��'��!�����Ծa龣�����������/��Ӿ�ĸ������w�@;�c�$����+������<�J =�(a=�؇=�3�=��=:S�=#ß=F��=;��=��x=�TO=�=���<�u�;�   �   �d� o��l�꒧��ؽH���X��I(�~F2��s5�E�1�ap(�(��J��������2�����J�zf*��R�O6������r��N�о� ��~�/�����r徻оT���N��&s��a8�Ev��ޥ���)����5�<=0;^=�$�=L�=G��=��=�=i�=�J�=�yq=��G=��=�F�<pۣ;�   �   �����$xu�PY����սBL �����!�(�)��+���'�j��X��:J콌�ڽ�;׽��-��aa��/E�t;s�Y5��B��<Kž��ؾ&���-꾭�徶Vپ4�ž;���u�����g��00����`���zE$�������<"�=f"U={߀=�e�=��=҇�=���=>�=��}=T[=��/=('�<�ق< _���   �   Pܼ��8��{���{��p�ҽ; ����
�tk���T���������>�b齅�нc�������cɽ�轍�1���[�\[���b��ғ��ģž��Ѿ~־�nҾ�-Ǿ�i��]ݞ�����.�V��#��Ⳗ�D��B���p<��	=��D=�=o=��=���=�܋=e��=�xx=��Z=�4=$=
m�<��;�"!��   �   ��"��d�Q������@cҽh� J�

��p�[�n��P�����޽�|Ľ띭��R��ۡ��O٥�\½��)P�7X=��g�
L��V1��8y��yb��⵼���������K���ԍ���o� B��m���׽����JZ�p�4�H�3<T�<�m,=@�S=��k=P
v=�s=�Bd=��J=P(=P��<���<P)�;X��p�ż�   �   �n�I���K����ý�Nؽ�`�*��������2�����]pͽ>w��o_��Aх���n��Ig�6z�R������2&��z0�D�?�Fge�H��s��/I��x����垾�����B��b�v��aR�:U,����9ǽA��@���$r����;\�<H>
=F>.=ZC=��I=��B=nF.=Xy=�~�<�`L<@�����z������`5��   �   �񪽃U��b�ѽ�޽���z��N��:b��޽�`Ͻ()��}3��ޗ���a��8������(�#���L�qU��D������*���6�kT�Wam����⃾�o��Ҷ|���j�MRR�+6��7�������%���+�0���`(`� �9<.�<��<_=��=��=���<ȣ�<�;�+� ռ�E+� �i�]����   �   h��R��|��v��֭�q���T��ܽ�RȽ��4M�� x���A�FM�ϼ�d��4����C���ܼ�\&�xEs��{���ܽ6	��e"�8�H�o?Q��S�5�M��	B��|1�я��������W��[؋��G��k��`�u� ���x�<p��<�<�N�<�Zw<@�;i������N�0h�����ź�ڎ׽�   �   \p �T%��$�BR�
A�uM
�
����bڽ����/����s��4������`��  ���=;;�|�:�袻�Ă� 
 ���L�}����1���"�9x��g�Tm �z%�w�$�P�Q?�@L
�����Nbڽp����0��֤s� �4���@ ����� �� �:; Ϫ:���dт�^ ��L� ���%7��*(�8{��j��   �   �BQ�S�3�M�RB��~1�f�������	X���׋���G��e��8�u��/�� �<4��<0�<|X�<�ow<@C�;P5������E� 'h��迺���׽V��^M��e��������_o���S�D�ܽ�SȽ���OO���x���A��R��ϼ�o��pƄ�@O��p�ܼ�c&�HMs�T�����ܽ	��h"�p8��H��   �   �䃾�q���|�ƒj��TR��,6�H9�ʂ�����.���+� �����_���9<
�<4��<U=ٟ=-�=z��<அ< w;X�+�ռ�=+���i�������Q���ѽ��޽��罒��9���b�Y�޽�bϽ�+��@6��Ú����a��8�f ����$�#��L��X��K������ͳ���6�gnT��dm�h��   �   X����瞾;���AD���v��cR��V,�
���:ǽ}A������r��Ч;�`�<�@
=,A.=.]C=$�I=x�B=�J.=�}=Ȉ�<hwL<������z�$���Z5���n�`������ܒý�Mؽ~`齊��������4��R��a�@sͽ;z��ob��3ԅ�^�n��Og��;z�x�������"*���2���?�?je�����t��K���   �   ����L�������M���Ս�Űo��B��n��׽Y����Z�@~4��4<^W�<�o,=x�S=2�k=v=�s=Fd=H�J=t(=N��<@��<�R�;@�� �żƷ"�|	d�����؂���bҽb�OJ��

��q�~���� �����޽�Ľ�����U������ܥ�B!½���Q�NZ=�{�g�iM���2���z��8d���   �   �־pҾ /Ǿ�j��wޞ�Ȉ����V���#�o꽷�������A� �p<�	=(�D=D?o=��=~��=�݋=���=`{x=��Z=<�4=�'=�t�<���;(!� 	ܼL�8��z���z����ҽP ��B�
�l����R��ġ���@����нpe��ڱ��(fɽ������1���[�^\���c�����,�ž	�Ѿ�   �   /�����Wپ)�ž���)�����g��10�%�����0F$�8��@��<��=:#U=�߀=`f�=��=���=h��=8�=��}=�	[=�/=�,�<D߂< ������$��$vu��X��B�սBL � ��!���)���+�j�'�k��Y��L�f ۽|=׽����\b��0E��<s�6���B��)Lž��ؾ:���   �   &0��(��	�Iоӥ������&s�Sb8��v�ߥ�:�)� ��5�<>=�;^=�$�=TL�=���= �=��=�i�=mK�={q=�G=,�=J�<��;��d�Bm���l�A�����ؽ$���X��I(��F2�t5���1��p(���JK�2���"��X�0����K�g*�JR��6�����ds��ȭо!�i��   �   <�>�ǀ;��X1���!�����~���^���n�Y�o?��=��֟+�����<�&0=�Uk=��="�=r�=��=�D�=��~=<Q`=x�;=�%=>.�<@�H< #P�Xo��f�2�H�l�I^���f��R๽�|ĽX�ǽ��Ľ~���h���������½�n�5����;���t�����ƾ�~�K��!�7i1�
�;��   �   &�;�/B8��H.�\��
#�#j�+i���9����U�6��ﰽ��'������~�<��.=��h=�
�=eʐ=�:�=l��=D�=үu=��U=�{0="'=���<8�<`m�,r��\��K9�hMq�P]��-��P����(½�Ľ���������@���Rb���ƽ�������y�7���o�g���Wd¾����&��FJ.�:8��   �   l2���.��j%�Q����r�޾�񳾾�|NK��X
�����~P�@F���V�<��*="�a=΁=���=�Ê={m�=\Tv=�Y=�6=|=d,�< �H< �!9P�I��ͼ����N����ꕽ�� ��`����廽�d��FF����������#럽J����н���O,���a�KΑ�����.K��P����~<%�5�.��   �   �#�[4 �����4
�Wu�-q̾�_������;�څ��d����f��z9�
i�<�"=^�S=P*q=(�|=0�x=�'h=�WM=L^*=g=<��<��
<��m������N�4r�lL���u���������౩�_��T޲�� ���������������/؊�%������*�C�f�K��������W]̾����	�a �����   �   "�m��vB� ��].׾����QF��Kd��K'�q��~w������ 7���<�=p?=��U=�iZ=�"O=�X6=�=�p�<4O<�k	��d���ܼ�[ ��M�pGu�(���x����p��@ݫ�����
������䠽�O���7��rqr��5a�T&`�j�v��U����ýb6��H/�se� ё�$���CԾ�Z��E�K1��   �   %�����ټ�Ҿl򸾳���L�~�oMF�E,�8Ƚ� s�����D��N�<F+�<J�!=X�0=��,=�=&�<,��<��;;�MM�p�鼺5��tp�������������UƽTǽ�ýX������ql�����䁽6k_�Ҁ?��)���#���4��a��4����ѽ�+��>�*�s���d���p;v�^��   �   �ʾ=�Ǿ���7r���O��@z���oW�
)�����zꮽP�X�ĎӼ�僻��L<޳�<L��<\[=P��<� �<�\<���(�̼�:6������a���̽�&轾����V���:	�.���<����ӽ���*����;��.d��=5��r��~⼨	˼f޼8��L�S�4q����ڽN���=B�{�r�Id���S���"���ž�   �   �8��8��^I�����=�z��W��!3������ؽ�˚�:vH�|�׼ ���0�;�o<⠘<$��<p:< p�8�R��V��p�����ݽ7������**�
3��r6�g:3�s�*�4��G���O����ѽ�������P(N�,3�P����q���%��D,�@ш����.�F�B!���ٽ'���V9���`�"|��1L��w����   �   {�t���t�X�l�:=]���G�j�.��%��5��%��
ʍ�~�D���� �o���f� �O;�ա;�'�:P��􈼼�e2�B;��8�Ƚ�Z�e2$�R�A���Y�<}k��t�)u�4�l��@]���G���.�:'��7��&��tʍ�"�D�����o���f���O; �; ��:h��T|��(^2��6����Ƚ�W��.$�H�A���Y��xk��   �   Z{3�o6�>73���*�������^M��*�ѽ����+����)N�"5�`����q�p�%� U,��ڈ����F�q%���ٽ0��XZ9���`�g~���N������_;������K��������z���W��#3�`��k�ؽ�̚��vH�4�׼���A�; %o<@��<���<�:< ��8DE��N���p�M誽P�ݽʛ�B��'*��   �   ޳���S�o��!�݆�����:�ӽY������<���/d�0@5�|u�4��˼xn޼$�� �S��t����ڽ����@B�F�r�wf��$V��=%��\ž�ʾڦǾ���[t��xQ���{��rW��)������뮽j�X���Ӽ�ރ���L<��<���<�^=4��<�	�<hs<�j�@�̼R16�����/\��$�̽� ��   �   ���槶�t ���Rƽǽ��ý��������l�����@偽�m_�ރ?�:�)�z�#�Ȣ4���a�Z7���ѽ.�7>�`�s��Ö��f��s;�x�<a�����?�N��1ҾH���7�����~�,OF�t-�~9Ƚ6"s���ἠ>��P�<p.�<Z�!=��0=�,=�=v�<$��< X<;�0M�D���5��kp�����   �   ��M��Au�����y����o��nܫ������
��E ���堽"Q��=9��Ttr�9a��)`��v��W��T�ý�7��J/��ue��ґ��%���EԾ�\�G��2�k�����C�,��0׾���nG���d��L'����Qx�����`5��<�=�?=��U=ZlZ=�%O=2\6=N�=�z�<JO<����d�X�ܼU ��   �   LF�tn�TL�^�u�𲍽�����������߲�{!��Ҹ��3���[���]����ي���������,�tD��K���������^̾?���	�n!�����#�f5 �����5
��v�br̾�`��e���;� ���#���"g�`|9��i�<x"=t�S=�+q=�|=X�x=N*h=�ZM=�a*=P=���<�< �m������   �   ؎I�� ͼ
��N�����ꕽy���������滽�e��G������\���	쟽K��,�нN��P,���a�ϑ�����NLྏQ����B=%���.�52�S�.�Dk%���o�H�޾��:�+OK�Y
�&����P�0F���V�< �*=ća=�΁=4��=xĊ=En�=<Vv=D�Y=P�6==�1�< �H< j$9�   �   @�l�(q�����&K9��Mq��]���-����@)½d�Ľ���y���n�������b��ǽ�N��_����7�a�o�Օ���d¾n��������J.�w:8���;��B8�II.����H#��j�ri���9��)�U�\��%ﰽ��'����<��.=�h=�
�=�ʐ=;�=Ĭ�=vD�=��u=��U=}0=7(=���<�<�   �    TP�x!o��h��2�.�l��^��Zg���๽�|Ľi�ǽ��Ľ`���h��f��r��ֿ½�n�.����;��t�%����ƾ�~�K��!�:i1��;�7�>���;��X1���!�}���~���@���9�Y�B?��=��f�+��쳻�<�&0=�Uk=��=�=`�=��=mD�=d�~=�P`=�;=Y%=.-�<��H<�   �   ��l�4o��t���I9�Lq��\��c,�������'½�Ľ����&���"��T���fa���Ž���ག����7� �o�����c¾P�O������I.��98���;��A8��H.����"�pi꾎h��	9���U�������'�P馻��<��.=��h=�=�ʐ=*;�=ڬ�=�D�=��u=�U=X}0=�(=���<X�<�   �   ؈I���̼��.�N�r���蕽W��\�������㻽 c���D��!������韽~H��T�н���N,���a��͑�ʬ��-J�SP�J���;%�j�.��2���.��i%����:�9�޾����MK�tW
�����\M��1���Z�<t�*=��a=�΁=u��=�Ċ=tn�=�Vv=��Y=��6=�=3�<��H< �%9�   �   8B��k�$L���u���������������۲����J�������筐���֊��������B(꽼A���K����a����[̾Ձ�)�	�X�����#�93 �����3
�ys�o̾�^������;�����ţ��*b� B9�o�<Y "=��S=�,q=��|=޹x=�*h=D[M=<b*=�=2��<P
<`�m������   �   F�M��>u�ɛ��0����l��M٫�^���#��3���ᠽ�L��5��lr��0a�R!`�\�v�&S����ý�4��F/��pe��ϑ�T"���AԾJX�D��/�����)A�����%,׾�����D��td�kI'����Ft������� �\�<=�?=��U=4mZ=�&O=�\6=�=�{�<�LO<���`�c�h�ܼ6S ��   �   ����B���f���.Pƽ
ǽ"�ý����]��eh���������d_��z?�$�)�:�#��4��a�K1����ѽ�)��>��s�8����b��/n;Ss⾦[�8�����	��`
Ҿ𸾒�����~�OJF��)��3ȽZs��������W�<j3�<0�!=D�0= �,=e=��<|��<`c<;�-M�X���5�Fjp����   �   ����.S�g����܃��Z��_�ӽ&�������j7��h&d��65�l�|r���ʼLZ޼����S�Ym���ڽ���z:B���r�b��<Q������ž�ʾL�Ǿ����o��3M��x���kW��)������宽Z�X�<�Ӽp����M<,��<:��<�_=(��<��<0v<e��̼�06�����[��Z�̽���   �   �z3�Jn6�H63���*�������I���ѽ��������d N��+� ��0�q��%�`-,� ň�|�８�F����hٽ��!S9�\�`��y���I������6��j���F��k���}�z���W��3�����ؽ�ƚ��mH�0�׼@{��\�;/o<ʪ�<T��<�:< $�8�C��^M��p��窽��ݽ�������&*��   �   ��t�G�t��l�-<]���G���.��#��1��!���ō��D�Ď�so��<f��JP;0 �;�n�:k��m���U2��1����Ƚ*T��*$���A���Y��sk�[�t���t�U�l�u8]���G�d�.�"�@/�7 ��1ō��D���h{o�@if� P;���;�׮:����z���]2�[6��j�ȽXW��.$��A�_�Y�bxk��   �   �8�����I������*�z���W� 3�f��>�ؽ1Ț��nH�t�׼ v��m�;@:o<���<��<(1:< V9(6��>E�V~p�c⪽��ݽ��'���"*��v3��j6��23�o�*�������F��0�ѽ����z���H!N��-������q���%�H?,�0ψ�D�０�F�� ��hٽ���V9�f�`�|��L��N����   �   �ʾ�ǾB���q��8O���y���nW��
)�����w箽�X���Ӽ𱃻�M<���<��<ic=r��<��<��<P-滠�̼2'6�ڬ���U��,�̽o�9���$P����n����A��7�ӽ����0����7��(d�N95�To��y�\˼�c޼b����S��p��O�ڽ.���=B�\�r�:d���S���"���ž�   �   ���t򾦼徾Ҿ�M���_�~�fLF�!+��5Ƚ�s�`�� ���Y�<�6�<W�!=�0=d�,=y=b�<ث�<@�<;XM�\�鼀�4�p`p�� �������������tLƽǽ�ýF������mh������ၽ�g_�@~?�
�)���#�4�R�a�@4��j�ѽ�+�z>��s���d���p;�u�i^��   �   �a��eB�� ��".׾e����E���d��J'���㽉u������`� �D�<> =D?=�U=�oZ=�)O=�`6=[�=v��<�dO<����c�@�ܼ�K ��yM�f7u�����f����j���׫�t����������⠽N���6��~or��4a�V%`���v��U����ýN6��H/�se��Б�$���CԾ�Z��E�D1��   �   �#�S4 �����4
�/u��p̾�_��v���;����������c�@J9�No�<!"=��S=8.q=��|=D�x=�-h=�^M=,f*=L=暦<�<@>m�<x�� 7Ἤf�lL���u���������������"ܲ����g������o��������׊�㊘�����*�C�W�K��������T]̾z���	�^ �����   �   i2���.��j%�H����T�޾�񳾔�NK�6X
������N��6���Z�<Đ*=t�a=\ρ=" �=xŊ=no�=�Xv=D�Y=��6=�=Z:�<��H< h)9�yI���̼~��l�N�@��蕽���\�������份�c���E��Q���/����ꟽ�I��ܚн���O,���a�FΑ�����,K��P���|<%�2�.��   �   #�;�.B8��H.�Y��#�j�i��w9����U������'��즻�<��.=��h=X�=ː=�;�=`��=$E�=d�u=��U=(0=�*=Ȕ�<�<`�l��j��h	���G9��Jq�\��,��l���(½b�Ľ*�������������6b���ƽ�������t�7���o�e���Ud¾����&��EJ.�:8��   �   󮉿>���$��! j�N� �.�~��ݾE2��x�h�>�My��ԗ� <�8�>�<|�9=8�i=n��=|B�=H��=�q=��W=E8=�=Ь�<��<@�< 90:�Pⅼ��¼�������2&��]2�X8�p9���8�;��2G���e��T������ k�ƞ;��P���)��������-�/���N��bj�.��(>���   �   d^������D�{�Z0f�-�J���+�̡��پ�O����d��_��«��I��[:(8�<�48=\�f=J~=��=��z=D<g=P�K=He*=��=�5�<x�a<�9�;ৈ�_K�|�����ݼ���$��,�&�5�(`9��x8�~	6���6��A�`_�Rb���⼽�a��7��}��⪾܊߾�`�2�,��K��\f���{�M����   �   #���c�|�o���Z�Mx@���"� ��r�ξ����g�X�p"��)��� ��X�:~.�<v�2=|7\=�o=b�o=�\a=�H=#�&=�C =�.�<�p0< _/:��P]��@�̼ X�����)�^�6��n>��@��W=��`6���.��J+��g2��)L�;�֮����],�d�n��_���uӾ����#���@��Z��To��|��   �   �<l�!#h�V�[��H�۷0�p���W�캽�� ���CF�;� ����Y輠�d;���<�=(= 
J=l�T=�M=<�5=E=|��<�=a<���:�Y.��Գ�2���%�&	@��S�R0`�*f�:�e�.>`�>�U���F�:�5��Y%�����|��3/�|9^�sԘ�-dٽ~����W�Ê������{��v��Tb0�mH��[��g��   �   1zQ�9�M�8&C��<2���������׾F���$z�:P/�h�ὺY{��ɾ�@�;v��<o�=��.=��.=�e=�<�<���<�@d;X{?��f޼V�+��a�ra��������3?��hY��ȵ���;���Ԋ�T�x�XY�"�9�<`�n��W �����`1���y�|�������:��s�rȨ�1�־��� ���C1�cB��~M��   �   9C3�gS0��/'�����l���@F���|��:�V��,�]���hR�L�����;���<���<��	=p�<z�<�+<p<�ĂӼZ;�#���/�����ͽ���@p���s���K��t�����ʽ����vz����y��WG�t����Њɼl;ʼd����9:����%OԽ�j��T�I獾m���X�߾��� '��&���/��   �   �����jG
�������޾���?����p��3��E��ن��>,���l�0%�;LԐ<���<�C�<�On< �:0���\����>������qa�M�"���1�X4:�̞;�W6�x3+��u�l��W1�����=���>b���!�\(ݼ���@��������G��,��Vb��(��c�YE�� l��3�ؾ�/����A���   �   �U�4���ܾvʾ�ݲ��.���y�hKC����N̽f^��d�h�G�  G;@7:<`5R<p��;�d亼�@�FV���ݽK
���4��T�n�M��<}��E��ѳ}��Dk�P�R��6�x���3��?��Æ���4��hۼ�k��X������rb�d�缰VQ�Nᨽ�%���\-��c�>K��f`��J�þ�7ؾH���   �   +���g���N��hɜ�T2��0>n��@D�2���齅F����U�0y�БF�@w�� �G; r�9�����ټ~!Q�"ר��l��Q�%���R��N��ѓ��1���P��I.���j��|Q��̜��4���An��CD�e�ҕ齋H����U��z�0�F��H����G; 4�9�t�@�ټ�Q�Ҩ�Zf����%�\�R��I��Γ��.��IM���   �   z������}��@k���R�~6���
0�[=������J�4��hۼ�k�h�����x�b����v]Q��娽<+��`-���c��M��Nc����þy;ؾ���4Y뾱7�/�ܾyʾHಾ�0��A
y��MC�����P̽�_���	��G� /G;?:<XAR<���;�Ē�`ֺ� @��P����ݽr�)�4��T�<�m�����   �   �/:���;�3S6��/+��r����-�b���;���<b��!�P)ݼl��H����h��L
G�v0���f��(���c��G���n��Mپ,3��̙�6��y��α�4I
������޾?
����Y�p��3��H������@,��l�)�;Dא<��<�J�<bn<���:|���V|�����櫶����q]��"���1��   �   ui��hm���E��1��#�གྷ�ʽ����x��J�y��VG�������(�ɼD@ʼ���>:�ѽ���RԽ*m���T� 鍾�����߾L���(��&���/�1E3�PU0�s1'�V��>n�9�� H��c~��R�V�3.��^���jR�$�����;ƾ�<F��<�	=�!�<��<XC<P�|qӼ�O;�s|�����ͽ����   �   	��ڞ���:���U������19���Ҋ���x��VY���9��`�6o��Y �J���c1�f�y����Y���:��v�-ʨ�R�־���u��[E1��dB�n�M�|Q���M��'C�>2����ȵ���׾WG���&z��Q/�4���[{��˾���;���<ɓ=��.=d/=oi=�E�<���<`�d;�\?�TU޼��+�(�a�[\���   �   �%��@�6�S�<+`�f��e��;`��U��F�X�5��Z%����~��5/�<^�֘�Dfٽޘ�l�W�������}������c0�inH���[���g�}>l��$h���[�Z�H��0�V��DY����y!��
EF��� �����[� �d;`��<�>(=�J=t U=0M=��5=I= ��<�Sa<�s�:x?.��Ƴ�(���   �    U��x�̼�T�"��l�)���6��m>���@��W=�Ja6���.��K+��h2��*L�'�׮�_��^,���n��`���vӾ}����#���@��Z��Uo��|�����r�|��o���Z�y@���"����3�ξ}���+�X��"�!*���!��T�:�.�<�2=l8\=0o=�o=
_a=H H=�&=�F =n6�<h�0<�r0:����   �   𙈻�XK����`�ݼ���~�b,�$�5�X`9�4y8��	6�d�6���A�"_��b��d㼽�a���7�ɐ}�㪾�߾a���,�yK�%]f�5 |������^��������{��0f���J���+���j�پ�O��׻d��_�ë��I��\:�8�<<58=Ԑf=�J~=+�=��z=z=g=��K=�f*=o�=�9�<�a<�H�;�   �    �9`<��ㅼ@�¼̦��(�^3&�^2�XX8�Np9���8��;��2G�t�e��T�����	k�ٞ;�Q��*��ε����?�/�¦N��bj�	.��*>��񮉿>���$�� j�N��.�f��ݾ 2��8�h��=��x��r�� ��8?�<��9=<�i=j��=pB�=<��=�q=x�W=�D8=�=0��<��<��<�   �   ����0VK�0~��x�ݼ���^}��,���5��^9�lw8�6���6���A�_��a��⼽#a���7�z�}�=⪾p�߾o`�ގ,��K� \f��{����^��2�����{��/f���J�:�+�b��g�پ'O����d��^�����H���:J:�<�58=@�f=K~=K�=��z=�=g=֜K=g*=��=:�<@�a< L�;�   �   S���̼*S�P��F�)�4�6�k>���@��T=��]6��.�@H+�&e2��&L��쀽hծ�H��$\,�?�n��^���tӾ?��>�#�ʣ@���Z��So�Т|�����A�|��}o���Z�]w@��"�L��G�ξ�����X�F!��'��� ��:T2�<>�2=J9\=�o=��o=l_a=� H=i�&==G =47�<8�0<��0:����   �   h%�� @�(�S��(`�f���e�*8`���U���F���5��U%�����x�L0/��5^�Ҙ��aٽ.����W�����Ƞ��:z��|��.a0��kH���[���g�f;l��!h���[���H���0�T���U�`���h���AF��� �����Q��e;,��<X@(=�J=NU=�M=�5=�I=���<hUa< ��:�<.�(ų�"���   �   O��ᝢ��9��T��ܰ��#7���Њ��x�hQY�>�9��Z�*i�VS ����\1�̕y��������:�rq��ƨ�<�־k�����)B1�caB��|M�TxQ�a�M�r$C��:2�%��c����׾.D���!z��M/�����S{������;~��<ӕ=D�.=X/=-j=�F�<ʺ�< �d;�Z?�(T޼>�+�B�a��[���   �   �h��`l��`D�����4��J�ʽ���u��n�y��PG������H�ɼ|1ʼT����4:�����KԽ�h�?�T��卾I�����߾<��n%�� &���/�3A3�eQ0��-'���9k����C���z�� �V�'*��X��bR�Xv��@?�;Ŵ<η�<�	=$�<��<�E<���dpӼdO;� |������{�ͽ&���   �   �/:��;��R6�,/+��q���!+轞|���8��b6b���!��ݼ, ����~�������p�F�+)���]��(���c�.C��fi��.�ؾE,����E��x����yE
�����r�޾�����z�p�_3��@��w����6,���l��N�;�ݐ<R�<N�<�fn<���:$����{�m�������7��D]���"�@�1��   �   Qz��d��O�}��?k���R�p6���d-�:��������4�d[ۼ��j�p,���{��[b����HOQ��ܨ�( ��&Y-��{c��H���]���þf4ؾ��徦Q�H0�(�ܾ�rʾ�ڲ��+��%y�tGC�����H̽�Y���x�G��wG;�K:<HJR<��;�����Ժ��@��P��X�ݽR��4��T��m�n���   �   �*��Ng��KN��ɜ��1��A=n��?D�����C����U��l��wF� ���`-H; ��90\�0tټQ��̨�`����%���R��D��˓��+���I���'��
d��7K��HƜ�~/��'9n�Q<D�~�|��SA����U��jＸxF�@¢��H; 9�9o�L�ټ�Q��Ѩ�f��h�%�C�R��I��Γ��.��,M���   �   fU��3辥�ܾ�uʾ_ݲ�R.���y�cJC�����K̽�[����p�G� �G;HS:<(VR<��;0���0Ǻ��	@�RK����ݽ����4��T���m��	���w������ �}�!;k���R�6�)��M)�7�������4��Zۼ�j�p;��В黠kb�����UQ��਽n%��p\-��c�4K��Y`��<�þ�7ؾ2���   �   w��د�XG
�`���t�޾��������p��3��C�������9,�ؗl� P�;z��<�<�T�<�xn<���:�~���r����S�����@Y�t�"���1��*:���;�[N6�d++�On�0���&�uy���6���3b���!�Tݼ�����l������G��,��b�{�(���c�PE���k��*�ؾ�/����9���   �   2C3�_S0��/'�����l�����E���|���V��+�J[��eR�8y��@=�;�ƴ<B��<Ĭ	=h+�< ��<�]<���_ӼFE;�av��.�����ͽ��va��ge���=�����&��"�ʽJ𱽐s��r�y��NG����P�𼴃ɼp6ʼ�����8:������NԽ�j���T�>獾e���P�߾���'��&���/��   �   0zQ�5�M�3&C��<2���������׾�E��F$z��O/����V{�Xþ�P�;T��<�=L�.=>/=�m=>P�<&Ǝ<`e;x;?�xB޼t�+���a�YV����������4���O�����4��=Ί���x�|OY�t�9�([�Rj�*U ���0_1���y�,������Ԓ:��s�kȨ�+�־�������C1�cB��~M��   �   �<l� #h�R�[��H�ѷ0�c���W�ú��x ��|CF��� ����U���d;p��<$A(=2J=\U=�M=t�5=�M=���<�la<�Q�:� .����V���
%�l�?��S�l"`��f�F�e��4`���U�Z�F�h�5�>V%�ܣ��z�~2/��8^�!Ԙ��cٽl����W���������{��t��Sb0�mH��[��g��   �   "���b�|�o���Z�Hx@���"����Z�ξ����"�X� "��(��r����:.2�<��2=$:\=,o=H�o=�aa=l#H=��&=K =�?�< �0<��1: ���H�� �̼xN�"����)�N�6��h>� �@��S=��]6���.�:I+��f2��(L��퀽�֮����],�X�n��_���uӾ����#���@��Z��To��|��   �   d^������C�{�X0f�+�J���+�ȡ�
�پ�O��p�d�y_��«�I���:�9�<68=��f=�K~=��=��z=?g=��K=i*=Ϡ=�>�<��a<�a�;���HKK�y����ݼ����{�� ,���5�4^9�Xw8�R6��6���A��_�*b���⼽�a��7� �}��⪾؊߾�`�2�,��K��\f���{�M����   �   O8��4���O���X���4����ss��uG�P���n�f̩�<f�������|��p��;FH�<��8=t<X=X�`=hlX=<<C=��%=<�=bӻ<��e<��;�NѺ0'����K�h.��@��<ۜ�9���햼���\=���Us�l=����!��:�.(���[�z�-��j}�&�������@�I�Δt�YI��K桿���������   �   �#��z�W������򘌿lo��D��=��Y��Φ�>�a����G���$ڼ�V�;���< >5="eR=�X=��M=�;6=p	=���<�B�<��< D�������c_�86������lj��XϿ�]���	��pA���Ӌ�#����������缄�5�WY����: *��}x��?��B��.o�m�E��hp�����6��ᨭ�D�   �   �.��h+���P��	p��;ȅ�W�c��c:��~���ܾ$��8�U���C��>ż���;��<�**= �@=5@=`.=��=
��<�1h<�=;�s���@aӼ���|H�Vr�$��R����	�4J���Ҽ,!����剼������ռ�j&�]��`�ѽ���1j�����
��hA�>~;��Jd��ᅿ}e��I6������   �   �%��zf��5=���j��i/v��UQ�92+�yj� ʾެ����B�4Q���{�P~��X�
<�u�<0�=*5"=R6=�s�<��<��;�M�����wE�3k��e��V̈���������@s�x_X�89�tc��z�����l�������=������h����RM�-�S�I�����;����+��[Q���u�\*��,����=���   �   G:���Ύ�Ɔ��Vx��Z���9���RH�.ܲ��u�?B+�(ѽ�AV�@d��PT<x�<���<b��<P*�<�&<�:������y,���y�p���Nݾ�/\ս<�⽊�潲�@�ӽ�`��}���R����_�N<+��_��ܖ��P���hs���^鼐�>�.�������7�Ez��n���x�� ���K9�Z�Q*w���������   �   ��y��u��i��?U�\<����V>��̾o蘾��Y�S������W.��D�@W�;Xi�<83�<p]h<�;�Zz����{�ZN���L���
�u�5h,���3���3�X-��� �	������8�̽��n�s� A-��,� Ԣ�8΋�@�����f�t���ŽRz�9�[��f���]ʾ����}:�V�S���g�;u��   �   ?O�\�K��bA��0����PD���׾�ᨾ��|�*3�(�콑t��������F�;`�*< ��; �����eB�(ԝ���὞b�QO7���V���p��B��^���o��Ba}���i�rO��[1����������(p�P.���¼쯁�H��ż�M/�H��T ��1/�Tv����L!Ӿ���m�� /���?�rK��   �   É%�v�"�I����������Ӿ]Ƭ�m.����I���� ���^8Z��Ѽ`��@ԃ: u�9(���lݼ\�Y�ha��QH�Pw.���]��$��� ����(~���M���$��[S���̢�����}:u���H�^>�Jg��C��l�T��&���8���*2��d���ټ.�J�����h�>�<�>������;W�� �T��"��   �   ����� ��c��X�ھ(����᣾�х��wQ�h7�@�۽���^~%�����P6�����8�D��T��O[��^��T��X�<�#�w�ɚ�����pԾ�g����:����$������ھn����䣾ԅ�0{Q��9�ܕ۽t����%�|����3�����h�D��I�PH[��Y����)�<���w�ƚ�����lԾ�c꾕����   �   �I��� ���O���ɢ������5u�ڦH�|;�c��@����T��"��8��0/2�X�d�h�ټN�J�0����j��<����󣥾;W���"����"�Q�%��#����ߘ�`���'�Ӿ�Ȭ�`0����I�É�㟺��;Z� Ѽ`����: �9(��D_ݼ��Y��[���D��r.���]��!�����n��Wz���   �   �Z���l���[}�h�i��mO�X1����Z�佪󪽢p��+�l�¼l������żR/�����$��4/�:
v�����`$Ӿ������|/�p�?�K��!O���K�AeA�A�0�����E���׾�㨾��|�J,3�/��qv����� ��0O�;�*<���;��������V\B�:Ν�j��W^�hJ7�Q�V���p��?���   �   ,�3���3��S-��� ����N�����̽���l�s��=-��(�$Ӣ��ϋ�����0���t�=ƽ�|�6�[��h��_`ʾR�� �=:���S��g��u���y���u�i� BU�P<�d���?�̾�阾ҵY�� �
����Y.�ȳD�p\�;�l�<d9�<@oh<�j;(<z�|��2{��G��JE潎�
�vp�oc,��   �   "�⽪��J�z}ӽ�[��P�������_��8+�[������$���(u��`b鼞�>�^�����ƈ7��{��G���Ժ���M9�Z��,w����ϓ���;��Ў�凇�a x���Z�H�9�F��>Jݲ��w��C+��	ѽDV��e��xU<�z�<|��<0��<�3�<P*&<` ��t��bo,�0�y�
���y־�Uս�   �   �`���ǈ�h��������9s��YX��39�`�(v�d����k������?�������h�����N���S�}�����;����+�&]Q�j�u�K+��*����>���&��wg��#>���k���0v�(WQ�:3+�Ck�/ʾ������B��R��{������
<�w�<͵=�7"=�9=8|�<�<�:�;�0��Ἴ��nE�0)k��   �   ����B��l�P��0��(�	��D��}Ҽ���0피p剼H���L�ռPl&�
^����ѽ���2j�t���?��,B�+;��Kd�Cⅿ,f��7�����s/��,��pQ���p���ȅ�2�c�8d:��y�ܾ�$����U�e���C��?żP��;2��<�+*=��@=07@=.=�=��<8Dh<`j=;0]�����TӼ�   �   pX_��0��䔮�(f���˿�8Z������?��Ӌ��"�����8�����V�5��Y��f�� *��~x�@����o���E��ip�Iጿu6��E����"$���󶿪���8��/���flo�D� >�$Z�Ϧ���a�;���G���$ڼ�W�;4��<�>5=�eR=�X=��M=�=6=Y=J��<�G�<X�< `u������   �   @*��8�K�P/���@��,ܜ��9�������=���Vs��=����!�.�:�M(���[潛�-�1k}�F���$��A�(I��t�eI��T桿��������O8��/���F���J���%����ss��uG�3���n�<̩��f�T��������ἠ��;�H�<��8=�<X=\�`=\lX=4<C=��%=�=ӻ<ȏe<� �; XѺ�   �   W_�$0��ܓ���d��\ʿ��X������=���Ћ�, �� ��\���̜�l�5��X�����*�>}x�3?��ہ��n��E�whp������5��������^#���򥭿�������_ko�=D�q=�Y�CΦ�Z�a�h���F���!ڼ�`�;П�<?5=LfR=X�X=�M=�=6=t=���<H�<�< �t������   �   ���A��k���̒���	�8A��yҼP���蔼\���Ў��4�ռ�h&��[�� �ѽ;���0j�՗�� ���@�}};��Id�ᅿ�d���5��&���-���*��P��[o���ǅ�<�c��b:��}�q�ܾ#����U�ΰ�fA���8ż@ <0��<�,*=H�@=�7@=n.=Y�=���<,Eh< n=;\�`����SӼ�   �   R`��ǈ��������7s��WX�19�P]�p����d��`�,7�������h����L���S�B�����;����+�^ZQ�4�u�)��9����<���$��qe��7<���i���-v�qTQ��0+�ri�_ʾ������B�<N�D�{��v���
<�{�<B�=�8"=O:=0}�<��<�=�;�/��༼����mE��(k��   �   ����潄὆|ӽ�Z����������ʼ_�,5+�hS��<��������j��LV�4�>�����������7�y��ʷ��_��М�GJ9�<Z�;(w����_���	9���͎����� x��Z��9�����E�Eڲ��r��?+��ѽ~<V�4[��(d<��<���<���<5�<�,&<�������o,���y�֩��,־��Tս�   �   �3���3�\S-�;� ���߮���̽������s��9-���ɢ�ċ���������t���Ž-x�q�[�e���[ʾX �=�{:��S��g���t�D�y�d�u�i�=U�2<�ܓ��<�[
̾^显^�Y����7����Q.�X�D��|�;�r�<*=�<dth<�y;�9z�����{�hG��E�p�
�Pp�@c,��   �   �Z��`l��:[}��i��lO�[W1������佮�Np��&��¼���� �~�D�ż�G/�������./��v�����fӾ<��a����.�X�?��	K��O���K�,`A���0����kB���׾5ߨ�R�|��&3���~p��|z�����p�;��*<���; ���<����[B��͝�0��=^�LJ7�7�V���p�z?���   �   �I��� ���O��bɢ�����65u��H��:�&a��>��(�T�����,��`2���d���ټ �J�����Re���<���Q���Y ;w��m�����"�)�%���"�Ϻ�t������s�ӾQì��+����I���
���(0Z�xѼ�������: c�9����\ݼ��Y�c[���D��r.���]�x!�����_��Dz���   �   ����o ��>��(�ھ�����᣾�х��vQ��6�_�۽����y%����H�0b����D�$<�@[�}T��ɭ��<��w�Ú�v���hԾQ_�������������2�ھl����ޣ�υ�,sQ��3�8�۽?���nv%�@}��@��p��0�D�`F�0G[�DY�����<��w��Ś����lԾ�c꾇����   �   ��%�m�"�<�����}�����ӾƬ�.����I���N���@4Z��Ѽ����@��: ��9 ��HPݼL�Y��U��/A��n.�u�]����=�����pv���E�����	L��Ƣ�����:0u��H�r7�]\�b;����T����,+���2���d���ټ��J�z����g��<�2������;Q�� �P��"��   �   <O�W�K��bA���0����9D���׾�ᨾ�|�e)3�����r��}�h��0v�;8�*<��;`a��ﺼ�RB�@ȝ�-��Z�zE7���V���p�]<���W��Di��VU}���i�;hO�XS1�t��p�����p��#���¼����@���ż�K/�����콢1/�8v����D!Ӿ���j�� /���?�nK��   �   ��y��u��i��?U�O<����@>��̾4蘾�Y���������T.�`�D�p~�;�u�<�B�<0�h< �;(z������z��@��u=�.�
��k�c^,���3���3��N-�� �Y��������̽������s��5-��@Ǣ��ċ�Ȣ��ҭ���t�{�Ž*z��[��f���]ʾ����}:�U�S���g�;u��   �   H:���Ύ�ņ��Rx��Z���9����0H�ܲ�Fu��A+�ѽr?V�$^���c<���<"�<��<�=�<�C&<�ë�h��d,�,�y�^���0Ͼ�jMսD���}潦�?vӽ�T��V��������_��0+��M��X���@���8l���Y���>���������7�<z��f���r�����K9�Z�R*w���������   �   �%��zf��6=���j��f/v��UQ�/2+�nj��ʾ����J�B�lP� �{��y��p�
<�|�<��=�:"=�==���<B'�<p�;@�(м�^~��cE�*k�[����������P���0s��PX��+9�8Y�@j�0�c��l񔼨8��.����h����2M��S�A�����;����+��[Q���u�]*��+����=���   �   �.��i+���P��
p��:ȅ�T�c��c:��~���ܾ�#�� �U����{B��0;ż�  <���<x-*=ʨ@=�9@=(	.=��=���<lXh<��=;�C�x鐼xFӼ6��$;��e�P�����,�	�<:���sҼt��H攼`߉� ���d�ռ�i&��\���ѽ����1j�������fA�<~;��Jd��ᅿ~e��K6������   �   �#��{�X������񘌿 lo��D��=��Y��Φ�"�a����VG��L#ڼ�]�;ܟ�<|?5=�fR=f�X=��M=|?6=�=p��<zM�<8�< xg��n��(I_�D)��<����^���Ŀ��S��,���:���΋�������t���|�� �5�(Y��v�0 *��}x�~?��B��-o�l�E��hp�����6��ᨭ�E�   �   �8�����;��"�տ����C��[ƅ���S��!��꾌Ρ��*R�Ĩ���u� ��T�U<$��<�X&=��0=o�&=@t=�<�<X��<��;�P�P�:��0��HH����ȼ��ɼ ~��Ds��8	y��J(��p��@CҺ  �8@��Ƚ���ü|YI����/��SKf�������F�#�VV�;������������տ
��R���   �   �;��M���\ҿ����᩟�����yP�[�}�e�PN����o������!Q<��<ax=\%'=G�=P��<�Q�<�"0< @/�P�%��:��8�ѼDN��`��p�����,�м�쥼p�l�0+��ڄ���̺ 61� ����ēD�����9��h�a��禾���~!���R��t��/L������U�ҿ����   �   ٩�'��GbڿI�ȿ�б�����{z�v:F��n�bSھ&����C�;��<`��|n�B<���<;}
=bC	=���<Tb�<�s�;�ʻ���:} ��*��J�(c]���c���]���L�Ā2�s�l߼�N��0�=���ۻP6���-&�T���%7�t�����T�>Ý���߾����G� �{��t������zȿ<ڿ����   �   V�׿lԿk�ɿ������'��ӈf�w,6�B
�4Ⱦ~����1���ϽZ�H�0�R���"<;�<��<�\�<��=<����f����B�V�c���{a�������;Ľ��Že/����������if��0�J���t�ʼ�����4���E�U���l#��������@�n���Y̾]���/7��g�[-���֣�+���O9ɿS�ӿ�   �   �����t������G���Y����y�tM�D�!����� ڰ�˵r�L��yP���|,�p�:�@;�;�bb<=F<�B;��F����X�]������Ͻ�%��!_����N�!��9!�g7���H����@ҽ��������5�t�䢟�pր������hz� ,ӽ0O'���z������"����!���L�z
y�Qґ������j!���   �   �R��x������������O|���V��0��
��AѾז��N��5�����>���K1���:�:);�
���E����3��Ⓗ'ӽl>�~K,�S'J��Zb�W�r��z��w�2l���X�,�>��w!����?ɽ�T��<�G�BI�P���禼���rK�����1�
��jR������о�
�i/���U���z�fҍ� ښ��G���   �   ����w���Ԯ��תm�|�Q���2�R�Bo微����x��s(�:�Խ�Ar�$���A�Pdػ�H�l�
�U�9笽����4*�hTX��т��@��m��������?����~��J����^wk��e?�L���9۽�`���{G�\���,S����ʼ��O��6Kڽ e(�G�u����?e�f,��p0���O��k�D逿����   �   
_���[��yP���>�9e(���h���.�������D��t������)=�dȼ��t�d!���J���9b��H��hi	���>��^z��X���ߺ�S`־?s�<	���^ �����`��ܾ0���xp�����NQ�څ�c�ڽ@����R4�D�⼰f��4��r#@�� ��(��L�=�.��`?���J��L�_�%�\�<���N�\�Z��   �   ��,���)��\!�����/���ܾ5�������R���J
Ƚ~�x�����*��@ȧ�p���(�Y�l���>�	���E�����:���8־�O���+����)��,���)��_!���.2���ܾ(8���	��~�R�����Ƚشx�����*�� ħ�����|�Y�������	�=�E���l7��u4־@K��)�?���)��   �   �[ �����[��۾h���Gm��x�<Q�ʂ���ڽJ���$O4����h�����L(@�_$��r���=�r0��uB���N�O��%�P�<���N���Z�h_�D�[��|P�h�>��g(���ٝ龞1������D��v�,���\,=�|ȼ��t����h?��Z1b�C���e	��>��Xz�@U���ۺ��[־`n�$���   �   �;���鴾���̗���늾5rk��a?�����4۽f]��wG�@����Q����ʼ��Q��8Oڽ�g(�'�u������h�o.�:s0�e�O��k��ꀿI��w���/���t���ͭm��Q�2�$�r�ؼ���x�	v(��Խ�Dr�<�h�A� Oػ�H�����U�.ᬽ@����*��NX�E΂�=��{���a����   �   �z���w�Gl�{X�v�>�s!�̩��:ɽ�P����G��E������榼(��� K�@���8�
��mR�鯗���о�
�t/�h�U�u�z��Ӎ��ۚ�bI���T��(���)���!���AR|��V��!0���
��CѾ�ؖ��N�;7�5������hJ1�@B�:�t);�߮�7����3��ܒ��ӽ
:�qF,��!J��Tb���r��   �   ��!�5!�
3����J~��;ҽ5���T����5���$���xԀ�4Һ�Jlz��.ӽQ'�k�z�r����$��~�!���L��y��ӑ����G����"������v����KI���Z����y�M���!�z����۰�ŷr����R��$~,�h�:�@F�;lmb<xMF<�hB;H�F�L��"�]�����_�Ͻ ���Z�����   �   Y5Ľ�Ž[)�����ʲ��Fb��v�J�4���ʼ<~��ȭ4���E�V��Zn#�� �������@������Z̾l���07�*g�Q.��أ�_����:ɿ��ӿ��׿�Կ��ɿ1��}	��[(��(�f��-6�
�[ȾL����1�ɛϽ��H���R�H�"<�>�<��<.e�<�=< ���V�������V�}���)[������   �   �Z]�ʹc� �]��~L��z2��m�(߼0H����=�@�ۻ�/�� -&������&7�������T�$ĝ���߾�����G�9�{��u�������{ȿ=ڿ���ͪ���cڿ�ȿ�ѱ����|z�+;F�'o�&Tھ�����C�
���<`��|n�|B<8��<7
=F	=z�<�j�<P��; �ɻ�����u ��*�tJ��   �   �F��������L��̿м襼@�l�p%��҄�@�̺ 11�8�� ����D�~���ĝ�0�a�2覾H���!�B�R��t���L��l���щҿi忊�v<�����C]ҿᓺ� ���E����yP�O[��澕�QPN�@��<�o������#Q<L��<dy=�&'=��=���<�V�<X.0<  ��(�%�<3��t�Ѽ�   �   �H���ȼ��ɼ�~��t���
y�(L(�`s��@MҺ ��8��纐��@�ü�YI�?���V���Kf�������e�#�-VV�M�����������տ��V���8�����.���տ�����C��Hƅ���S��!���`Ρ��*R�h���u�P���@�U<���<�X&=��0=y�&=Mt=�<�<Z��<p��;�P��:�D1���   �   F��h��������ܾм�楼��l��"��̄�@�̺� 1������ҒD�>������a�a禾,��=!�R�R�lt���K�������ҿw忍�u;����1�j\ҿ���w��������xP��Z�����?ON�ʿ�2�o���P'Q<���<�y=�&'=&�=�<�V�<�.0< ��ж%��2��0�Ѽ�   �   �Z]�L�c�n�]�~L��y2��l��߼xE����=�p�ۻ  ���#&� ����"7�B綠\����T�����߾\���G�	�{�;t��W���zȿ@;ڿ�����1��Yaڿk�ȿб����{zz�u9F��m�#Rھ7����C�)���8`�rn��B<���<�
=�F	=,�<bk�<��;��ɻ$����u ��*�(J��   �   5Ľ��Ž�(������+����a��ցJ�V�|�ʼ�y��Т4��E�\N��\i#�7��������@�x����W̾����.7�"g��,���գ����8ɿ	�ӿ�׿Կ%�ɿ���t���&��4�f� +6�3

��ȾF���9�1�ʗϽ��H���R�x�"<^B�<b��<�f�<�=<����pU�����Z�V�`���[��䦹��   �   i�!��4!��2�����}��+:ҽ6�����z�5��򼔗���̀��䣼ƴ�Pdz�0)ӽgM'�X�z����e ����!�/�L�ly�ё�����J���������ds�����F��NX��Y�y��	M���!����<ذ���r�&��6M��~w,�(�:�0_�;�ub<�RF<�vB;ȭF������]�ث��>�Ͻ���Z�����   �   kz�j�w�	l��zX��>�s!�D���9ɽxO����G�4B�t��ܦ���K�P���.�
�(hR�1�����оi
��/���U��z��Ѝ��ؚ��E��9Q������醛�!����L|�e�V��0�h�
�)?ѾՖ��N�|3�텖�<��(61� ��: �);�Ӯ�5��L�3��ܒ��ӽ�9�_F,��!J�pTb���r��   �   �;���鴾��������늾�qk�
a?�d��j3۽�[��hsG�����,G��L|ʼ�	��K�� GڽFb(���u��~��7b⾂*��n0���O��k��瀿���ﶊ�����&�����m���Q��2�@��k�����x��p(�d�Խ,:r�,����A� 3ػ��G���ΠU��ଽ���j*��NX�<΂�=��t���W����   �   �[ �����[�u�۾:���m��8򅾨Q�$��~�ڽ�����J4�8���Z���輈@�v�����Ԅ=��+��}<��BG侩J���%�~�<�|�N��Z��_���[��vP���>��b(�d�{�龻+�������D�|q�ֵ���!=���Ǽ��t���� ;���/b��B���e	���>��Xz�8U���ۺ��[־Zn����   �   ��,���)��\!�~���/���ܾ�4��T��H�R�r���Ƚ��x�ȅ�T�����������zY�������	�$�E����.4���0־�F���&�l����(��,���)�Z!�ת��-���ܾ�1�����A�R�{���Ƚ^�x��� ��캧�����|�Y������	��E���c7��o4־=K��)�>���)��   �   	_���[��yP���>�*e(���:�龵.��̅��c�D��s�򸥽t%=�d�Ǽ��t� ���0��d(b�w=��)b	���>�bSz��Q���׺�kW־�i����`Y �b���V���۾B����i��k7Q��~���ڽ����F4�8���Z�� �輼 @��������=��-��V?���J��L�]�%�Z�<���N�[�Z��   �   ����x���Ԯ��Ъm�t�Q�{�2�A�o�{���Nx�Ns(�ӪԽB>r����A��!ػH�G�`���U�۬������*�LIX�˂��9������4���g7���崾������n芾Blk��\?�ʞ��-۽�W���mG�(����D���}ʼt��M���Jڽ�d(�$�u�	���7e�d,��p0���O��k�E逿����   �   �R��x������������O|���V��0��
��AѾ�֖�*N�B5����r��X71��ݟ:��);@���('���3��֒�l ӽ�5�lA,�J�ZNb�q�r��z���w��l�+uX��>��n!�����3ɽ'K��|�G�>��貼Xۦ���K������
��jR�筗��о�
�g/���U���z�fҍ�!ښ��G���   �   �����t������G���Y����y�lM�<�!�h����ٰ�u�r�ܫ�\O���y,���:� f�;�~b<bF< �B;x�F������]�^���ƖϽ����U������!�0!�@.�y��v���3ҽ稨������5���񼬑���ɀ�x䣼���fz�R+ӽ�N'���z�����}"����!���L�z
y�Qґ������j!���   �   X�׿mԿm�ɿ������'��Έf�n,6�8
�Ⱦ^�����1���Ͻ,�H���R�8�"<~E�<���<\n�<��=<�����E��4|���V�r����T��*���D.Ľ�Ž�"����⬙�]��>zJ�R�D�ʼ�r��ؚ4���E�tN��tj#�O��L�����@�b���Y̾[���/7��g�[-���֣�,���R9ɿT�ӿ�   �   ک�(��HbڿJ�ȿ�б�����{z�p:F��n�PSھ����C���彞:`��tn�HB<z��<��
=I	=�
�<�s�<���; �ɻ�����m ��y*��J��Q]���c�4�]�vvL�s2�g���޼�=����=���ۻ����!&� ����#7��綠�����T�8Ý���߾����G���{��t������zȿ<ڿ����   �   �;��N���\ҿ����੟�����yP�[�u�Y��ON����l�o�����&Q<>��<�z=.('=��=ڟ�<�[�<�:0<  ����%��*����Ѽp=����������طм�ॼX�l�x�п����̺@1� �����D�����'��^�a��禾���}!���R��t��/L������T�ҿ����   �   �������B���w�bϿ�䫿���M�Q�\��m׾R��!c1���ĽT�,�OɻV��<���<��<��<H�<�*&< 
����M�d���]��M�t�*���,�n#�J����� ᥼��A��]���F�:�E�;���:` �ȩ�f;�����A��V���޾����T������(���lп�3�F#��&����   �   ��t�L�����^��e'̿�,���憿'{N�iM���Ӿ9���$.�D����)���л As<e�<b��<Fg�<�C{< �;؏�8���N���p(�`D�t�R�:|T��I�fm2����l�ۼ�����
�@Vɺ@D�: ��80����鼠�{��~�I>�d���ھr@��AQ�n1���O���Ϳ�O�p��T���n��   �   v���,�^�
��B��;��!�¿�=��Tp���\D�=����Ⱦ /��B�$����~�!��8컄�:<N�<�<��D<�2>:��[�8E�H5�lcn�(���i(��6n�������h���jfr�pt@�������(D��
������09��J��n�3Oؽ�]3�]����ξ�=��F�Lm��:	��jBÿ��e0����
�@��   �   L!	�����O �����ѿK㳿7����l�&4�����
���s��A�֟��~����P��;H�<@�y;�� ���Ǽ�,4�j���W�� �սo���0���	����=�����{b̽	 ��e쁽ƛ:���� K���YU��^{�d���d[�HEĽe�"��~�ǀ�����6�V�m�����쳿�dѿ�r�> ����   �   �A��)i񿥷�Bӿ"���Qˠ�������R��D �	��l�����V�*��P��F	�pL�`C���LԻ���n��d,z����f0�?��Y,1���F�U��A[�ضX���M�~�;�{0$�L	�L�ڽf]��NCh��V��Ҽ�۳�@
뼚F� Ϋ��0� �^��¥����R� �}�R�댄��X��5^eҿ���K���   �   3�Կ\;ѿ>ǿ���h���犿��d� �4�%`	�F�Ǿl���g6����hS~����`����w��8�߼ qB�u`��j�⽊����C�_Lm��K��sK���E���L��P
���ś�V��z�#�R�r*�5���þ���`V2�H��lK ��2�ӭ����Mt;��B����Ⱦ,I	��[4�J�c�r���Z����*ƿ��п�   �   ���F_���Ӧ�7������$�g��,>���5�̹��r�c��i����EY�V����ڼ����`^�h������.3�8k��䒾����;�ɾtC޾�뾭J񾤾���hξ�������3�y�93B�7��S=˽۴���8<�����e%��<q�>t���T���c��壾Hᾅ���\<�F_e��t��T���Lӥ�\ή��   �   \	���ҍ�A҆��Pw�$�Z��(:�Ku�F��(#��Sق�=<4�������;�L��F��g�Ҡ��i&���@�����⏨��dоW\���0�G2�ac$�q�'��P%�����0/����־���䈾F�L��:�DLǽ3'���w8��[!�^�E�4���f:��1�x������v������7�8�W���t�\օ�]H���   �   K`���\��Q�J+@�z�)�"��{�aϸ�z����G����f����\i�v�(�,�$��v]����ߐ��@�Hm��/�������0���&�8�=���O�4�[��N`�s�\���Q��.@�\�)����뾊Ҹ����l�G����n����_i��(���$��q]��������?��j������e��1.���&�ج=�B�O�e�[��   �   !�'�SM%�����G*��˳־��nሾ3�L��7�8Hǽ�$���u8��[!�F�E�����>�G!1�Pz�����e��W���7���W�s�t�_؅�uJ��z���ԍ�7Ԇ�BTw�T�Z�N+:��w�����%��Dۂ��>4�6�뽯𓽤�;�����B��g�˛���"���@���2����`о4W���-�(/�`$��   �   IE�`���ᾔcξ
���������y��.B�����8˽�����4<�n���f%�$@q�jw��W�!�c�F裾��ᾠ��j_<�[be�Pv��H���dե��Ю�$��ma��֦��8��1�����g�/>�r�R8�ۻ��Q�c�vk�9����FY������ڼ@���X^������*3�<k�����ϛ���{ɾb>޾����   �   �H��=�������R���z���R�%*��������a��bQ2�����J ���2�����7���v;��D���Ⱦ�J	��]4��c�����\���𵿛,ƿ#�п\�Կv=ѿ;ǿQ��Uj���芿�d���4��a	�R�Ǿج���h6�5��dU~�V������o��(�߼
hB�wZ�������]�C��Em�H���G���A���   �   �;[�ڰX� �M�S�;��+$�H	�ހڽIX���;h�@Q���Ҽ\س�(
�^F�Ы�@2���^��ĥ�'���� �y�R� ���eZ���ﺿ%gҿ���E��C��k�u�忼Cӿ�����̠� ���@�R�F ��龵���a�V�&+��Q��x	�xL��)���$Ի4���Z��� z����(�s��'1�-�F��U��   �   ��	����U�����&\̽�����災��:���hC��HPU�@Z{� ���f[�GĽ��"�~�E������l6�
�m������3fѿZt� �ھ�""	�z��fP �U���ѿM䳿���;�l�,�4�������)�s�iB����������`��;��< )z;X� �(�Ǽ�"4������P����սe��� ��   �   �h�����9z����^r��m@�$�������C�0��� ���09��K�x�n��Pؽ�^3�,����ξu>���F��m��
��OCÿ�㿃1��`�
�����j-���
��C����ӻ¿k>���p��1]D����:�Ⱦs/����$�������!�p3컄�:<�<v�<��D<��?:�[�X6��5�Zn����,#���   �   z�R�^wT�&I�>i2����ۼ|����
� &ɺ�d�: ��8����鼬�{����>�瑓��ھ�@��BQ��1��KP��oͿ`P�������o�8 �jt����������'̿�,��#熿o{N��M�>�Ӿ`���B$.�=D����)���лpDs<^g�<���<~k�<`N{<��;h���������k(�hD��   �   ��*���,�Zn#����L���᥼�A�@`���<�:@C�;���:����뼨;��p� �A��V���޾���T������(���lп4�P#��&��������~�:���w�bϿ�䫿���%�Q�8���l׾'���b1���Ľ��,�`Lɻƺ�<��<&�<>��<~�<+&<�	����M�����]��M��   �   X�R�:wT��I� i2����`�ۼ�����
��ɺ�|�: � 9�����鼬�{�[~��>�-����ھ8@��AQ�81���O���ͿcO�2����pn����s����8��з��&̿,���憿�zN��L�F�Ӿ����R#.��B����)���л\Gs<vh�<V��<�k�<�N{<��; ����������k(�XD��   �   �h�����z�������]r��l@�P�䓴�8�C�P������9��E漘�n��Mؽ�\3�ˈ��*�ξ =�6�F��l������Aÿ��i/��:�
���ئ�6,���
�~A��>��B�¿=���o��|[D�u��_�Ⱦ&.���$�)���b�!��!�h�:<��<��<��D< �?:h�[�6켪5��Yn����#���   �   ��	����5��T�뽼[̽���U災@�:����?��GU��N{�8��`a[�DCĽ�"�2~��������6��m���y볿�cѿvq�z
 �4��t 	�����N �|�뿕�ѿ⳿4���7�l��}4����c	���}s��?�B���.�����pƭ;��< 6z;H� �h�Ǽ^"4�x����P����սR���� ��   �   w;[�°X���M�!�;��+$��G	�:�ڽ�W���9h�O�0�Ҽ8ѳ�� ��F��˫�
/���^���������� ���R�ڋ���W���캿�cҿ��\��?��1g����R@ӿ�����ɠ�Ű����R�9C ���龤����V�&(��M������K����pԻD������| z�����'�n���&1�$�F��U��   �   �H��1������gR���z���R��*�`������(��VN2�����E �x�2�ƪ��6���q;�?A��b�Ⱦ�G	��Y4��c�	��SY���쵿�(ƿ�пԿ89ѿ/ǿ�	���f��
抿�d���4�{^	���Ǿ����1d6��~�dL~�6��ĕ���i����߼�fB�"Z�����΢�N�C��Em�H���G���A���   �   CE�T����|cξ駵�j���M�y�p.B�b��J7˽����0<�"��d_%�6q�Lp��R�;�c��㣾M|ᾘ��lZ<�e\e��r��t���Bѥ�6̮����]���Ѧ�5��õ��	�g�*>�v	�(2�>�����c��f������=Y�b��p�ڼ����V^�'������)3�,k�����˛���{ɾa>޾����   �   �'�NM%����	��)*����־���:ሾ��L�7��Fǽ�"���p8��T!�t�E�8���o5齹1��u�����뾞�ց7��W��t�eԅ�JF��=��fЍ�:І��Lw���Z��%:��r�?������ւ��84���>ꓽ��;�����>�b�f������"���@�����,���|`о2W���-�(/�`$��   �   K`���\��Q�A+@�n�)���{�5ϸ�F��n�G��������Xi���(��$�&j]�	������?��g��d���I�徵+���&���=���O���[�8G`���\�l�Q��'@�f�)�x�ew��˸������G�(������Si���(�j�$�2n]���������?�j������_��0.���&�ڬ=�B�O�f�[��   �   \	���ҍ�?҆��Pw��Z��(:�<u�"���"��ق��;4�<�뽸쓽β;�>��t;�n�f�p���z���@������B\о>R��+�,��\$���'�J%����#��%��<�־D ��Rވ�<�L��3�Bǽ����m8�NT!�x�E�����d9齨1��w������l������7�8�W���t�]օ�]H���   �   ���G_���Ӧ�	7�������g��,>���Z5㾟�����c��h�W���J@Y������ڼ���NO^�ٟ��f�X%3�yk��ݒ������vɾ_9޾m���?�������^ξ����׶��a�y��)B�����1˽J��� ,<�����_%��8q��r��0T�T�c��壾<ᾂ���\<�E_e��t��U���Lӥ�^ή��   �   5�Կ^;ѿ=ǿ���h���犿��d���4�`	�$�Ǿ=����f6����pO~����䒔�xb����߼�^B��T��f��R����C��?m�vD���C���=��PD����Ž���N��0z��R�+*����Ʒ������H2�*��6D ��2�,���ݯ��s;��B����Ⱦ(I	��[4�J�c�r���Z����*ƿ��п�   �   �A��+i񿦷�Bӿ!���Pˠ�������R��D ���G���J�V��)�BO����H�K������ӻ\������z������򽼊��!1�`�F��U�B5[���X�&�M���;��&$��C	�Jyڽ�Q��1h��H���ҼT̳�8���F��̫�E0��^��¥����P� �|�R�댄��X��5_eҿ���M���   �   L!	�����O �����ѿI㳿5���ލl�4�����
���s�/A�����V��8��Pԭ;(<�z;�� ���Ǽ�4�����J��6�սH������P�	�`��!������T̽E���n⁽V�:������6��;U��G{�\��@b[�fDĽ�"��~��������6�U�m�����쳿�dѿ�r�> ����   �   v���,�`�
��B��;��#�¿�=��Rp��{\D�6��x�Ⱦ�.���$�_���z�!��!�H�:<��<��<d	E<��@:�z[�h'�@�4��Pn��������^c��+���t��뜎�RUr�~e@��	������C��յ� z��p9�PE�0�n��Nؽ`]3�P����ξ�=��F�Km��:	��kBÿ��e0����
�@��   �   ��t�L�����^��e'̿�,���憿%{N�fM���Ӿ-����#.��C����)�p�л�Hs<j�<
��<�o�<�X{<`�;�r�П��"���f(�D���R��qT��I�8d2�n��دۼ8�� �
� �Ⱥ@��: �9��8�鼼�{��~�5>�`���ھq@��AQ�n1���O���Ϳ�O�p��T���n��   �   ��E���A� ~7�R�'�ĝ��N���IԿiH���B����A�$��{J����j��
�G����ּ �z84�\<�l�<x�_<���;�@ӻx����P��6�ڳ]�ny�f����lr���T���,�L���T8���@���˺ ��: -��lp�`v$��ߨ�7��ayv��0������E�6��������տ#d ��(��(���7�J�A��   �   |$B���>�2k4�<%�\L��b���ѿq����"����>�^��U���wf�m���Z����ؼ X���7<��a<��< ���b[�8��
�+�D�`��녽����{��,白Z?���"�0S�� ��ټ�r�����@Vº��~��m���9$�j_����Qr��ʺ��z	���A������7����ҿ<�������F%�&t4�6�>��   �   fA8�85�"�+�NG������� rǿ�ğ�=�u��H5������⫾��Z��� �X���!߼`᧻ ��;`>e;`���	��>���>X��搽�!��R�̽�$߽�罥Y��=׽)��rB���:��p$B�b$�Λ�P�5�h5'��i��*=$�1Z��:�G'e����X���7�$rx�����ȿP��ּ�;�s+���4��   �   �R)���&�2)��@����޿]���l���gb�`�&�0��񆝾&aH�^�������UF���(�h�`6缼�D��L��B�Ž��������$��1�A6���3��*�'��y��ܽ�g��VWz��'+�0�� R����ɼҭ&��C���� ��VQ�V����~�Ru(��d�����ʸ�8޿�� �������A&��   �   ��R���l�v��z翛�ƿc錄͍��{I������ϾQk��1�I�Խ��o���4��� jռ�\$�����,ɼ�\� �;;%���H�j�h��\���找WM���C��N����p��bR��40����n�ս=D���V����le
���.�C��R��8��{��xҾ���?J�����¤�	aƿ1濬~�����K��   �   ���Z� ��j����ῼ�ȿ7{��o����b��#-�N~�������an��������~d�tD�0E���O��*��w
�T�PM����Pڙ�z���/�¾3�ξ�Ӿzо�žL������`�����X�0�'�����;��l�x��A���@�e����)ǽBm��-r�����,���-�{-b���Yl��e�ǿ�j࿄���u ��   �   ��ۿٗؿ\Jο
ս�����e��,n�%�<�s���Ѿv�����D�����~ a��F�D�n�Ei��Z>����.��}l����Pa\�� �O���7�.d�Z��r��J��}�\o¾K���Dw��9�b��<V��&��`�P	v�{������fF��ϒ��о���O;��l�{������:��x�̿�׿�   �   ���J�������U���-w���i�v�?��F����5"���i��g���Ͻ@/���3j�@�~�dz���d����5�U�|�䟨���׾1������2��KC���N���R�҄O��#E���4��T��V�� ݾ�����?%=�N,��!������z�u����y�нb��=}g��L��B�⾘j�=�,f������k��3K��.P���   �   @gЉ����xup���T�P5��Y����鴰��O��DF3�h��@ȧ�ٓ��#Q����}r���.���z�����>徖���.2�;�Q�P�m������<�������҉����}yp�+�T�[5�K\����췰��Q��LI3�@��Dʧ�;����O��2���m�N�.���z����@:����+2���Q�.�m�Z���i:���   �   q�R�ҀO��E��4��Q�&T�vݾ��������!=��)�^��&�����u�c�����н#��K�g��O��
��m�=��/f��↿�m���M���R���������������� y��6i�<�?�!I��徦$��M�i��i�(н0��X2j���~�Zv���^��c�5���|�:����׾t�w��:2��GC��N��   �   �`���o��G��x�k¾�G��?w�X	9�W��R���#��
`�H
v��������iF��ђ�)�о"��=R;��l�[��!��&=���̿��׿*�ۿt�ؿ�LοK׽�����g��n�r�<�6����ѾE���W�D�x����N~a���F��|n�Rd��l7��V�.�	xl�m����鼾9W�� �*���4��   �   ��ӾuоM�žꢴ�6����G�X���'�����7����x�:A���@�1���,ǽ<o��0r����0���-�0b�C���4n����ǿ�l���.w �:���� ��l���῰�ȿ�|��ՠ��V�b�L%-�܀���ñ�Gdn�a��	���~d��A�&@��O�%��8ή�RJM�����R֙� ���Q�¾�ξ�   �   �I��@��� ���p��\R�00������սR?��ҞV�2���b
�l�.�D����̥8� }��%zҾ}���AJ�ĵ��}ä��bƿ%�������M�������m�v�G|��ƿ��Ύ���|I�����Ͼcl���1���Խ��o�`��܇��h^ռ:T$����6¼�� �#6%��H���h�)Y�� ㉾�   �   6�g�3���)����u���۽b��TNz�� +�H�㼠K����ɼ��&��D���� �\XQ�����a�v(�3d����0̸��޿�� ��������B&��S)���&�$*��A�i��޿^��jm��4ib�P�&����·��5bH�r��V���hKF�0����h��&�ތD��F��$�Ž����t����$�X1��   �   =�FS��7׽�#���=��K6��hB����ś� �5��-'�Hh���=$�[���:��(e������Y���7�gsx������ȿg��v���;��s+���4�6B8��5�ԝ+��G���h���rǿ5ş��u�CI5�ݧ��㫾��Z�� �z��  ߼ ӧ�0��;�{e;P镻 �������5X��ᐽ���$�̽U߽�   �   x��+䙽�<�����S�� �(ټ��r����+º��~�tm��T:$�`�����-r�}˺�e{	�$�A�����e8����ҿۨ��R��PG%��t4���>��$B��>��k4��%��L��b���ѿ�����"��ި>��������wf�����Z����ؼ@:���7<L�a<��<���S[�t���+���`�
酽�����   �   z�	Á�mr���T���,�ܹ��9���A� �˺���:�6�(np��v$�N਽p���yv��0�����'E�O��������տ1d ��(��(���7�P�A���E�|�A�~7�D�'����rN��rIԿMH���B����A���DJ��F�j�F
��F���ּ �{8�\<�l�<�_<���;�?ӻP���~P��6��]��y��   �   �w��!䙽v<��g�`S��� ��ټH�r��鿻�º�s~�<k���8$��^������r��ʺ��z	�F�A�g����7����ҿѧ������F%��s4�Ύ>�
$B�H�>��j4��%�L��a���ѿ����6"���>�������vf�����Y����ؼ@���
7<رa<��<���S[�\���+���`�
酽�����   �   6�6S佷7׽l#��V=��6���B�
��Û���5��''�d���:$��X��X9�M&e���SX�6�7�>qx�C���V~ȿm��N��f:�Xr+��4��@8�l5�`�+��F������7qǿ�ß��u��G5������᫾u�Z��� �����߼�ŧ�ઇ;��e;�啻����h���5X��ᐽ���&�̽N߽�   �   �6�Z�3���)����u���۽�a��PMz��+���TG����ɼ֩&��A��|� �(UQ�O���}�St(�6d�����ɸ��޿�� �0�����v@&��Q)��&�2(��?���(޿�[���k��Ofb��&�R�꾔���(_H�X����x� BF�(��ؖh��%缈�D��F���Ž����r����$�T1��   �   �I��@��� ���p��\R��/0����h�ս�>���V����d_
�x�.�h@��X���8�?z��>vҾ���*>J���������}_ƿf}濨}�d���J�H���hk�b��x���ƿ������yI�s����Ͼ�i��k�1���ԽX�o���@����Zռ&S$�����¼�� �6%���H���h�)Y�� ㉾�   �   ��ӾuоB�žڢ�� ������X���'�,����5��*�x�`A��@�?���[&ǽk��*r����K*���-�-+b�A󍿦j��m�ǿth����t ����� �h����ῢ�ȿ^y��ܝ����b��!-�2{�������^n�h������wd�*=�=���O��$���Ὓ�BJM�����Q֙�����P�¾�ξ�   �   �`���o��G��x�k¾yG���>w��9�����P���!��~`�<v��������cF��͒�`�оF��HM;��l�����	���8���̿p�׿��ۿ7�ؿ�Gο�ҽ�율�d���n���<�f����Ѿ$�����D�o���ꢽ�va���F��yn�Xc���6��,�.��wl�g����鼾9W�� �+���4��   �   q�R�рO��E��4��Q�T�Wݾe�����!=�)�|��|�����u��{����нo��Uyg�"J�����Xh�A=��(f��ކ��i���H���M����������.����u��@i�l�?�uD����A��x�i�0d�l�Ͻ�*��4+j��~��t���]���5���|�.����׾t�w��;2��GC���N��   �   AfЉ����rup���T�F5��Y�ߥ龾����O���E3�����ŧ�H����K������ h��.���z�u��26�^���(2���Q�/�m�,���8���닿Ή�\
��Jqp�֠T�
5�W����n���M��2B3���.ç�[����L�� ��Pl���.�k�z����8:����+2���Q�0�m�\���k:���   �   ���K�������R���)w���i�l�?��F�n��"��c�i��f���Ͻ,���*j�L�~�Zq���X��>5�B�|�����׾�|�i���2�DC��N�Z�R��|O�E�|�4��N�XQ��ݾ��������=�$&����h�����u��|����нΈ��|g��L��4�⾔j�=�
,f������k��5K��/P���   �   ��ۿۗؿ[Jοս�����e��"n��<�e���ѾA���`�D������뢽Twa��F�tn��^��w0����.�Wrl�崘��弾;R� ���Y1�{]���ll��D��s徊f¾�C���8w�`9�o���K�����|`�v����,�xfF��ϒ��о���O;��l�z������:��z�̿
�׿�   �   ���\� ��j����Ώ�ȿ5{��k����b��#-�2~������qan�>������xd��;��8�zO�v����:��DM�V~��rҙ�������¾��ξ��Ӿ�oоY�žS�������D�X���'�����0����x��A��@�y����'ǽ�l�A-r�|���,���-�{-b���[l��f�ǿ�j࿆���u ��   �   ��T���l�v��z翙�ƿ`錄ɍ���zI������Ͼ!k��6�1���Խ��o�8��T|���Pռ�K$�����h����� �,1%�?�H�T�h��U��@߉��E��F<��!���U�p��VR��*0�Z��|�ս09���V���\
�2�.��@����o�8�g{���wҾ���?J�����¤�
aƿ2濬~�����K��   �   �R)���&�2)��@����޿]���l���gb�X�&���φ���`H�6��t���8:F����P�h���&�D��@��$}Ž��������$�$1��6��3���)����q�{�۽�[���Cz��+����l?���ɼ�&�:B��� �XVQ�A���|~�Qu(��d�����ʸ�7޿�� �������A&��   �   fA8�<5�"�+�PG�������rǿ�ğ�9�u��H5����v⫾��Z�V� �<��߼�������; �e;p��������,X��ܐ�5����̽�߽�罠L�n1׽���8��x1��B�������h�5�@'��`��:$�*Y���9�'e����X���7�$rx�����ȿQ��ּ�;�s+���4��   �   ~$B���>�4k4�<%�\L��b���ѿq����"����>�[��J���wf�B��*Z����ؼ@���7<(�a<��<�G�8E[���(�+�<�`�慽|����t������b9����(S�� ��ټH�r��Կ����� ]~�pi��R8$��^�����<r��ʺ��z	���A������7����ҿ;�������F%�(t4�6�>��   �   r��m��_�hWJ�Z�1��'�x����˿ѝ���j�:�&���⾔z��{,2��Vƽvo=�DU��  !��; ��8�j�,M����THW����2��:���W����� �������p��C8�������������������ɼp`a��ؽ�";�A4��0��4�)��n�)ȟ�@�Ϳ(%���$���2���J�X8_��%m��   �   �dm�:�h���Z���F��/����P���rȿ�O����f��	$���޾����R/�{�ý�6>��苼��5� �g90���脼h���,�A��/���7��%^��*�Ƚ,OϽ$̽�\���B���ߎ�$�_����˼�g�`���A�,aԼ�~a�\Iս�
8����������&��j��#���iʿ������/��%G�[�r�h��   �   J`���[�^O�>�<���&����9��nD��[����[�����Ӿ�ӈ��$'��T���NA�����/1�@C>�,��j�"|d�;6��8�ǽ���%�Q�t��1�&�	�H���Խ�2���Â��w8�P"�������ԟ�4@���b�Ĉͽ]//�����@	ؾ\��P^��u��ۼ���*�Bo�Z�&�t�<��#O�8�[��   �   p^L��H�H>���-�����E��ܿ�ǰ�S��FJ��;�I@¾C�{�\����
�H����C˼a�L�F�␒�z�ʽC��� ��;��4P�|0^�i�c�F7`��T���@�`'���
��6۽"Σ�pfi���%����d��Xg�zl½��!��C���ž`�L�}q��2�����ܿ*O�|��\K-��y=�`H��   �   �4�� 2��
)� 1���	��R�3Uſ���qs���3��A���^��|�_����x!����X��/*��:���~�)��,����'�R�� |�����q(���"������@I���W�����Բ���Z��{/�,����ƽ�i���Y�|�F�@s��l��Fu�je�F����\ ���4�FIt�J���ſ-���H	�`a�TD(��1��   �   �����C���a���4οF!��2���m�Q��Y�Gھ�򓾧�A�z�������G�t�71q�2����hӽ���BbG�r�(���뽾�پ�������.�[���S�:�ܾ� ¾���S����O����#⽖<��Uք�i��R��U< �;iE�󇕾�;۾ ��գQ��U��<Y���̿"�����e�F"��   �   ���z�M�����5�ɿ�6��R��Td��Y.�����=�����u�[C#�~dڽ�ʟ���������7��] ��p]�b������O�4/	��*��O+��65���8��6���,��D�1��L�� d��㻗���d�/�&�2�ｳ������?���N�߽^I%�� w������Y��N�-�y�b��0��4���|�ǿ��lK��ʓ ��   �   2iտ?Nҿ[_ȿnq��sޣ��X��Fmg��x7�z����̾Ӑ��BF����½ݣ�~����a潓-"���d�1����ϾK�ć!��2>���W�� l��by�"T~��wz�}n��[Z�`�@��C$���K�Ӿ���Ïj��&���5��\ڧ�E`Ľ�`�}�E�����,˾X�
�2�5���d�)����	��ן����ƿ�wѿ�   �   �𧿀s���{��s���=����Z��3�� �m�׾G�v�_��f�Tbݽ�ݰ� ����ڽ*��<\�������Ծ���Q1��W�T:}��)��~B���Ǥ���7v��6~��ӷ��$?��F�Z��3�Z#��׾����#�_��h��dݽް������ڽ='�P8\�������Ծ�PN1�H�W��5}�1'���?���Ĥ��   �   LO~��rz��n��WZ���@�t@$�N��6�Ӿ���B�j��&�B���3��`ڧ�)bĽ�b���E�*���k/˾��
��5�-�d�D���G��������ƿ�zѿ4lտ3Qҿ'bȿt���ࣿ�Z���pg��{7�~����̾ᒐ��DF�d��½Lܣ�ё��]�*"���d�����H�Ͼ��~�!��.>�T�W�ll�^y��   �   ��8��6�>�,�tA�0��.���_��������d���&�.�ｬ������������߽�K%�c$w�,����]����-���b��2��h�����ǿџ�iN��Z� �V���7�����⿒�ɿ�8���S��d��[.����k�����u�E#��eڽ8ʟ�����3���,2��Y �k]��{��=�����,	�d'��K+��25��   �   �+��T���M��ܾ3������P���O�ʚ�Z⽸8��Ԅ�^h���R���= ��kE�ǉ��z>۾ٲ�F�Q�9W��[��2�̿���X���f��#���@��JE�4������6ο�"��������Q�[�nھR���[�A����萢�u�t�j+q������bӽ����\G����?潾)پɹ������   �   ���D���S�����j���Z��v/�Q���ƽ�e���Y�f�F��?s� n���v�]le�����] ���4��Kt��K��b ſ3���I	��b��E(�p�1���4�62�J)�X2���	�dT�VſC���ss��3��C��2`���_�Ź��!����X��+*�:�:��~�#�������'���Q��|�����'$��r���   �   $�c�"1`� T�8�@�T['�x�
��/۽�ȣ�.^i���%�����b��Xg��m½��!��D����ž|��L�xr��j����ܿP�����L-��z=�paH��_L�l�H�|>���-�r���F�#!ܿ�Ȱ����cJ��<�SA¾��{������H�����9˼4Z� �F����\�ʽ�>�̟ �;�/P�N*^��   �   .p��-���	�����yԽ�-�������p8�����y��@П�0>��X�b�ƉͽY0/�U���t
ؾ�\��Q^�yv��ǽ���+��o��&�X�<��$O�J�[�\`���[��^O� �<�.�&�F����E�������[�}��ϜӾRԈ�%'�
U��NA�����"1��1>�h����b�sd��0���ǽ��P"�IM��   �   �KϽx ̽XY��d?��(ݎ�f�_�����˼��f����0�A��`Լ6a�Jսr8�������V�&��j�7$��Mjʿ&��z����/��&G��[��h�|em�ĕh�4�Z�2�F�$	/�,�����1sȿP���f��	$���޾����4R/�p�ý6>�|拼��5� �i90��4ᄼx�����A��,��G4���Z����Ƚ�   �   �W��%��������ދp�D8�d���������0�������ɼaa�+ؽ�";�q4��p��]�)�"n�Fȟ�`�ͿI%���$�ʭ2���J�b8_��%m�r��m��_�XWJ�H�1��'�V����˿ѝ�h�j��&����fz��7,2�bVƽo=��T�� � ���; �8j��L����<HW����2��>���   �   �KϽw ̽PY��W?��ݎ�2�_����D�˼ �f�����A�`^Լ�}a��Hս~
8�b�����㾖�&��j��#��viʿ��ڣ�6�/��%G��[��h�Ldm���h�.�Z�P�F�h/�������drȿnO���f��$���޾"���JQ/�=�ýt4>��䋼��5� "j9�������`�����A��,��I4���Z����Ƚ�   �   .p��-���	�����yԽV-��P���Np8����pw��,͟��9���b�V�ͽ�./�����vؾ�[��O^�4u��-����)￼n���&���<��"O�2�[�6`���[�]O�`�<�ҹ&�$��)��C��� ��ל[� ���Ӿӈ�H#'��R��KA�����1�P.>�����Rb��rd��0���ǽ��R"�JM��   �   $�c�1`��T�(�@�=['�Z�
��/۽Xȣ�]i��%�����_�TTg�>j½M�!��B����ž���L��p��2���[�ܿjN����LJ-�tx=��^H�
]L���H�>���-���� E��ܿxư�_~���J��:��>¾��{��������H�D��6˼:Y���F�슒�D�ʽ�>�˟ �;�/P�P*^��   �   ���D���S�����\����
Z��v/���`�ƽ�d��dY���F�*:s��i���s��ge������[ �T�4�ZGt��H��%ſ[�쿰G	�&`��B(�d�1�z�4�.�1�z	)��/���	��P�Sſ����os�Դ3�[?��]����_��������X��(*�N�:�֭~��"�������'���Q��|�����)$��v���   �   �+��T���M��ܾ$������P��=�O�s��b�T7��҄�`e���N��Z: ��fE�D���z9۾f����Q�TT���W���̿������c�� �~���TB�������2οn�������Q��W��ھ�𓾭�A�����������t��'q������aӽ}���\G�����>潾,پ͹������   �   ��8��6�<�,�pA�)�����_��q���a�d��&�ʷ､�����B����߽�F%�Tw�+����V��"�-���b�=/��)����ǿd�࿇H��A� �.����N����⿯�ɿ�4��4P��?d�$W.�;���~�����u�H@#�u_ڽ�ş�򦐽v���1�pY ��j]��{��8�����,	�g'��K+��25��   �   NO~��rz��n��WZ���@�k@$�A���Ӿل��͊j�Z�&�P���0��֧��[Ľ9^��E�s����(˾E�
���5�L�d�.������I���#�ƿ�tѿ/fտCKҿz\ȿ�n��ܣ�vV���ig�v7�*��E�̾7���%>F��
�� ½0أ�(���e[潀)"���d�����?�Ͼ��~�!��.>�V�W�ol�!^y��   �   �𧿁s���{��q���=����Z���3�� �H�׾��_��e��_ݽ�ٰ�+�����ڽ$�4\�����5�Ծ��NK1���W��1}��$��P=��1¤��p���x�������:����Z���3�Q�H�׾ ��_��b��\ݽlذ�����6�ڽ{&��7\�c�����Ծ�QN1�I�W��5}�3'���?���Ĥ��   �   2iտ@NҿZ_ȿlq��oޣ��X��=mg��x7�j����̾����MAF���4½ أ����RW�O&"��d�����(�Ͼ��b�!�+>�:�W��l�dYy�vJ~�!nz�an�tSZ���@�=$������Ӿw���΅j���&����l.��kէ� ]Ľ�_�ڢE������+˾R�
�0�5���d�)����	��ڟ����ƿ�wѿ�   �   ���|�M�����2�ɿ�6��R��Jd��Y.��������D�u�eB#��aڽCƟ�����<����+佯U ��e]�wx�������")	�$�#H+��.5���8��6�q�,��=�
�����a[��ⴗ���d���&����{����������߽�H%�R w�l����Y��K�-�x�b��0��6���}�ǿ��oK��˓ ��   �   �����C���_���4οC!��/���d�Q�uY� ھ���A�&���g���>�t� #q�����\ӽ���wWG��뀾����὾�پ
�������(��N�� H�x�ܾN������M����O�)����2��Pτ�d���N��:; ��hE����;۾���գQ��U��=Y���̿%�����e�F"��   �   �4�� 2��
)�1���	��R�2Uſ���qs���3��A���^����_�������X�"%*�F�:���~��������'��Q��|�����������hﭾ=@��1O������˫���Z��q/������ƽ�_���Y���F�z8s�Xj��rt��ie�$����\ ���4�GIt�J���ſ.���H	�ba�XD(��1��   �   r^L��H�H>���-�����E��ܿ�ǰ�R��@J��;�(@¾݋{�����r�H����\.˼�R�F�v���|�ʽ�:�� ��;�@)P�$$^�֥c��*`��T��z@�MV'��
�}(۽�£��Si�6�%����\�DSg��j½�!��C����ž[� L�}q��3�����ܿ*O�~��\K-��y=�`H��   �   J`���[�^O�@�<���&����9��mD��Z����[����
�Ӿ�ӈ�1$'��S��TKA�`���1��>��^[�jjd��+��+�ǽj���rI�@l��)�ͽ	������sԽ�'��º���h8��
��xn���Ɵ��5��Z�b���ͽ //�m���3	ؾ\��P^��u��ۼ���*�Do�X�&�t�<��#O�:�[��   �   �dm�:�h���Z���F��/����O���rȿ�O����f��	$���޾�����Q/���ý�4>��㋼��5� �k90Xڄ�<���
�A�*��1��(W���Ƚ�GϽ�̽�U���;��ڎ�܆_�L����˼��f�@��@{A�0\Լ�|a��Hս�
8����������&��j��#���iʿ�������/��%G�
[�r�h��   �   �v��q+�������n���O�j=0����=�p඿����sC����o��%TX�CT��<6��T��� SR���(�L�,���N����`��=������d"ɽ�?ٽR�߽{�۽7�ͽd���窚��t�2�1���ز���#_�����m��������_��W�����5RF�2j�������n�0��o1���P��so����0���   �   �X���-��<���_j��:L�g-����Im�>���s��P7@��]�������T�Ą���������,��HK�|��������4B������tͽ�;轃���	p �����v1�&lԽ�����y��FbW����L�ü$	��(������"���P�ǚ[�XN��K���B�+��������鿴���m.�:�L�f�j��F���'���   �   Ҕ���~\u�P�]�:�A��<%�D&	���ܿ����<��Z�6�<���`(��boK�"�������l�ʼ4�Ҽ\��6�\��ꚽ�v˽�G��:�$E$�ߍ/��3���0���&�����/�ĭս�Х���r�~+�h����Z���,�(��� ���Q�厦�����"9��e��>8��|�޿��	�`�%��7B�Ԏ]�Nu�y����   �   �xq���l�p_��J�Vc2�H�������h̿������k��(�*|�V@��c�<��y彃��r�:���%���G��8��Z�������"���C�*�a�;�y������������X�|�o�e�1�H�u�'�Ӭ�<�˽����]�*0;��~O��"��U�ｱ4B���6�辻�)��m����sOͿ�������2��J��b^�Sl��   �   l�S�L�O���D�@�3�$I������} ��:����R�%c�@�˾�,���\+�"�ٽ�y��/�r�悽�ܩ�ċ�}��WK�س|�L���7J��׫��ɾ�S;�ʾX���ή�y���x����Q���"�������ꌽd����g��+S�Ȧ/�V\���?ξU���*S�
��&Q���㿼j����
�2�f�C��NO��   �   ��4�:2�:*)�j�d4
������ſ驞��yt�9�4�BT ������i�����^н�ᢽm&���Ž��5� �p�C��ߤ���z�����q]�҅����
)�̋��r�,侚J��L����w�=�:���	�8Eν�p���b���=׽Q��k�f䰾�� �>5��ft�#K��+ſ|��2	��B��(�(b1��   �   ����\�������Fȿ�3��|���I�K�L.��'վu��E���3{̽ۖ���R׽(���NC��섾�|��F߾���E !�l�6��aH���S�f�W�v�T��I�s�8�vU#���
��F㾺���⇾BH��"��E޽�r��kiѽ�	��2G������>վ����J�T�����	�ƿ�濞��D���Q��   �   �'��B��b=�տv����Ǣ����g$V�#�#����,:���{m��$���kнr`߽���!�D������\��g��y<��F=�C^���{��k��)���œ�=����p���1~��a�Y�?�������P��/H���rH�zf�"`㽸Cӽ^P��%��m�2���:�ﾻ�"�!OT��N�����6����ӿK��ަ��   �   ~G¿�m���U�������~�]�Q�$]&�����9���4��L�;�x�*<޽`�ݽш��:��΃�;�������Wr$�rO���{��@��W��^��ٲ���J¿�p���X���ç�}��~���Q��_&�ϰ��N���V!���;�ry��<޽ؠݽ��a	:�t̃�Ƌ��#���Wo$�UnO�6�{�=>�����b�������   �   P�����n���,~�� a���?� ��Z���BM���E��]oH�<d��]㽲Cӽ~R��S%��m�����$��Y�"�zRT��P��$�������ӿ���H��D+�����@�	տ����ɢ�����r'V�z�#����<���~m���$�C��jнf]߽��	�D������X��S��Q9�C=��>^���{�Gi��m����   �   ��W��T���I���8��Q#���
��A�����$߇��=H� �dB޽q���iѽ3�	�O5G������Aվ)����J�������ƿ��6������S��������������rHȿ�5�������K�0�	*վ�v����E�؞��z̽����tN׽����IC��鄾�x���@߾x���!�l�6�a]H��S��   �   #���%�s��wo����E�������w���:�2�	��@ν*n���a���>׽����k��氾M� �_5��it��L��Hſ�~�J4	�fD�j!(�d1���4�2��+)��k��5
����ſp��� |t���4��U �M����i�����^нLࢽ&#��� Žd��*�4���p�P�����uྵ���Z�E���   �   aN;�ʾm����ɮ�u��Du���Q�q�"�:��(���X猽����Ng��dT�G�/��]���Aξ̊��,S�V���R�����k�����2�0�C��PO�b�S�.�O�L�D���3�bJ��������!��K����R�Gd���˾�-���]+�r�ٽ~x��b�r�8₽ש�k��ƶ�3QK�ج|�:����E��ݦ���ɾ�   �   ���~����|�E�e���H�ƌ'����˽;����]��+;�p|O��"�����6B�2������)���m�!����PͿ��������2�PJ�*d^��Tl�dzq���l��_�L�J�dd2� �������i̿�����k��(�d}�A��$�<��y�����:��%��G��3����������"�~C��a�j�y������   �   ��3���0���&���I,��ս�˥���r�x+�ؘ���U����,�^�����
�Q�ҏ��p����#9��f��9����޿T�	�(�%��8B���]��u�,����������]u�H�]���A��=%��&	���ܿ���������6�����(���oK�^��"�����<�ʼ �Ҽ����|\��嚽�p˽�@��T��@$�t�/��   �   �m �g|���-�hԽ΄���v���]W�\���üH�� ���z��]"��^Q���[��N�������B����l���E����n.���L��j��F��'(��OY���-���<��`j�*;L�\g-�ī��m�z��t���7@�^�	�����T������������()�� K�Ђ��X����/B���� �[pͽ�7�L����   �   \�߽��۽W�ͽ~������t���1���뼐���H%_����`n�����<��2 _�X����eRF�Pj�������n��0�p1���P��so����!0���v��l+�������n�j�O�T=0�����P඿�����sC�����n���SX��S���5��|����QR���H�L���������`�l=������]"ɽ�?ٽ�   �   �m �k|���-�hԽ�����v���]W�$���ü0��\���@��q!���P�t�[�N��"����B��������O��|��Xm.���L���j�=F��e'���X��?-��!<���^j�B:L��f-�2���l�����s���6@�]�B�����T�X���ڍ��x���'��8K�X�������/B�����^pͽ�7�V����   �   ��3���0���&����@,�ѧս�˥�L�r�lw+�����`R����,����������Q�B���$���"9��e���7����޿2�	���%�"7B�ҍ]�u�̡�����X���6[u�6�]�N�A�8<%��%	���ܿ#������`�6�Ҷ��^'���mK�Ȥ�u��v����ʼx�Ҽ<��~|\��嚽�p˽�@��W��@$�x�/��   �   ����~����|�;�e���H���'�Ψ���˽������]�|);�2yO�@ ��ڠ�93B�
��ԣ���)���m� ���RNͿ���ڲ��2��J��`^�HQl��vq��l��_���J�&b2�J������og̿�����k��(�Qz�?��c�<�Ev�~�� �:�D�%���G�x3����������"�~C��a�p�y������   �   gN;�ʾl���~ɮ�u��8u���Q�=�"����N���挽����Zd���O��/�[���=ξ��K)S�����O��\�㿰i�R����2���C��LO�x�S�b�O���D���3��G�|��%�����򘍿�R��a��˾J+��yZ+�&�ٽ�u��Ղr�%Ⴝx֩��轮��*QK�Ԭ|�=����E��㦽��ɾ�   �   %���%�s��to����E��o����w�Z�:���	�X?ν
l���^���9׽�2�k�{ⰾj� �f5�^dt��I��Cſ�y쿄1	�<A��(�J`1��4�T 2�n()�nh��2
�a���ſ.����vt��4��R �Y���8 i�U���Yн@ݢ�8!��X�Ľ
����4���p�I�����uྼ���Z�I���   �   ��W��T���I���8��Q#���
��A������އ�G=H�P�8@޽:n���dѽz�	��/G������;վ,��{�J�����������ƿU�������P�2�������^��6�迚Cȿ�1������}�K�*,�V$վ�r��H�E�8��v̽�����L׽A���IC�z鄾�x���@߾w���!�o�6�f]H��S��   �   Q�����n���,~�� a���?���>���M��XE���nH�4c��Z��>ӽbK��%� m��~���~�X�"�LT��L��{�������ӿ�必��`$��ו�:�տ����)Ţ� ���!V�z�#�~��.7��Pwm���$�S��
fнrZ߽��{�D������X��J��P9�C=��>^���{�Ii��p����   �   �G¿�m���U��
�����~�S�Q�]&�u���������^�;��v��7޽�ݽ���:�ʃ����������l$��jO��{��;�����x�������ZD¿�j���R��=����딿v�~���Q�Z&�Ч���~��|��/�;��t�p6޽��ݽ����:�6̃��������Uo$�VnO�8�{�?>�����e�������   �   �'��D��b=�տs����Ǣ����^$V��#�]���9���zm���$�N���eн#X߽ɴ���D�����T�����W6�k?=��:^���{��f���󐿌���ȃ��ok���'~�6�`���?��|�%���-I��rB���jH��`��W�.>ӽ�L���%�Em����� �ﾶ�"�!OT��N�����9����ӿN�����   �   
����^�������Fȿ�3��x���>�K�<.�M'վ�t����E�s��xv̽쏻��H׽P��=EC��愾�t��<߾���?!���6�"YH���S�4�W�e�T�j�I�v�8�YN#���
�}<㾢��ۇ��8H��<޽l���dѽ]�	��1G�Z���l>վ����J�U������ƿ	�濠��F���Q��   �   ��4�<2�8*)�j�d4
������ſ穞��yt�-�4�.T �g����i�����ZнPܢ������Ľ���g�4���p���������oྤ����V��~�����!�	��Nl� ��A��p���5w�h�:��	�7:ν�h��6]��:׽�G�k�1䰾�� �:5��ft�$K��+ſ|��2	��B��(�*b1��   �   n�S�N�O���D�>�3�$I������{ ��7����R�c��˾�,���[+�9�ٽBu��r��݂�oѩ�8}�<���KK��|�H���.A�������ɾI;wʾh~���Į��p���q����Q�{�"�>��̉��8⌽D���Xc��NP�ܥ/�\���?ξM���*S�
��(Q���㿾j����
�2�h�C��NO��   �   �xq���l�r_��J�Vc2�H�������h̿������k��(�|�!@����<�kw�l����:���%���G��.��V�������d�!��xC���a���y�f���c����z����|���e���H�ć'������˽x�����]��#;��uO����D��	4B�����辷�)��m����uOͿ�������2��J��b^�Sl��   �   Ӕ���~\u�P�]�8�A��<%�D&	���ܿ󫫿:��T�6�*���@(���nK�ҥ���,����ʼ��Ҽ.���t\������j˽ :�����<$��/��3��0�z�&�	���(���սkƥ���r��p+�����K��H�,�'��4���}�Q�Ȏ�������"9��e��?8��}�޿��	�`�%��7B�Ԏ]�Pu�y����   �   �X���-��<���_j��:L�g-����Im�>���s��O7@��]�ч����T�"��������h%�� �J��|������+B�V����쫽�lͽ�3�"����k �"x��j)�dԽF����s��^XW�̐�<�ü����|������!���P���[�JN��I���B�,��������鿶���m.�8�L�f�j��F���'���   �   yZ���U��I���L��&nl�<xF��A#��>���̿������\� ��Ǿg�y���1ߦ���0��ü��������*�P�S��
����5սW���t ����jX�d����ٽ?����N����`����$qܼP����6�0�?�<���>:�s�~��4ʾ�y�@_�"��|�ο�m�Ό$�|�G�fsm���������[���   �   匥��������������h�^C�� �l;��xɿ�����X������þf"v�NK��1���7��5޼�ʿ�$�����2�5}�����r�нD���	���P4���`�
�|����Kֽ�/��\��\�@������ۼ�^���`F��׮�
���{�
�ƾ��fU[� ���T˿nO�0�!��-D���h����~���i����   �   �Ś��F�� F���=}��[��9��@�����5���ꏿ�bN����F^���Zk����$���f�M�\��$����K�dO���z�� ��RK�W�+��>�i�J���O�VL���@��.��{�?���W�Ž쑔��Z��)�6j%���[���������o����+N�5pP��*��v���Y�����:���[��*}�T���#���   �   �݊�1����~�X�e���H�t�*�.���[�O���b���7�=�"C��ҫ�c�Z�Lv�`Ȭ��u��*^�7����>�����6��=�%b����s������暾�R��4��DU����e�>A��9�،｝���?����k��/������D�<�^����z���q?����"���I;�D���*���H��Xe�p6~�ಇ��   �   ��p��Zl���^��J�y2�����?����̿�ٞ���l���(���羝����,G���ܿ������bȣ��Ͻ�T
��P7�r7k����*���Qľ��׾j?�
����+پ�Wƾ�e��������o�s�;�FH��=ֽa���$��V���0��zVJ�gl��4�龁�)���m��A��~�̿����c�r�1�N�I�l�]�R�k��   �   ��K��cH���=�\�-�:P����E	ݿ����V����K�*O���Ǿ�҅��U2�>����WƽĮĽ���o���KR��j���-����׾�������M��
�'��'+��e(���n;�7� �;�ھ��t݌�2�V��& �C�IFʽp˽|Y����4�?���p�Ⱦ���"L��M���M���6ܿ��M���,�~�<�p�G��   �   �)�~&��k����h���߿4깿�ꔿINe���)���h#����c������r:�:' �lx&�\b��w���$Ⱦ�������%6��|N�^�a��Pn��r��o�,c��BP��8�	��f} �0�ʾ����e��l)�ɑ�F��&��(N ��e�����2��e)�Ğd�=���ɸ���ݿ�� ����|o���%��   �   �V	�zR�� ����ӿ���%�p��8��R���¾ ����>�������9���&��c�O᜾�6Ծ���/��U��Gz�g��>��q���ؙ�����/��������|��W���1�z��p�־����(f���(�(��Z����@��)?�qӇ�E¾����7��!o�����M���ѿ��뿖& �����   �   %ٿu�տո˿��������񎿉l�/�;�r]�o�Ӿ闾�0X�N)��������+�V�(喾VҾ�0���9��i������2�����xʿGտ�
ٿ��տ�˿�����¦�E�dl�G�;��_��Ӿ{뗾�3X��*�5�����}���V�m▾xҾ,.�9�9���i�����/������uʿ�տ�   �   ǖ�����1,������|���W�c�1�ғ�e�־����f�2�(���E����A�$,?��Շ�a¾��٠7�:%o����������ѿ��h( �t���X	�\T��� �U��˽ӿ[��/𖿊�p���8��T�F�¾�����>�(�����8���&�O{c�ޜ��2Ծ����/���U��Bz�Td��;��k����   �   ��r��o�?'c�$>P��8�����z ���ʾŻ��*�e��i)�ԏ�qD彊'���O ��e�󍧾����g)�ߡd�?��4̸�S�ݿ�� ����tq���%��)��&��m���������߿[칿P씿Qe���)����E%����c����ʲ��7��$ ��t&��a�
t��F Ⱦ&���v���!6�bxN���a��Kn��   �   �#+��a(�W�� 8�1� ��ھT鲾ڌ��V�)# �@ �hCʽ�o˽�Z��T�4�������Ⱦ���|$L�yO���O���8ܿr�(O�`�,���<���G�2�K� fH���=�"�-��Q�޸�[ݿɨ��X����K��P���Ǿ�Ӆ��V2�Z����Uƽ(�Ľج�`|�FR� g��0)����׾����l������'��   �   ��後%پ�RƾMa���}��s�o�|�;�|D�8ֽr]���"������ڷ�$XJ��m��y��&�)��m�C��L�̿���d��1�0�I���]���k��p�]l���^�ޚJ��z2���xA��|�̿�ڞ�g�l���(���羨����-G�������0�"ģ�uϽrP
��K7��0k��������Lľ�׾�9��   �   �⚾�N��X0���Q����e��@�N5���T���f	���k�Z.��䂳�����^�C��y��=s?�����a����<�8	���*�p�H�@Ze�v8~������ފ�B��d�~���e���H�n�*����\�C������>�=��C�]ӫ�B�Z��v��Ǭ��u��$^���:9��'�罎1�x=��b������ ������   �   ��O�oL��@�Ǒ.�0x�������Ž�����Z�B�)�<g%�d�[��������o�����N�OqP��+��g���DZ��r��:��[�,}�#���$��qƚ�G���F���>}��[�>�9�8A�����16��d돿WcN�h���^��9[k���������M�d�����L�K��J�� u��7��kG���+�5�>�{�J��   �   �1����1�
�|���2Hֽy,��zY��d�@������ۼd\��V`F��׮�����{���ƾ���V[������T˿�O���!�r.D���h�m�������椡�_�������������Bh��C�>� ��;��xɿ�����X������þ�"v�EK�@1����7��1޼$ſ��z���2��}�V����}н���	�����   �   ���oX�|����ٽ`���O����`����qܼ���\7�Đ?�����:���~�:5ʾ�y�v_�?"����ο�m��$���G��sm���������[��yZ���U��@���L��nl�$xF��A#��>���̿u���z�\��~��Ǿ�y�����ަ�Z�0�4�üP���������S��
�����5սP���t ��   �   �1����3�
�x���.Hֽm,��iY��,�@����l�ۼ�Z��_F��֮�����{���ƾ��� U[�픘��S˿>O���!��-D�|�h������������k���%���"���P���(h��C��� �;�xɿ=���X�J���þa!v��J�L0��d�7��/޼@Ŀ�0z����2��}�V����}н ���	�����   �   ��O�sL��@�ő.�*x�����ϰŽ`���6Z�0�)��e%��[�*���4����o�����M�oP�o*��ϫ��?X��*�:� �[�t)}�����"���Ě��E��UE��D<}���[��~9� @�����4��4ꏿ�aN�*��$]��Yk�~��ϫ����M��~����ƽK��J���t��.��pG��+�;�>���J��   �   �⚾�N��Y0���Q����e���@�55����֭�������k��,��>�������^��������p?�B���(���:�z���*���H��Ve��4~�α���܊���~�~���e�.�H�R�*�B��1Z����p�����=�B�ѫ�2�Z��t�Ŭ��	u��"^�N��8����罃1�s=��b������ ������   �   !��徐%پ�RƾGa���}��T�o�K�;�5D�:7ֽ\��� ��ι��g��fTJ�k��K��(�)�܏m�W@����̿���jb���1���I�\�]��k�J�p�lXl�~�^�>�J��w2����r=��6�̿M؞�h�l���(����䴙��)G��������B��£��Ͻ@P
�zK7��0k��������Lľ�׾�9��   �   �#+��a(�W���7�.� ��ھC鲾ڌ�ʄV��" ����*Aʽl˽8U��F�4�����M�Ⱦw�� L��L��L��i4ܿ���L���,�z�<�8�G���K��aH���=�|�-��N�:���ݿ0���.U��K�K�fM�L�Ǿ�Ѕ��R2�.����Rƽ�Ľ��� |��ER�g��,)����׾����p������'��   �   �r��o�A'c�$>P��8�����z ���ʾ������e��h)�����@�'"���K ��e�s���%��oc)� �d�W;���Ǹ���ݿr� �
���m���%��)��{&��i������&�߿�繿�蔿.Ke�"�)����� ����c�������4��# �t&���a��s��; Ⱦ"���v���!6�gxN���a��Kn��   �   ˖�����2,������|���W�Z�1�Ɠ�@�־����rf��(�E��#����=�Y&?�Kч�V¾���E�7�o������|��/�ѿn���$ ����U	��P�<� ����ӷӿ)���떿h�p��8��P�B�¾������>�W�����u6���&��zc��ݜ��2Ծ���/���U��Bz�Vd��#;��m����   �   (ٿy�տָ˿���������񎿁l�&�;�c]�>�Ӿ�藾�/X��'������z���V��ߖ�� Ҿ�+� �9��i�ԋ��&-����mrʿoտ�ٿ�տ��˿����3���`l��|;��Z�f�Ӿ旾X,X��%������J|���V�,▾WҾ$.�7�9���i�!����/�����uʿ�տ�   �   �V	�zR�� ����ӿ����p�ا8��R�W�¾����^�>�t�����25�:�&��vc��ڜ�y.ԾA �,�/���U�0>z��a��K8��p����������G)��Z���)�|���W�Ή1���ݒ־H����f�)�(����E����>�\(?�Ӈ�¾����7��!o�����P���ѿ��뿘& �����   �   �)�~&��k����h���߿0깿�ꔿ>Ne�t�)����#����c�/������2��! ��p&���a��p���Ⱦ����+��#6�tN���a��Fn���r�x	o�e"c��9P��8�7���w �&�ʾ���w�e�Be)�X���>��!���L ��e�^�����}e)�Þd�=���ɸ���ݿ�� �¤��o���%��   �   ��K��cH���=�Z�-�:P����D	ݿ����V����K�O���Ǿn҅�VT2�����Qƽ�Ľ���Hx��@R��c���$��`�׾����	�����$�'��+��](����z4�� ���ھ�䲾m֌�GV�� ���=ʽnj˽kU��a�4�����7�Ⱦ���"L��M���M���6ܿ��M���,���<�p�G��   �   ��p��Zl���^��J�y2�����?����̿�ٞ���l�x�(����M����+G�O��5���6@���5ϽtL
��F7��*k����3���Gľ��׾�3�0��4��پrMƾ�\���y����o���;�@�1ֽ�W�����������zUJ�l����y�)���m��A����̿����c�r�1�P�I�n�]�R�k��   �   �݊�1����~�X�e���H�t�*�.���[�N���_���/�=�C�Mҫ���Z�,u�Ŭ��u�}^�v큽�3����6-�B�<��b� �����������ޚ��J���,��AN��g�e�x�@��0�<~����T����k��*�����$���^����n���q?����#���K;�F���*� �H��Xe�p6~�ᲇ��   �   �Ś��F�� F���=}��[��9��@�����5���ꏿ�bN���&^��8Zk�������8�M��{�����K�DF���o�����C���+���>���J���O�{�K�!�@�\�.�6t�����
�Ž�����Z���)��a%�r�[�����T��P�o����$N�4pP��*��y���Y�����:���[��*}�T���#���   �   挥��������������h�^C�� �l;��xɿ�����X������þ0"v��J��0���7�p-޼Կ���s����2�w}�D���!zн
��l	�`���/�Z����
�7���QDֽ)���V��^�@�Ĺ���ۼ|V���]F��֮�����{���ƾ��dU[� ���T˿nO�0�!��-D���h����}���j����   �   �̼��S��}���S��F1��<�X��1�2��zrݿ;���\p��s%�gfھR$���8'������
[��u�@�޼���H�8�"f�~f����ν������	��[������C���h,ҽ�'��򟃽 |@����X����o�c�Vƽ�)��ً���ܾ.�&��q�_ħ��߿����2�h�Y�����x���}����X���   �   я���2��/�������;��T��0.�$���ڿI㣿�l�P�"���־��z%�����Rnb��w��0�6� �9�\����������d�C&
����#��A'��1$�����������ŽN	���d��(��<�����j�v�ƽ�/(�b�����ؾ�$���m����uۿЙ�J /�ԹU����xA����-���   �   pa��v^��Uڜ��݋�ֲp���I���%�@\�п�+���`�k��v�̾;��ԗ ��]ýʗy�L�?��=D�:�w�������ڽ4�	��#&�Fa?��oS��r`�.e�
%a�s�T�QA��+(��#�s߽GW��� ���qL��G����V�ǽ�#�̾���sξp��4b�����%ѿP��v�&��]J�j�p��Ջ�I���Z@���   �   ��������̌��|��1[��[9�27�1����F��?
��
�N�o_�亼���r�����ǽ���������ϙ�$8ǽ���ْ)�~ER��3z�����A������+ک���X�����O�|���T�x!,�S ��˽���U���q���n�˽x��=u�]J��yR�#�O�ϴ������1t��v�0f9���Z��|�I|��_r���   �   믄�-���&Gt��]��A��@%�4F	�kEݿ�������}8�#������
]��)�K�н����߽�v|콓��$=L��!��\ڟ�����׾{��c���?���������N�ؾl����x��-����O��:����j����ڵ�B�Խ��$!_�Q2��P�����8�N߀�M^���iݿ�.	�L�$��A��*\��ls�칁��   �   ��^�ڊZ���N��<�d�&��>����p��'䔿Z�]��y�F�ھ�a���SF���d����.��4/��Qi�����������U�C)��-���6�E:��27�Z�-�-��b�����hþK��xl�4�1�����>余��<��f�G��)����۾�����]�wݔ��ֿ������,�%���;�>�M���Y��   �   �N7�W4��U+� h�@�x6��ȿ8���x� �8�2���A��dx{�'1�YM	�w����N��9��"z�8˧�(r۾�
��	)��{F�n�`�rgu�tc��ʃ�����#pv��b�(�G�a*�����eݾY��x�|�h�;�-��M� ��e
��2��I|�ӊ����;t8��_x������ǿ���~1����*���3��   �   |[�n��%��1 ��p�`�Ŀ~K�������H�Đ���Ծ]s��:lS��a��+��a�.�9��v{��s��Zm�`���r?�?sh������m���*����V4���k���⧿"S���房�(j�L�@�����󫭾14}�#;��F�J�����~�S�qU��qwԾ�"���G��ꁿSb���oÿU�������
�����   �   �e�����ۿ،ʿ5�����������K�����䀦��dn���0�ɿ�L���0��m��ϥ�@��=:�ToJ�82~�����|��G^ɿ�ڿ�M�[i꿝�濒�ۿ�ʿ�7��0������ܫK� ���|���hn�H�0�0��h���0� �m��̥���m7��kJ��-~�������Zɿ��ڿ*J��   �   1���h���ߧ�OP��[䈿�$j���@�����Ũ���/}�b ;�6E�?�����6�S��W���zԾH%���G��쁿�d���rÿ���m��� �
�ƺ��]�|��'�j3 ��s��Ŀ�M��֊��q�H�ے�{�Ծ?u��WnS�pb�+��_���9��q{�tp���h�N���n?��nh������j���'������   �   Xǃ�𩁿 kv���a���G�p]*����0aݾ�U��Q�|��;���h� ��e
�s2��L|�M���g��v8��bx�(�����ǿ���83���� �*�H�3�Q7�NY4��W+�j���?9��ȿ�9���x�2�8�����C���z{�)1�-M	�����PL��9�z�eǧ�0m۾г
��)��wF���`�>bu��`���   �   �@:�[.7�P�-�y��_�"��WdþzG���l�7�1� ���;佘��ͤ�(�G�X+���۾���!�]�!ߔ��ؿ�@������%���;���M�*Z�H�^�b�Z�J�N��<��&�@@���?���唿~�]��{�L�ھ�b���TF� ��b���� �=0/��Ki�矘�S}��5�쾺Q�|%�s-�6�6��   �   C9��M�������ؾ�����t��Ψ���O��6� ��x����ص�ԕԽ���"_��3������|�8������_���kݿ�/	���$��A��,\�Pos�H���O���� ���It��]���A��A%�:G	�Gݿ�������8�����;���]��)��н���Z۽��u�-��v7L�<��֟�����x׾q���\���   �   �թ���E�������|�U�T��,����d�˽����������r�˽8���>u��K���S���O�׵��� ���u��w�|g9���Z��|�w}���s�����Ӫ�� Ό��|�d3[�]9�8������G����(�N�0`�ѻ����r����*�ǽ�����}��*˙��1ǽȍ���)��?R�2-z������=��-}���   �   �(e��a�o�T��A��'(�* ��߽�R��E���lL�ިG�l��ǽr#�x����tξF��J5b�����&ѿ���B�&��^J���p��֋�8���YA��ob��g_��.ۜ�Uދ��p���I���%��\��пC,����`����̾R;���� �4]ý$�y� �?��7D�S�w�������ڽ��	��&��\?��jS�m`��   �   <?'�|/$����f�����Ž�����d���(�L:������j�Րƽ#0(�����d�ؾ8$���m����;vۿ.��� /�p�U�����A��u���.��Z���:3���������n<�|�T��0.�V���ڿ{㣿@l�|�"���־ ��z%�|����lb��u�v-�F� �/�\���������y`�$
������#��   �   �[������]����,ҽ�'�� ���x|@� ��(��h���c��Vƽd�)��ً���ܾ\�&�N�q��ħ�&߿����2���Y��������������X���̼��S��}���S��71�� �X�x1���Srݿ���"p��s%�(fھ"$���8'�B���w
[��u���޼@����8��e�cf��|�ν������	��   �   @?'��/$����f������Ž���x�d�d�(��9����-�j�ǏƽQ/(�2���j�ؾ$���m��
��Uuۿ��� /�n�U�V��A��{���-��H���02��������$;���T�,0.�Ƚ�ڿ�⣿Al�ǳ"���־~��2y%�r����kb��t��,��� ��\�|�������z`�$
������#��   �   �(e��a�w�T��A��'(�" ��߽rR�����~kL�8�G���ǽ�#�B����rξ���X3b�B��%ѿ���ڌ&��\J�N�p�)Ջ�n���g?��p`��y]��iٜ��܋���p���I�8�%��[�п�*����`����<�̾ :��j� �>[ý��y�v�?��6D�Ąw�������ڽ��	��&��\?��jS��m`��   �   �թ���H�������|�G�T��,�t���˽��|���F�����˽
��S;u�5I���Q���O���������r��0u�e9�j�Z��|�-{��!q��S��Q����ˌ��|�V0[��Z9�06�����SE��;	����N�R^�K���Q�r�؛�k�ǽӯ���|���ʙ��1ǽ����)��?R�6-z������=��4}���   �   O9��T�������ؾ�����t��¨��cO�~6�&������ֵ���Խ���_��0��A���F�8�Rހ�]��(hݿ�-	� �$�A��(\�pjs��������������Dt�~]�>�A�*?%�
E	��CݿH��r���8�����:���]�W'���н���ڽ�/u����Z7L�7��֟������׾{���\���   �   �@:�_.7�R�-�y��_���HdþcG���l���1�c��r9��������G�(��6�۾��b�]�ܔ��Կ�{��4����%���;���M��Y��^�F�Z���N�ڕ<���&�`=�,��a��┿̜]�x���ھ~_���PF�X�F_⽧��p��//�mKi�ٟ��O}��6�쾼Q��%�x-�=�6��   �   [ǃ�󩁿kv���a���G�l]*����aݾjU��܊|�*�;������ �c
�2�F|�u���� ��q8��\x�,�����ǿ	���/��}�چ*���3�VL7��T4�~S+�(f���z3�)�ȿ�5����x�p�8�K���>��Ft{��1�aJ	�@���0K�_�9��z�Kǧ�$m۾ϳ
��)��wF���`�Dbu��`���   �   1���h���ߧ�NP��Y䈿�$j���@�����꾎���#/}�D;�uC���������S�"S��GtԾ� ���G�避`��mÿ?��N���~
����dY�\��#��/ �>m係�ĿI�����n�H�X����Ծ�p��2hS�Y^�S(�H^���9�Uq{�Ip���h�J���n?��nh������j���'������   �   �e�����ۿڌʿ5���������}�K����羗����cn���0�R�����u|0���m��ɥ�*���4�ahJ��)~����������Wɿ�ڿ�F��a�;�濄�ۿ��ʿ2�����7���K���~�澥}���_n���0�x�����?~0��m��̥����f7��kJ��-~��������Zɿ��ڿ/J��   �   ~[�p��%��1 ��p�]�Ŀ{K�� �����H����O�Ծ�r���jS��_�>(��\�,�9��l{�m��&d�m��Tk?�ejh�z��g���$�������-��{e���ܧ�eM���ሿ j���@����<����9*}�;��A������*�S�U��8wԾ�"�z�G��ꁿTb���oÿY������
�
�����   �   �N7�W4��U+�"h�>�v6��ȿ8���x��8���LA��Fw{�`1��J	�n���I�ڲ9�xz��ç�yh۾߰
�F)�]sF��`�&]u�^���ă�9����ev���a���G��Y*�~��\ݾ�Q��4�|�6�;�]��H� ��b
�#2�}H|�������3t8��_x������ǿ���~1�����*���3��   �   ��^�ڊZ���N��<�b�&��>����n��$䔿Q�]��y��ھa��bRF���6^⽂�ཾ���+/��Ei�=����x�����{N��!�r-���6�l<:�*7�6�-���%\�G��s_þ�C���l�Z�1�R���5�$�����G�R)��E�۾�����]�wݔ��ֿ������,�%���;�@�M���Y��   �   믄�.���&Gt��]��A��@%�6F	�kEݿ�������q8���������	]�(�^�н���$ֽ�Ao���2L����ҟ��׾��뾅V���2���������Dzؾ����Vp��4���� O�2��������ӵ�L�Խ,� _�2��&�����8�N߀�P^���iݿ�.	�L�$��A��*\��ls����   �   ��������̌��|��1[��[9�27�3����F��=
���N�a_������r����b�ǽl����y��gƙ��+ǽ���J�)�:R��&z�-���u9���x��cѩ�[馾	�����ݠ|�d�T��,�}����˽b��@���P����˽I��O<u�&J��lR��O�ϴ������3t��v�2f9���Z��|�J|��_r���   �   oa��u^��Vڜ��݋�ֲp���I���%�@\�
п�+���`�b��T�̾�:��� �s[ý4�y�4�?��1D��}w��×ڽ�	�t&�X?��eS�9h`�G#e�ga�U�T��A��#(�r�R߽`M�����~eL���G��쀽�ǽ#������sξi��4b�����%ѿP��x�&��]J�j�p��Ջ�I���Z@���   �   ҏ���2��/�������;��T��0.�$���ڿI㣿�l�N�"�}�־����y%�����$kb��s��*��� ���\����������\��!
�R���#��<'��,$�:��������Žv��l�d�b�(��6�z����j�W�ƽE/(�D�����ؾ�$���m����uۿЙ�J /�ԹU����xA�����-���   �   �������ey��������Vgd���9�D�����3����,|��=.���澜���[P3���ӽj"x�J$ �D�>�;�S������ⷽХཎ��F��64��{�_t�gg��+�"�����e���NW��l!�b��#��{��սP�4�Sw����)�.�9}�78���迀�pY:���d�E(�������������   �   �9��륿��d��rc������.`�
�6��H�@�Zի��x��Y+�r��&����x1�*�ӽg���.�,��tw;�p�y���ďӽ�N ��q�6^$��.�?2�Q�.���$�j���n?սح���}���>��!�2�����q�սk�2��J����㾮,���x��g�������07�P�`�9G���|��mj��V����   �   Ub��d�������S�� <~��:T�,�-�·���ٿ����Gl���"��'ؾ�Z���O,��Yսۋ��`[��F`��Ԋ�`���ӂ�����1�,L�P�`�J0n�[�r���n�da�~�L�1�2����nq�Μ��
����c�Z�^�؟���I׽�p-�Q���
پ�#�n�l��6��Pڿ���4).�,}T�r]~��O����������   �   ���������A���}����f�`B��I ���@ɿ(	���SY�����Ǿ������$�Ēٽ�~���ٔ����dٽ\�c�5�Q`�tބ������N���ۯ��9��2���������n���Fa���6���]۽'ޫ�X����1�� \۽|�%�����w:Ⱦ�o��Y�?]��6�ɿ0��i ��eB�@�f��Z��������   �   ́��������J�h��$K���,��m�rG翚���Ć��A�*���Ĳ��4k�a�b��ýerϽ` �9'��Y�~<���N����Ǿ������hH�N��Kl���l���xȾ�������,[�U(���,ѽ�Ľ^��.���'l�6Q�������A�y�E@��Z�
b�t�,�p�J�h�-����[���   �   .lj�\�e�r�X���E�J].����L&����ȿ䛿�h���&�V����yIS���0�����'g�cx;�>Cx�jʡ��̾إ�����&u&�x6��@�V�C�T6@��\6���&�3Q�����tv;������y���<�`D����5u��=���S�%b��I���&��h�᛿8�ȿ9����F���-��E��vX�d�e��   �   �%@���<��*3�a$�z�ͬ��u�ѿ앨��\����A���
�-`���F��6�<�`u�8F	�.���IF��ڄ�[������6�l�1��P���k����ަ������ʇ�� ����l�^Q��2�*��k��R���g���"G�ě�@�	�&��sQ=�>w��6�����
�f�A��<��U��(Kѿ���Ү�(�#�"�2��<��   �   ��F��":�����K��CͿ��������pgR����%ྂ蝾&�`�?*�=����6F��m��)^���4������\I��3t�h����ڠ�����8���l���k���t���K��&��yu��J��| �*���*x҅���F��U�Ą��m*���`�F۝�K�߾e���R��N���/����̿o�� X�����h��   �   ����g�B��fӿQ&��T����ԅ�[U���#�������ig|��P<� �����7"<�b|�C���g�,a#���T�n��t ��������ҿ��������:���piӿM)��餡��օ��^U�p�#�l�򾽕���j|��R<�������<�R|��?��5c�<^#�(�T��k����������ҿ�����   �   �i���h��Pq���H��f#���u�
J��y ������궾1Ѕ���F�(T����3o*�^�`��ݝ���߾���&R��P��U2����̿ؓ��Y����k���p��(<�λ�OFͿप�����gjR����(�~Ꝿa�`��?*��<����2F�k��}Z���/��`���XI��.t������נ�l���5���   �   ����Ǉ������l��YQ�^�2������NN���d��KG����N�	�q��S=��x��ʅ��m�
�	�A��>��MW���Mѿ������>�#�r�2�f�<�:(@�@�<��,3�c$�2�����߻ѿᗨ�H^����A�9�
�Mb���G��F�<�4u��D	�����EF��ׄ�Z���ݰ羝3���1���P���k�f�������   �   ʃC��1@��X6��&��M�ʚ���q;̉���y��}<��A��
��)t���=�{�S��c������&���h��⛿a�ȿ����*H���-�E�yX�0�e�oj��e���X�ΌE�_.�(���(����ȿ�囿[�h�A�&�x��X���JS����P������c��s;�=x�fơ���̾ʟ��s��3q&�0�5�i�?��   �   �� i��������sȾ�	��p튾'[��P(����'ѽ�Ľ������)l��R�����k�A����A��\�Hc���,�Z�J�lh�����O]��Q���]���7��x�h�T&K���,��n�%I�����ņ��A�$���Ų�6k���$��ý�mϽ� �z4'�%�Y��8��J����Ǿ�������E��   �   /5�����ܪ�������k���@a���6��W۽�٫�����60��\۽C�%������;Ⱦq���Y�Q^����ɿ�0��j �gB��f��[����e��g���3���C���~��&�f�LaB��J �\�Aɿ�	���TY�����Ǿ#���)�$��ٽ�|��6֔�����]ٽ8 �F�5�5`��ڄ��~��zJ��&ׯ��   �   ��r��{n��^a���L��2��~�ik����V���ιc���^�����I׽�q-����پ�#���l�]7��Qڿ>��
*.�D~T��^~��P���������ec��f������vT��.=~�j;T���-�H����ٿ���l�f�"�X(ؾ�Z�� P,�-Yս�ً�l\[�z@`��Њ�$���f|���2�1�?L���`��*n��   �   �<2���.�0�$�(���<ս���A}�:�>�x!��2�Ȳ����ս�2��J�����;,���x�&h�����v��V17���`��G��J}���j��飿�B:��q���e���c��'��/`�T�6�0I�c@俏ի�x�Z+����8���}x1���ӽ�����.����Ns;�5�y���ӽ�L �`o��[$�j�.��   �   �{�et�tg��+�("�����e��4OW� m!�tb�`�#���{�v�ս��4��w��2��Y�.�t}�[8���还��Y:���d�V(������������������Yy��������8gd���9�,���������,|�j=.�F��i���P3�P�ӽ�!x��# �������S�f���nⷽ��ཅ��>��24��   �   �<2���.�5�$�)����;ս����}���>��!��2������ս�2�QJ�����{,�~�x�qg�����ܷ��07��`��F��d|���i��Ϣ��$9��X���d���b��q��.`���6��H�y?��ԫ�x�[Y+���⾐����w1���ӽl����.�p��s;��y���ӽ�L �co��[$�o�.��   �   ��r�|n��^a���L���2��~�Jk�Η�������c�S�^�Ν���G׽�o-�����	پx�#���l�6��[Oڿ���(.�L|T�B\~�O��������Fa��U�������R���:~�x9T�Z�-�*����ٿ����l���"�m&ؾ�Y��cN,�WսR؋��Z[��?`�bЊ�����U|���4�1�GL��`��*n��   �   65�����᪦������k���@a���6����V۽!٫�^���b.��Y۽��%�̏��C9Ⱦo���Y�m\��"�ɿP/��h �zdB���f��Y������ߟ�����z����@���|��Թf��^B��H ����>ɿ���QY�����}Ǿh�����$��ٽ�z��Ք�N��0]ٽ �8�5�3`��ڄ��~���J��-ׯ��   �   ���i��������sȾ�	��h튾�&[��P(�z��&ѽ��Ľ���=��[%l��O������A�t��>��VX��`��,���J��h�ᫀ�aZ��J���o~�������h��"K��,�jl�vE����Æ��}A�Й��²��1k����㽸ýSlϽ� �@4'��Y��8��J����Ǿ���ʕ��E��   �   ЃC��1@��X6��&��M�Ś���q;������y�_}<��@�?��jp���:���S�k`���
�#�&�ƛh��ߛ�Q�ȿ����$E�$�-��	E�tX���e�Vij���e���X�p�E�f[.�"���#����ȿO⛿qh���&�q�����:FS������2��>c�es;��<x�Vơ���̾ȟ��t��6q&�4�5�p�?��   �   ����Ǉ������l��YQ�[�2���s��*N���d���G�_��l�	�����N=�ku��������
��A�Q;��*S���Hѿ�����0�#��2�~�<�0#@�V�<�0(3�_$�������Ҷѿ����[����A���
�I]���D����<�Hr��B	�`���DF�fׄ�<���Ѱ羛3���1���P���k�i�������   �   �i���h��Sq���H��e#���u��	J��y �u����궾�υ�¿F�]R����j*��`��؝���߾%���R��L��v-���̿4��,V�����f�\���8���ZH��@Ϳ��������"dR�!�"��坾�{`��;*��9�E���1F��j��OZ���/��Z���XI��.t������נ�o���5���   �   ����i�E��fӿQ&��R����ԅ�[U���#�T�򾻒��gf|�5O<������g<��|��<�� _�[#���T��i��)��������ҿV	�I������񿍆忥bӿ3#������@҅�DWU���#���򾦏��Yb|��L<�������B<�T|��?��c�3^#�%�T��k���������!�ҿ�����   �   ��H��$:�����K��CͿ��������ggR����%�蝾�~`��<*��9�����.F�nh���V�� +��]��UI�|*t�����Ԡ�A��E2��&f��%e��n���E��� ��0�t� J��v �����涾Fͅ�n�F��P�j���k*�+�`��ڝ��߾W���R��N���/����̿r��X�����h��   �   �%@���<��*3�a$�z�̬��s�ѿ镨��\����A���
��_��(F��c�<��r�
B	�$��HAF��Ԅ������羈0���1�4�P���k�����=�����Ň�a�����l�7UQ�s�2�ο�=��)J���a��jG�����	�V���O=��v�����q�
�]�A��<�� U��)Kѿ���Ԯ�,�#�&�2��<��   �   0lj�\�e�t�X���E�J].����M&����ȿ䛿�h���&��澠��HS��������p`�:o;�7x��¡�2�̾������\m&���5���?�HC�i-@�{T6� �&�AJ������l;�����zy��x<��=�?���n���:�9�S��a�����&�
�h�᛿9�ȿ=����F���-��E��vX�f�e��   �   ΁��������J�h��$K���,��m�rG翙���Ć��A���iĲ��3k���D�xý3hϽv
 ��/'�s�Y�C5���E����Ǿ�⾑����A�����e�����㾖nȾK���銾� [��K(���!ѽŮĽ@��z���&l��P�������A�z�H@��Z�b�v�,�r�J�h�.����[���   �   ���������A���}����f�`B��I ���@ɿ(	���SY����NǾB�����$��ٽ�y��JҔ���HWٽ?��e�5�R`�zׄ��z��>F���ү��0��,�����������g���:a���6���4P۽Oԫ����T,��VX۽C�%�O���A:Ⱦ�o��Y�?]��9�ɿ0��i ��eB�B�f��Z��������   �   Vb��c�������S�� <~��:T�,�-�·� �ٿ����Dl���"��'ؾHZ��O,�ZWս�׋�tW[�,:`��̊�'���Nv�n����1�zL���`�2%n��r�kvn��Ya���L���2�{��dｒ���ݙ����c���^�k���BG׽	p-����
پ��#�m�l��6��Pڿ���6).�,}T�r]~��O����������   �   �9��륿��d��rc������.`�
�6��H�@�Yի��x��Y+�b�����'x1���ӽ��Z�.����o;���y��륽��ӽ�J �!m�6Y$�ә.�):2��.���$�����B8սʧ���
}���>��!�x2�F���O�ս	�2�eJ����㾬,���x��g�������07�P�`�9G���|��lj��U����   �   �x��;����/���e��b���D�g��G<�N��m�꿭��U��
1���꾙ԕ�pD8���۽DY���-��g���+��a�N
��b���.������:8��^!�[(�v��tn�j1轔��O���aa���*�j����,��䂽\۽��7�����`��"�0�b���ܰ�+��rl��$<��zg����L\���+�������   �   ����i������������Cc��9��'�:�0��2�{��.�s�b����b6�P!ܽ�/���j<�M+��PI����<���~�۽�p�����(�Z�2�oW6�a�2�Ӆ(�����?��۽������vH�bu*�g�;�6�����۽�6�3t�������-�dz{����������8��%c�E��'���p���j���   �   
��������|l��؀�B�V�.�/�z@��ܿP���m�o�P�%�kܾ5\���1���ݽK:��քi�v~n��8����������� � �6���P���e��s�P�w�Ds�B�e�·P�sP6����6d�����đ���m�ةh��ɒ�uݽ��0��0��}�۾�s%�PTo��ץ��aܿ,���/���V�Ԁ��m��� ������   �   o#��>���F��7����i�l�D��!"������˿�
���w\��b�z'˾у���)�N��`��<D��Һ��$�ὲ~�
�:�Spe�`���Y��� b���벾�1���޲��I��6c������$e�ID:�j9����E��L֛������7έU)�ګ����ʾ�E��T\� �����˿�|�@"���D��i�|@���Q���E���   �   u���L���y���0k�TWM�F�.������鿞B��c���|FD���������p�h}!��&뽒�ʽtf׽9X���+�/@_�	?��Ш���c˾��澇����I�3��}@�~����S3˾x��	��i�^���+�q�r�ֽ�tʽ���4H!�GGp��������0D�G|��e9����n��:�.�RmM�rNk�c���-V���   �   �em�ġh��F[��G�t0���c����ʿ����k�)��m�f���.X�H��#������`��f]@���}�f���aо'���m6��)�F�8���B�bF� �B�ʒ8���(�p�����c'о&⤾��}�_@����N��������X�瞾OW�W�(�5}k�O����˿�����V)0�$�G�le[���h��   �   ^B�T�>�X�4���%��l���O�ӿab���⃿�KD����C�ľ�懾!bA�j���Y�9D��)K�������������:�4���S��\o��~��d������Z��Jn���2o���S�~�4������!״�ޑ��s�J�0�6��v�UGA�xۇ��ľ����RD��냿�s����ӿI.�����T&�r5�b�>��   �   ����$�H�����;q�-ϿMT��8��H�T���x�����e�f.��?�0#�n�J��0��#���6`���"��nL���w�j�������W��s��#����e��A@��O袿"���~�w�E@L��]"��*��㗹����J��#�O-�[.��e��������|'���T��(��jr��VϿ��*	���J1��   �   ߑ��À����=`տ�齿�3���4��x�W�5�%�I8��hO�����ai@�f� �O� �3y@�;����h���`����%�r�W��R���X��;���տ7��-��Օ������翚cտ�콿6��7����W���%�C<��(R��ޅ��>k@��� �f� ��v@�0����e��}\����%���W�5P���U������տw��B���   �   ����cb��
=��X墿~����w�{<L��Z"�&���������2�J�n#�>-�S\.��e����:���)� U��*���t��YϿ�������3�����&�T������t�f0Ͽ�V��$��F�T�L��{�����!e��f.�?�V#��J�N.��n���1[���~"��jL�-�w�����x���T���o���   �   &����W���k���-o�V�S���4��|�Џ�`Ӵ�&�����J���5� w��HA�݇���ľ���BUD�\탿%v��I�ӿq1��f��p&��
5���>��`B���>���4���%�dn�����ӿ\d��.䃿.ND�8��n�ľ�燾8cA�A���X��A��%K��������o�뾺��F�4�9�S��Wo�4|��.a���   �   �F���B���8���(��������"оTޤ���}�*@�(���K��t�������X��螾�Y�I�(��k����˿J�����@+0�l�G�
h[�b�h��hm���h�4I[�2�G�>0�2�Ŭ���ʿ����k��)��o꾳���O/X�`��0!������*���X@�s�}�U���\о����2��)��8�t�B��   �   Ϫ�+=��w��^��D.˾�s��z����^�S�+�S�L�ֽ�rʽ0���H!�'Ip�0���J��{2D��}��;���鿮��ƹ.�DoM��Pk�ŉ���W���v��:N���z���2k�YM���.����[���C��i����GD����
����p��}!��%뽝�ʽ�a׽�T�8�+�-:_�L;��O���t^˾���"���6F��   �   �,��"ڲ�ZE��G_�������e�c?:��5���vA��wӛ�����7�{V)������ʾG�,V\�5���W�˿�}�X"��D���i��A���R���F���$��f?���G��8��V�i���D��""�r����˿����x\�^c�x(˾�у��)����N ���@��������ὅz�ވ:�$je�ȶ��Q���]��G精�   �   ��w���r���e��P�+L6���^��<��$���N�m�p�h�,ɒ��ݽ��0�71����۾�t%��Uo�aإ��bܿ�,���/���V��Ԁ��n���!��0�����������Em���؀�&�V���/��@���ܿ����7�o�֘%�ܾ�\��&1�-�ݽ�8��d�i�*xn�b4��X���6��������6���P�6�e��s��   �   �T6���2�X�(�H���=�v۽4������<sH��r*���;������۽b6��t��I��}�-�({{���Q�V��8��&c����������k��7	��Xj��M��鿠�Q��^Dc��9�"(�i:�K0��|�{�.���v���|b6�� ܽ�.��_h<��I+��LI� ������|۽�n�>��|�(���2��   �   �^!�^(�����n��1轷��|����a��*�В��,�0傽o\۽�7�񢕾���S�0�����ܰ�U�꿊l��$<�{g����\\���+�������x��5����/���e��R���$�g�|G<�6��B�꿉�����	1����eԕ�$D8�V�۽�X����-�`g�$�+���a�&
��>���������48��   �   �T6���2�Z�(�I���=�s۽,��œ���rH�rr*��;�U����۽�6�t��D�澽�-�z{�^��e翼�B�8�~%c����¸�����j����<i��?���������FCc�9��'�{9翕/��n�{�Q.���ɣ���a6��ܽ.��zg<�`I+��LI�������|۽�n�A���(���2��   �   ��w���r��e��P�,L6���^��������G�m�ʤh��ǒ��ݽ��0��/����۾Ss%��So�ץ�aܿ�+��/���V�gӀ��l�����������멵����k��U׀�&�V�V�/��?�ׄܿ~���0�o�f�%� ܾB[���1�~ݽ�7���~i�"wn�4��&���&��������6���P�@�e��s��   �   �,��(ڲ�bE��K_�������e�V?:�d5��὿@��Tқ�>����4�6T)�����R�ʾE�[S\�N����˿B|�V"�l�D�X�i�w?��\P��5D��"���<��=E���5���i��D�� "���?�˿�	���u\�aa��%˾�σ���)����x����?��B���8��gz�͈:�je�ɶ��U���]��O精�   �   Ԫ�0=��w��e��F.˾�s��t����^��+�����ֽhpʽ���@F!��Dp������ /D�@{��8��I��X��ֶ.��kM�:Lk�����T���s��=K��'x��X.k�dUM���.�������A��"����DD�e������p��z!�"�n�ʽL`׽^T���+�:_�D;��L���w^˾���+���<F��   �   �F���B���8���(� ������"оBޤ�{�}��@�o��:I���������\ X�a垾�T꾨�(��zk�̹��  ˿G������'0���G��b[���h��bm��h�D[�G��0�$�������ʿַ���k�)��j�G����*X�q��f��:���l��YX@�4�}�C���\о����2��)���8�z�B��   �   *����W���k���-o�V�S���4��|����@Ӵ���J���83�.t�jDA��ه���ľ���;PD�ꃿ�q��/�ӿ]+��Ԇ�R&�,5���>��[B���>��4���%��j�������ӿ/`������&ID����V�ľp䇾�^A�L���V�]@��$K�M������^�뾷��D�4�:�S��Wo�6|��1a���   �   ����gb��=��[墿~����w�x<L��Z"�&��R���q���J��#�p*�X.�+e�D���[��5%���T��&��p��JSϿ˞�P���/�J���"�2������m�*Ͽ�Q������T����t�D���`e��b.�3<��#���J��-��=���[���~"��jL�-�w�����{���T���o���   �   ���ǀ����@`տ�齿�3���4��r�W�)�%� 8��O�������g@��� �f� �Ws@������b��^X��1�%��W�N��_S����E�տ���k������|�:���\տ�潿�0���2����W�4�%��3��L������ee@��� ��� �4u@������e��V\����%���W�5P���U������տ{��G���   �   ����$�J�����<q�-ϿLT��6��@�T��lx㾡���6e��c.�#<�!#��J��+��߶��xV���{"��fL���w��������OQ��Dl��C����^���9��O⢿����$�w�s8L��W"�� �����������J���"��)��X.�me�C���q��m'���T��(��kr��VϿ��,	���L1��   �   ^B�V�>�Z�4���%��l���O�ӿab���⃿�KD�{���ľ懾K`A�����U�!>�#!K����� ���p�뾚����4���S��Ro��y��[^��E���U���h���(o�țS�Ǌ4�`y����6ϴ�􋇾��J���1�t��EA��ڇ���ľ����RD��냿�s����ӿJ.�����V&�t5�f�>��   �   �em�ȡh��F[��G�t0���c����ʿ������k��)�Gm������,X���V��������"T@�b�}�r���Wо"���j/���(���8���B�=F� �B�;�8���(�q�����rо2ڤ�7�}�@�8��,E������ˬ��X��枾W�G�(�0}k�O����˿�����V)0�&�G�ne[���h��   �   u���L���y���0k�VWM�F�.������鿟B��b���sFD�������s�p��{!��!�*�ʽ$\׽?Q���+�i4_��7������dY˾-������B�o���9�sq�����	)˾Co���	����^�r�+�z�'�ֽpmʽ��~F!�/Fp�9������0D�F|��g9����n��:�.�TmM�rNk�c���.V���   �   p#��>���F��7����i�l�D��!"������˿�
���w\��b�B'˾�Ѓ�q�)��������<���7�ὀv��:�-de�N���d{��VY���ⲾS(���ղ�A��E[�������e�,::�81���;���Λ�0����3�xT)�x���O�ʾ�E��T\� �����˿�|�B"���D��i�}@���Q���E���   �   	��������}l��؀�D�V�.�/�z@��ܿP���l�o�G�%�Jܾ�[��51�T~ݽ�6��R{i��qn�T0��K������I��e�6���P��e�Xs��w��r���e���P��G6����W���������
�m�X�h�|ƒ�ݽ�0�D0��Z�۾�s%�PTo��ץ��aܿ,���/���V�Ԁ��m��� ������   �   ����i������������Cc��9��'�:�0��1�{��.�c�D���%b6� ܽ�-��f<��F+��HI�����.}��Fy۽�l�����(��2�R6��2�ɀ(���a;��۽��� ����nH�:o*�Ë;�����l�۽z6�t��x����-�cz{����������8��%c�E��'���q���j���   �   �������=��+=�����ܷa�t8��v��>��~��O�z��-�M�澓b��j�5�T	ڽ�=��f=/�BS�F-��db�����q���>���y�v��H����TP��
�v佈��������A]���'�F4�P*��u��#�ֽ�3�:���]�,��ty�I����忤���M7���`�,���h���'���{���   �   ����0��t0��K���i���]�P�4������޴����v�۲*�M���;��N�3��Fڽ���;�=���,�?>J��ރ�������ٽ������:&�;0��S3�Ϭ/�]|%�H����B׽�橽�;��tE�
�'��]8�r=��.7׽�-2����d`�v�)��eu�\⩿/�� ~�BH4�f�\��ڄ�����w(���3���   �   ����ï������Ñ��fz�ޖQ��,��Q
��ؿ����P�j�@W"��	ؾo����.�b�۽�ƒ���i�B�n�$Α��F��Ut�e%��4�r�M���a���n��"s��cn��a�~�L�֧2�������l��=�� ei�K�d����N�ؽz-��	���־U�!���i�롿=׿�	�؝+��8Q�8z��ɑ�@���گ��   �   Oՠ�����~���*��/c��?����؋���ǿ�ޕ���W�=^��kǾ���G['��߽4��>���B���ڞ߽r��D
8��a�����pї�E��v{��{����-��H���{�������;`��T6� 5�#�ܽ�譽^���Y���N�ܽ��%��΀� Zƾo��$W�f����ƿ
���X�:�?��_c��]��ٺ��/0���   �   ;+������0}�P�d��H�Ё*�b������\�������.@������|�l��^����/ɽi�սg����)���[���������ͭǾ�w����~������W����%{�r�ƾ{���T뉾�Z��(� v�Y�ҽ��ƽb潨�@k�u�3���?�W^��K%��Ϸ�:��j�*�$zH��3e��}��E���   �   ��f��8b��PU�(SB�Ƴ+��x������vƿY@��vbf��q%���<��z�T����H���������=���y��F��5�̾�4���O�ӣ%��4���>���A��?>�U4���$�Ē�1���(Q˾#$��<x�<�ܠ�N����5�����\�S�m����4��4%��<f�\F��q�ƿ&s��
���M,��	C�L�U�ܟb��   �   L�=��:�lm0�Z�!����u��a�οZ��,瀿��?���	������q��%T>���\�����H��x��ұ�[o���"01�ՔO��{j�����t��5����@����~�@�i�E�N��=0�>��,澢���褄�r�F�t�H�
�/����=��+�� x����	�0@�����ަ���ϿL��"����"��1��w:��   �   �A����~(�j����꿯Mʿ�H���چ�`�O�U����޾�q���a�á+���J� ���G��م�hU��<���UP��]H���r�?ˍ�������ހ���l���6��o*��c��� ����q��XG���� j��|��A����F�f" �C���\+��`�����U�޾���̇P�zL����v/˿U��FN���p���   �   �.�c
l�haпj��XO������ӝR���!�n������%�{���<�)�A�
M=�L�|����X��щ"��S������I��nAѿ&�tu2�(�Dp⿳dп�l���Q�����D�R�R�!�Q��q����|�� =��)�3@��J=�M�|�}��	~��"�TS���������F��>ѿb"㿠q��   �   qi���3��M'��}��4�� �q��TG�����e�y���>����F�! �1���]+���`�K�����޾X��
�P��N��H�i2˿���(P�������C��z*�8�����sPʿMK���܆�O�O������޾�s��a���+�{�z� �n�G�jׅ��Q��U���&M��YH��r��ȍ�ﳟ�R����}���   �   _����=����~�k�i���N��90�5��Z�����?�����F�F�X�
�t���=�B-���z����	��@����ᦿ[�Ͽa������"� 1�>z:�ħ=�(!:��o0�P�!�Z��S����οM����耿�?�G�	�ɪ��s��8U>��������H��u��$α�4j����C,1�\�O��vj�#���q���   �   (�A��;>��P4���$�i��u���uL˾i ���x��<�������4����#�S����Y7��6%�:?f�H����ƿ�u�����`O,��C���U���b���f�L;b�jSU�>UB���+�z������xƿ�A���df�@s%�6�征����T����6F���������_�=�s�y��B��<�̾�.��[L��%���4�0�>��   �   ����T������uᾁ�ƾG����牾-Z�}(��r�D�ҽl�ƽ�a�_��Ak����r���?��_���&��ƹ�p����*� |H�D6e���}�G���,��W��3}�r�d��H�*�*�t��M��T^�������/@��²���l��^�r��),ɽ�~ս��&�)���[� �3�����Ǿ�q�̖��6���   �   񈲾^)��������L����5`��O6�P1�N�ܽ�䭽��������H�ܽt�%��π�n[ƾ����%W�+g����ƿ����Y���?��ac��^������1���֠�7������+���0c�0�?����:����ǿmߕ���W�_��lǾ�����['�N�߽*��瘛�}���q�߽U��48���a�~��͗��@���v���   �   ?s�!^n�Ua�ĊL���2�x����,h������_i���d�0����ؽ&-�M
��&�־/�!�ƚi��롿>׿��	���+��9Q�p9z��ʑ�9���$ۯ�����į�����}đ��gz���Q�(,�TR
��ؿ����j��W"��
ؾ����.�̓۽�Œ�r�i��n�ʑ��A���m�!�h�3���M���a�,�n��   �   "Q3�<�/��y%�������ֽ�㩽T9��E���'��\8�:=���7׽".2���a� �)�fu��⩿˓�b~��H4��\�0ۄ����)��z4��'����0���0���������T�]���4�,��������v�
�*�����;��D�3�tFڽ8����=�d�,�:J�H܃�b����ٽ������}7&��0��   �   H����_P��
��佧�������B]�T (��4��*�v����ֽU�3�P:��\徍�,��ty�n��� 忼���M7��`�<���w���'���{���������=��=�������a�X8��v��>濨~���z��-���`b��"�5��ڽ�=���</��R��-�kdb�v���N���>���r�p���   �   &Q3�A�/��y%�������ֽ�㩽>9���E��'��[8��<��z6׽P-2�h��"`�D�)�xeu�'⩿���}��G4� �\��ڄ�4���(��e3�����~/���/��˵�����F�]���4�����a����v�M�*���N;��k�3�dEڽ������=���,��9J�.܃�R����ٽ�������7&��0��   �   Ns�+^n�aa�̊L���2�r����h��Q���^i�Y�d������ؽ�-�	��C�־ɀ!�Θi��꡿_<׿��	�:�+��7Q��6z��ȑ�\���ٯ�����¯�������dez�̕Q��,�4Q
��ؿ�����j�\V"��ؾ���f�.�۽8Ē���i�
�n��ɑ�wA���m�!�h�3���M���a�6�n��   �   ����d)��������N����5`��O6�41��ܽ�㭽y���.��x�ܽ?�%��̀��Xƾ����"W�Qe��u�ƿ����W��?�\^c��\�������.���Ӡ����V}���)��`-c���?����'�����ǿ�ݕ���W�]��iǾɭ��JY'�t�߽Z������Ħ���߽8��8���a� ~���͗��@�� w���   �   ����T�����uᾆ�ƾF����牾Z�F(��r���ҽL�ƽB^潿��=k���'����?�W]���#��!��,���*�rxH��1e���}�&D���)��}���-}��d� H�P�*�*�����j[��c����,@��
�������l�F\����)ɽZ}ս����)���[��/�����Ǿ�q�Ֆ��;���   �   .�A��;>��P4���$�k��u���nL˾[ ��Tx��<�^��¡��,1��@����S�����d2�63%�a:f��D����ƿ�p������K,��C���U�2�b���f��5b�~NU��PB��+�$w������tƿ�>���_f��o%�:��&��B�T�	��yB��|���&���=�/�y��B��0�̾�.��ZL��%���4�6�>��   �   c����=����~�o�i���N��90�3��M�޻�����!�F����
������=��)���u��3�	��@�v��	ݦ�]�Ͽq��r���"��1�lu:�֢=�Z:�*k0�R�!����e����ο5}��u倿.�?���	�Υ���o���P>�~�&�����H��u��α�"j����A,1�\�O�wj�(���q���   �   ui���3��P'�����6�� �q��TG�����e�[y��w>����F�G �r���Y+�y�`������޾���لP��J��t�,˿"��xL���R��~?����v&����)���Jʿ~F���؆��O�׊���޾o���a�O�+����� �M�G�ׅ��Q��6���M��YH��r��ȍ�𳟿U����}���   �   �.�g
l�kaпj��YO������ҝR���!�G��x���/�{�a�<��&�C=�PG=��|�����y�;�"��{S�����A���C���:ѿ���m��*��i�^п�f���L�������R���!����n���+�{��<��%��=�I=�L�|�1���}���"�OS���������F��>ѿf"㿤q��   �   �A�����(�l����꿱Mʿ�H���چ�Z�O�F��l�޾oq��pa���+���V� ���G��ԅ�MN������*J��UH���r��ō�	���0���:z��f��D0��$��������t�q��PG��~��`��u���;����F�r ����Z+���`������޾���ćP�wL����u/˿V��HN���r���   �   L�=��:�pm0�\�!����w��a�οZ��*瀿��?���	�W���Bq��ZR>�R~�;����0H�s��Xʱ�Ne�����(1��O�)rj���/o�������:��Z�~�x�i���N�60� ��-	�뷰�"����F���(�
�f����=�"+���w����	�&@�����ަ���ϿL��"����"��1��w:��   �   ��f��8b�QU�,SB�Ƴ+��x������vƿY@��pbf��q%�ڼ�����T����lA��F���b��Ξ=�~�y��>��x�̾)���H��%���4�Ҁ>���A�/7>��L4���$���~���zG˾f��:�w�<�<��̝��Q/��U���S�����}4��4%��<f�[F��q�ƿ's��
���M,��	C�N�U�ޟb��   �   <+������0}�R�d��H�Ё*�d������\������.@������l�l��\�����'ɽLyս�����)�?�[�����󣩾��Ǿ1l⾰������_��UQ������o�m�ƾ䇨�4䉾9Z��(�4o�H�ҽj�ƽ]����>k�"����?�V^��K%��з�<��l�*�$zH� 4e� �}��E���   �   Oՠ�����~���*��/c��?����ً���ǿ�ޕ���W�0^�TkǾ����Z'�p�߽����������%�߽b��U 8�(�a��z���ɗ��<���r��o����$��ح�����Σ���/`��J6�!-���ܽ6߭�(���#}����ܽ�%�x΀��Yƾa��$W�f����ƿ
���X�:�?��_c��]��ں��10���   �   ����ï������Ñ��fz���Q��,��Q
��ؿ����O�j�:W"��	ؾ2���.��۽Ò�w�i�ɥn�Ƒ��<���g���9�3�װM���a���n��s��Xn�a���L�T�2�����~��b��A���Xi��d�����ؽ�-�a	���־M�!���i�롿=׿�	�؝+��8Q�8z��ɑ�?���گ��   �   ����0��s0��K���j���]�R�4������ߴ����v�ز*�>���;����3��Eڽ\�����=���,�g6J��ك�������ٽ���o��5&�0��N3���/�qw%������6�ֽ�੽�6����D��'�pY8��;��6׽@-2�|��U`�r�)��eu�[⩿/�� ~�BH4�f�\��ڄ�����w(���3���   �   ���±�ۂ���f���}�\�S�&�-����Fڿ�Z���\m�2@$�2Oھ����o�,���ν=�x���%�l�� �#�H�V��͍��b���qڽ|D���\�ެ��K����
�n����4ֽO����݈��gL��������j�Kn�>
ɽ�*)�F���a�׾�"�a.k��񢿟ؿԡ
�\�,�:�R��%|�;���b��[����   �   ���g���$ˡ��6���	x���O�X�*��x	���ֿ�����ni���!�u�־������*�X#Ͻ~���o3�s#��~?�+
z�^����nνW|����������&���)��	&��3�f�����ɽ��M�o��85�87��)��@u�"Zɽ�y'�h���:FԾ:���\g��]���(տ�����)�z�N�FFw�]������I­��   �   �@��rJ��5J���A����i�jE�Ƙ"����̿���^�����̾�̓�j�%�(XнH*���]�3+b�}D��>���罢l���*�C�mV�l b��e��Ia�D�T�d�@�C(�V��ޑ��'��w��W��BS�����r�ʽ��"�����&Mʾ.��B\�	ۘ��m˿�P���!�puD���i��J��p���k���   �   ˔�HR���ڇ��Nt�|�T��4�,�� ��ύ��6L�F�[Ƽ���u����bԽ�c������
���I7Խ#s	�U�.��OV��}�F͏�b��O����Ĩ��v��Wj��灎�3z��+S���+�js���νI���~��n���Ͻ���$�r��[*�#�J�@��#��{A� ��f�4��U�j�t�(4��a����   �   �{���M{��l���U�p<�>� ���l�ؿ�Ĩ���|�֦5�����	1��o=`�x�~�ܽ6ʾ�>�ʽ�q���!�r�P�T���� �J��mN־�,꾞��� ������H�辶�Ծ�-���Ӟ�p偾A?M�"����ŽD#��Q9ؽ�����]��̧���}�4���{��j��asؿ6/�rS!���<�p�V��m���{��   �   �EX�x�S��H���6� �!��a����j���-ϑ�M�Y�HM��.پǷ��'�I����H�"�Z���3���l��ƙ��������p
����e�*��4�f7�)�3��*�}���3	��r����@˗�K�i��1�����罢d�����G��ʒ�zFؾ?��iY�	ؑ�����n���F�"���7��I��}T��   �   �2��\/�>W&�*��Z������ÿ0Q���rs�k45��-����M�|��94�u���:�r����=���|��i���۾��	�9�'�lfD�,�]�K�q��C~�,+��e�}���p�yM\�C�B�&�R��,�ؾ����� z�Y;�����&L�:3�ʊ{�Tµ��&�Jj5�
t�-ꝿ5�Ŀ��������='���/��   �   ����[�\R�����ݿ(���잿-�~�":D�����'Ҿ�Ô�e�T��h"�����8�L"=���}�����,o�����=���e�X<���9��<q������m��eH��i���1��n(����c���;��d��o�� ���e{��;���l0�I�!�P�T�b锾*�Ҿ�U��E�����������#�߿���R�l���   �   �E��8Ὺֿ{�Ŀ� ��`���y���F�߬������&�m���2�b��o���3��o�,����a侀��$H���z�ؙ��T���0Rƿ�?׿G��}I�U<� ֿ��Ŀ�#��mb���y��F�_��o㾑���d n�<�2�Ѓ�����3���n�O����]�Į��H�r�z�G���d����Nƿ(<׿����   �   �i��AE��o���F.���%����c�O�;��a�jk����:a{�<�;�_�X0�x�!��T��딾l�Ҿ
X��"E�N��4���ϑ��W�߿����@�p������]�:T������ݿ�*�����~��<D�����*Ҿ�Ŕ���T��i"�B���6�0=��{}�=����j���ȏ=�:�e��9��7��-n��y����   �   }(��$�}���p��H\�4�B��&�u����ؾF�����y��U;�	�ת�hL��3���{��ĵ�k(��l5�Et�8읿��Ŀ�쿂�����@'��/�0�2��^/�HY&�������I��a�ÿ	S���us��65�c/������|��:4�O��o9�����=��|�:f��۾��	���'�/bD�s�]�2�q�f>~��   �   )�6��3��*����0	�pm龭����Ǘ���i� 1�{����罗c�N����G�̒��Hؾ	���kY��ّ��
��Gq�\���"���7�!I�j�T�*HX���S�!H���6���!��b����3����Б�m�Y��N�1پ����O�I����?F�b�W�L�3���l�Ù�8���V�뾈m
�ܦ�d�*�R	4��   �   ����������l�ԾF)���Ϟ�*⁾:M�'��I��0�Ž!���8ؽ���S�]�$Χ�l��/�4�;�{�l��=uؿZ0��T!���<�|�V�,m�,�{�,}��dP{�>l���U�<��� ����ؿ�Ũ���|�5�5�v���)2���>`���S�ܽxǾ�ȂʽQk��<!��P�ܼ��ƾ��q���H־'�o����   �   v���^r��bf��I~���z�&S�|+��o� �νE��|���l���Ͻ_����r��ﺾb+���J�=��h��C������4�\U�P�t�D5������C̔�wS���ۇ�BPt���T��4���r	�＿�Ѝ�8L��F�HǼ���u����Խb��p���{���:1Խ=o	���.��IV�	}��ɏ�^������   �   ��e��Da�e�T���@�?(����A��N#����W��?S������ʽ&�"�=���5Nʾ�.�D\��ۘ��n˿~Q���!�dvD���i�gK���p���l��xA��\K��K��nB����i�4E�^�"�z�_�̿+򙿈^�����̾�̓���%��Wн�(��Z{]�W%b��@��M��� 	�
i���*�rC�qV�5b��   �   "�)��&�51�K�����ɽ���%�o��55�
5��)�'@u�nZɽDz'�֯���FԾ����]g�=^���)տ ��D�)��N��Fw����)����­�����伭��ˡ�L7��:
x�*�O���*��x	�6�ֿ񰡿1oi���!���־������*��"Ͻ����m3�p#��z?�=z�^���"kνYx�����Q��H�&��   �   �K����
������4ֽu���ވ��gL������.k��n��
ɽ�*)�v�����׾��"��.k����ؿ�
�t�,�T�R�&|�J���b��b������±�Ђ���f���}�B�S��-�j���Eڿ�Z���\m�@$��Nھ����/�,�D�ν��x�.�%�����#��V�o͍�ob���qڽeD���\�ج��   �   &�)��&�:1�N�����ɽ�����o�T55�~4��)��>u�zYɽ{y'�:����EԾ���\g��]���(տx����)� �N��Ew���?�����������ử��ʡ�6���x�4�O���*�\x	�V�ֿF���2ni��!���־�����*��!Ͻ����l3��o#��z?�z�T���kνQx�����T��K�&��   �   ��e��Da�n�T���@�?(����*��&#����W�K>S�������ʽ��"����nLʾ�-�>B\��ژ�m˿xP�P�!��tD���i��I��Go���j���?��I��RI���@��`�i�nE��"�j���̿�𙿢^�)��Ʌ̾�̃��%��Uн�'���y]�N$b�?@��������h���*�sC�vV�>b��   �   |���dr��if��N~���z�&S�|+��o���νpD���z��k���νI��{�r�l��)��J�~��%��5@�0��X�4�rU���t�3��5����ɔ�Q���ه��Lt���T�ƴ4�,����V��΍�j5L��D��ļ���u�Ⱥ��ԽF`��N���đ���0Խo	�p�.��IV�}��ɏ�^������   �   ����������u�ԾK)���Ϟ�&⁾�9M���������Ž���5ؽ)��|�]�8˧����4��{�Ti���qؿ:.�4R!�d�<���V���l��{��z��HK{��l���U��	<��� �����ؿè�A�|��5����2/���:`�(��ܽVž�o�ʽvj���!���P�Ѽ������p�� I־'�w����   �   0�6�	�3��*����0	�rm龪����Ǘ���i���0����o��$`齚����G��Ȓ�ADؾ����fY��֑�����l鿔���"���7��I��{T�$CX��S��H���6�F�!�0`���c����͑�˥Y�kK�I,پε���I�����B��LV���3���l���+���M�뾆m
�ݦ�g�*�V	4��   �   �(��*�}���p��H\�:�B��&�t����ؾ-���x�y��T;������I��3�a�{����%�h5�'
t�W蝿�ĿM�<��*���;'���/���2�hZ/�(U&�F�������꿥�ÿ'O���os��15�,���D~|�X64�����7����)�=���|�f���۾��	���'�.bD�t�]�5�q�j>~��   �   �i��DE��r���I.���%����c�O�;��a�Sk徜���`{�1�;����-�w�!��T�"甾�Ҿ�S�E�$������a����߿����r�p������Y�tP���U�ݿG%��IꞿK�~�7D�I��M$Ҿ0���u�T�ze"����5�=� {}����jj�����=�6�e��9��7��0n��{����   �   �E��8΅ֿ��Ŀ� ��`���y���F�֬���÷��;�m� �2���ʪ�X3���n�����Y�8��W	H�c�z�ٔ���~���Kƿ�8׿��1B�*5�8ֿF�Ŀ��y]��@�x�$�F�����䴤�m�m�ˑ2�&��.��3���n����x]侷���H�n�z�F���d����Nƿ+<׿����   �   ����[�^R������ݿ(���잿.�~�:D�����'ҾbÔ��T��f"�����3�q=��v}�����(f�E��@�=���e�S7��Y4��3k��X����f��B��i���w+��t#���c���;��^��f�5���[{��;���<-�.�!���T��蔾�Ҿ�U��E�����������$�߿	���R�n���   �   �2��\/�BW&�.��\������ÿ1Q���rs�c45��-�u��?�|��74�Ο��6������=���|��b��k۾��	��'�^D���]�4�q�&9~��%��ޏ}��{p�:D\��B��&�p����ؾu�����y�Q;�p�Ч�I�{3���{������&�>j5�t�+ꝿ3�Ŀ��������='���/��   �   �EX�z�S��H���6� �!��a����j���-ϑ�H�Y�;M��.پ_���ɇI�z���A��뽭S���3�/�l�f����������Wj
�B��x�*�.4���6�܋3��*�?��Q-	��g� ����×���i�\�0�������\^齪����G�ʒ�9Fؾ.��iY�ؑ�����n���F�"���7��I��}T��   �   �{���M{��l���U�t<�>� ���o�ؿ�Ĩ���|�Φ5�s����0��g<`�����ܽCþ��}ʽ�d���!�|�P�������������C־Q!�V�������r	������Ծ{$���˞��ށ�q4M����1�򽅄Ž\���4ؽ^����]�Ŗ����r�4���{��j��asؿ8/�pS!���<�p�V��m���{��   �   ˔�IR���ڇ��Nt�|�T��4�.��#��ύ��6L��E�'Ƽ�<�u�����Խ�^����������2+Խyk	��.�qDV��}��ŏ�Z����5���-n��bb���z��:z�a S�Hw+��k���ν�?���w��i��P�ν���h�r�RL*��J�?��$��|A� ��f�4��U�j�t�(4��b����   �   �@��sJ��5J���A����i�lE�Ș"����̿���^����߆̾r̓���%��Uн'���v]�Gb��<������9罗e���*���B��V�b���e��?a�x~T�`�@�;(�b��4��@���ꄽC�W�%:S���2�ʽĽ"�^���Mʾ.��B\�ۘ��m˿�P���!�ruD���i��J��p���k���   �   ���h���$ˡ��6���	x���O�X�*��x	���ֿ�����ni���!�f�־w���>�*�:"ϽO��rk3�Jm#�bw?�� z������gν�t��p����߾&���)�&��.��!��G�ɽ"���
�o�u15��1��)�i=u�Yɽpy'�K���+FԾ7���\g��]���(տ�����)�z�N�FFw�\������I­��   �   ���Ü�AK�����T!c���?� ��H �ȿ�k����X����qǾak����>N����`����0����$���@�[���ܣ���ƽ��a���,y�'��r�1���e�9���j���p��Y0��5�(�ۼ��O�L#��8����y��ľA���3V�
���mƿ�����p�@�>��b�����++�������   �   ���M��m#��)]��8�^�ؠ<�h)����C�Ŀ�����HU�,|� 1ľ��{�z��{}���$g�,� �<���+��a�����`ֻ��p��T�a��H��v����ʦ�$��x�۽@;��6e����P�\���� �6x���U��w����v�����xp�=�R�;^��;�¿����h��Ѝ;��^�'��1���S���   �   $��쌏��E���q��R��"3����Z8𿘏���Ό��J��7�Һ�)�p��d�`���ѷ{��VG��K�1z��3��d�ҽH��I��2�HoC��IN�+�Q�xM�53A�]/��7�����ʽ΋����h���:�l�6���j����������k��ַ��l
�$�H��~��m
�������� �2��mR�n�q�_m��L����   �   3��C���r��[���@�^�$�4<	���ݿ���������o:�W� �f��%�`�b������rq������n��Y1��1������b�C��Fg��^��T���Ru���♾_���X`������Tc��O?����_��F\�����t�z����������;\��驾.
��v�8����������ܿ��ĺ$�0A��0\��Ys������   �   Rf��{a�d�T���A��)+�L�Z����^ƿ�X����f�C�%�v���w����L�E�	���Ƚ�F��N"���j����>���p������þn�վ��"��m7�Ծ�y���/��@D��O�k���9�{���ٽ�T���������\O��'I�򒘾`��,�$�;�e��왿q/ƿ����&���+���B�6�U��b��   �   ��C���?�\�5��&����6.��{տB���z.����F�߇��ƾ�̆��7������׽��ֽ��W;$���X��������Ȁ׾����M�y�]D$���&�s�#����֗�l���CԾe���Ή�~�S�� �/���F<н,�ѽ-�75�����k�ľ���BF��8��R��r�տ�R �����'���6�ޕ@��   �   #��  �0��������۰ֿ�粿���'^�*%�@J��� @f��;$��� �u�𽒴�3-��g��ޙ��$Ⱦ�����kb3�ˡJ�Y�\�t8h���k�=jg��T[���H�RT1����l���ž�Q����b�(�)�A��+������!�"���d������6�l%���^�g������cؿ���b������� ��   �   ̽�LW�Q���C��˿翮�#���#h���2����3m������*�A�2��x�5�
��v,��fg�=����PӾC�	�q$-�f�Q�_vu�U���u������u��׀��cx�������r��O��+�@���оq���]od�B*������ ���ܐA�J������v�2�3���i��]��h��g�̿�u��@���   �   !
ҿz<ο��ÿ���)����7����b���4��
���ξ�镾��X��M"����F�#���Y�o��dfо�D���6�^e�᱊�ۣ��·���Eſ�ο~ҿ�?ο��ÿ��������9��~�b���4�e�
���ξ?앾��X��O"�:����#�4�Y�����bоBB�K�6�Ze�����'���ô���Bſ��ο�   �   �r���}���u��$���r�&�O��+�����о����pkd��?*�v���� ���9�A�B���	���x���3��i�`���j��ZͿZ濠x�������Y�����c俏˿O®�)���&h��2�����o��\����A�������
��s,�Vbg� ���LLӾ��	�!-�P�Q��qu�eR���r���
���   �   ��k�keg�$P[�~�H��P1���Ig��hžN���b��)�W��|��>���z�"�9�d������9��n%���^��h��7��Wfؿ���������� �
#�� ���X�����Y�ֿ�鲿�����^��+%�	M�l��)Bf��<$��� �"��Q���-��g�ۙ�L Ⱦd�����^3�v�J���\��3h��   �   ��&���#�A���������>ԾZ
���ˉ���S� �N���j9н1�ѽ�-��85������ľ��.EF� :��*����տ7T ��T�'���6���@���C���?�D�5���&����0���տ鸫��/����F�B���ƾΆ��7����N�׽i�ֽ���h7$�X�X�:�������{׾�������	��@$��   �   n���1��Ծ�t��l+���@��U�k�0�9�_w�X�ٽ\Q�����g����O�e)I�O�����㾷�$�V�e�H$1ƿ����b����+�N�B�6�U�� b�@Tf�~a�R�T�D�A�F++�n�2���%`ƿ�Y��I�f���%�&���x����L�|�	���Ƚ4D��2��e���>�.�p�쒾����"�þ�վ7��   �   ߙ������\��k����c��J?�������*W��H�����z��������4���\��ꩾ����8���������y�ܿ���ػ$��	A�R2\��[s�����4��D��ܟr���[��@�T�$��<	���ݿ���������p:�� ��f���`��������o������B���+�����3��#�C��@g�1[������vq���   �   X�Q��M��.A�D /��3������ɽ������h��:�p�6�.�j�
��������k�z׷�Nm
�,�H�Q��M�����j���2��nR���q�n�������������F��&�q�̸R�v#3�"��-9�<��� ό���J�e8��Һ���p�e�䌽�b�{�$SG���K��)z�d/��لҽ������2��jC�9EN��   �   �s�������J���۽J8���b����P�k��~� ��v�x�U��w��\��v�T����p��R��^����¿x������N�;��^�b'�����OT������M���#��t]����^�,�<��)������Ŀ�����HU�U|�M1ľة{�s��}��B#g�� �l��A�+���a�ނ�� ӻ�Tm��R�0�� ���   �   &��r�C��f�9���j��+�p�.Z0�F6���ۼv���O��#��t���y��ľj���3V�*����ƿ����p�X�>��b�����4+���������Ü�8K��u��:!c���?���4 ��ȿ�k����X�����qǾk�����M��<�`�B��x����$�U�@��Z���ܣ���ƽ���N���&y��   �   �s�������N���۽K8���b����P�!��� �:v�N�U��v�����v�{���Mp���R�^����¿���.����;��^��&�����sS�����M�� #���\����^�V�<� )������ĿW����GU��{�o0ľ��{����|���!g�L� �����+�I�a�̂��ӻ�Mm��R�2�����   �   _�Q��M��.A�L /��3������ɽ�����h�+�:��6���j�M�&����k��շ�l
�z�H�,~���	��˓�>��x�2� mR�V�q��l������T����� E����q�ֶR��!3���<7𿲎���͌���J�,7��к���p��c������{��QG�w�K�F)z�(/����ҽ���v���2��jC�?EN��   �   ߙ������\��p����c��J?��������V��������z�6���&���J���\��詾���r�8����������ܿL��ع$�A�B/\��Ws������1�� B��8�r�r�[�Z�@�D�$�N;	�;�ݿ�������zn:�U� ��d����`����{����m���������F+���������C��@g�/[������yq���   �   t���1��Ծ�t��p+���@��L�k��9�-w���ٽ8P��4�x����M��%I���������$�~�e��뙿�-ƿ���
����+��B�L�U�|b��Of��ya�d�T�؟A�f(+�
�A����\ƿcW��^�f���%�"��=v���L��	���Ƚ0B�����2d�����>��p�쒾����"�þ�վ=��   �   ��&���#�E���������>ԾV
��yˉ�d�S��  ����d7н��ѽ+��45�6���b�ľx��@F�?7�����q�տ�Q � ��'���6�ʓ@�\�C���?�d�5�~&�"���+��<տe����,��r�F�+��bƾˆ�/�7�$����׽5�ֽ0���6$�	�X�"���{���{׾�������	��@$��   �   ��k�qeg�*P[���H��P1���Gg��^žgN����b�d�)�P��@��4�����"�m�d�i����3�j%���^�Se�����-aؿ������$���� �#����T�� �����1�ֿD岿#���*^��'%��F���J<f��8$�:� ����4���-�Lg��ڙ�4 ȾS�����^3�u�J���\��3h��   �   �r���}���u��'�� �r�)�O��+����	�оq����jd��>*����5� �����A�8���A���t���3�@�i��[���e����̿� 濯q��r����zU�������˿W�������h���2����j��I�����A�!�����
��r,��ag�ꓝ�(LӾy�	�� -�J�Q��qu�eR���r���
���   �   $
ҿ}<ο��ÿ���+����7����b���4��
���ξ�镾��X��L"������#�U�Y�>��1_о�?�J�6�KVe�H�������౵��?ſl�ο�ҿ+9ο��ÿ���~���\5����b���4���
�ʝξ畾5}X�xJ"����@��#�?�Y�����bо3B�B�6� Ze�����&���Ĵ���Bſ��ο�   �   ̽�NW�U���H��˿鿮�#���#h���2�����l��K�����A�F����ؐ
�qp,��]g����JHӾ�	��-�h�Q�"mu��O��p������o��{���r�����v�r��O�^+����ԥоT���{fd��;*�N���� �����A�⹇�����v�'�3���i��]��h��f�̿�u��B���   �   #��  �2�����#���ݰֿ�粿���%^��)%�J�M��?f�V:$�}� �$��P���-��g��י�Ⱦ���l��Z3�@�J��\��.h��k��`g��K[�8�H��L1�K��a���žK����b�ح)����������}�"���d�2����6�l%���^� g������cؿ���d������� ��   �   ��C���?�^�5��&����:.��~տD���{.����F�ԇ��ƾ�̆���7�����׽l�ֽe��d3$�!�X�鈌�i���v׾���� �:��<$���&�ޤ#����<�������8Ծ��ȉ��S���������3нS�ѽ+��55�H���*�ľ���BF��8��O��p�տ�R �����'���6�ޕ@��   �   
Rf��{a�h�T���A��)+�N�\����^ƿ�X����f�;�%�P�徥w����L���	�k�ȽD@��\���^�"��>��p�^蒾\���J�þűվ��¬�D,ྊԾ�o��'���<��	�k��9�>s���ٽL���諒V����M��&I�����2���$�5�e��왿p/ƿ����$���+���B�8�U��b��   �   3��C���r��[���@�`�$�6<	���ݿ���������o:�K� ��e��x�`�J��z����l��-����	��0&��������C��:g��W������m��&ۙ�����Y�����| c�RE?�<�����FQ��������z�g��n���|���\�^驾
��n�8����������ܿ��ĺ$�0A��0\��Ys������   �   #��팏��E���q��R��"3����[8𿙏���Ό��J��7��Ѻ���p�7d�B�����{��NG��K��"z��*��xҽ�������2�BfC��@N���Q�
M�?*A��.�/0�^���*�ɽ�����h�̨:�7�6���j���A��E�k�aַ��l
� �H��~��m
������ �2��mR�p�q�`m��M����   �   ���M��n#��*]��8�^�ؠ<�j)����D�Ŀ�����HU�*|�1ľ��{�$��p|���!g�� ������+�`�a�^���&л��i��P�������q�V�����B
��m�۽5��	`��I�P����F� �2t���U��v�����v�����tp�;�R�:^��:�¿����h��Ѝ;��^�'��2���S���   �   ��_ ���y�γa���E���(�8���/�xD��e��S?��=���ja���
��ꤽ�GB� ���t/ּ�����&�!�^�f쎽㭽�?ɽvf޽}T뽹�p轖�ؽ�Y��l������n�E�?���������H2ļ��&�������K�Y�漫�����g<��/��3��v���X���'�<�D�*-a�ވy�c���   �   �E��ud����t��s]��OB��&��N
��߿f�������<�7�t��/^� b	�f
��HH��	����l*�seC��i��)N��f}ƽ������}5�&-����g���ܽ�����Ԙ�|�i��(���������5ۼR�,�@t���t�8�V�����Z��mW9����]z��sqݿ�:	�v%�D�A��]�L�t�j���   �    �z�`ku�V�f��sQ��i8���V��dտ��ɺx��2�p0���¤��wT�~?��ܥ�h>Z��+�p�/��5Y���������#0	������+�X[5��8���3�h�(�n��J���Kڽ>F��' >���h���@�B���X���8�M������0o0���u�R���7xӿ���&)8���Q�^g���u��   �   ��c���^��4R�p�?�F})���g󿗝Ŀ� ����d�uP$��C�y���[�E����������{���g� ���@J��H�ܽ����,�	�K��g�=}�m[��t_��nx����y�M�b��VF��v&�!���)Ͻ�꛽#�n���N�Q�b�|ߜ�1
�#@��锾\�߾��"���b�C��ӽÿ��򿔵���)��,@���R��K_��   �   p_H�tqD���9��<*��9��a���ٿ#���,]��vK����&>ʾ���?4�6��Fz��
��ᠽԫƽ�~��<(��T�t���sc�����}W���?ƾ�Kɾ�1ž�[���ة��3��)y|� �M��W!�����-*����� 
�������Tt/�����=�Ǿ���\J��*z���	ڿv�����P)+��:���D��   �   ,���(��4 ��6����E�	����ї���j���.�����dj��sSm�ݚ!��=�Ʃ���Ի���޽����>��x�M�����X�޾�$��ρ	���� �����G�(����2۾(/��y��x�p��p8�Z�
��<Խ�4��P���Q_߽��j�����:���6�.��k�%0�������㿲��O��0!�m)��   �   E����j��S���ޯܿC,��P3��&�}���C�)W��о7	��v^J�v�(��[vҽK���A��K�\���^���C޾��)-�l�2��B�1�L���O���K��)A��0������9ھ�Ŭ�y��F���=���˽K�۽���)�H����S�о���eD�P�b��-׿���޿M�������,��   �   �|�m3��ۿ�ʿy���?u��P��0uL��F�5��<?��in���)�>6�����vq�K�K��䊾(I��ܢ�@��3>9�V�X��at��������^ҍ��%��6���q���U���6�RL�5���d����G��i�����߽C= ���)���n����뾴���QN��S���"������̿RݿF��   �   '��E����s���?��AF����q��G��	�Q8���v��5�����=���D�콜\�@��p�?�� ������.���	!�'`J��
u�\���O⠿&Į�l��)!��7����v��2B���H����q�K�G�)�Y<���y��D���:�=���� ��O[���k�?�@���ې��**��!��\J��u��􎿤ߠ�H���i���   �   �ύ�V#������^�q���U���6��I�������a��<�G�tg����h�߽4> ���)�3�n�A
���	�+���TN��U���$�������̿&Uݿ� �.�뿡6��ۿ�ʿ�³�fw����xL��H���龌A��nn���)��6�2�F���n�s�K�1⊾rE��	��=���:9�(�X��\t�-��������   �   v�O�x�K��%A�P�0�p������پU¬�Bv���F�4�����f�˽��۽���H����� �оݢ�}hD���d���ٿ�f�޿X���:��>.��F�@�����9���o�ܿ|.��/5��,�}��C��X���о�
��``J�P���TtҽF��>���K�\���w���$>޾� ��)���2���B���L��   �   ������D�b����-۾�*���u����p��l8�)�
�28Խ(2��i���`߽	��j��������3�.�tk��1��������PQ�T2!��n)��,�>�(�r6 �p8� ��G��¼�zӗ�%�j�]�.�4���l��hUm�қ!��=�`����ѻ���޽�����>��x�QI��d���޾���~	�P���   �   �Fɾ�,ž>W���ԩ��/���r|���M��S!����`%�����2��j���转u/�ļ���ǾE���]J���{��bڿ���6���*+���:�RE�:aH�,sD�\�9�:>*�,;��b�i�ٿz���8^���wK�����?ʾ���@4����Wy�����sݠ���ƽt{�18(�h�T�����_�������R���:ƾ�   �   \��u����y�x�b�dQF�_r&�o���#Ͻ/曽s�n���N��b�nߜ�K�b@��ꔾ �߾Ӂ"�0�b�L���ÿS�򿂶��)�.@�d�R�hM_�P�c�t�^��5R���?�J~)����_h󿭞Ŀ����d�\Q$��D�8���!�E��������w{���g�l���JE���ܽ���H�,���K��g��6}�X���   �   P
8���3�t�(�̀���DFڽ�髽jB��r>������W@�h���T���>�M������p0���u����,yӿ��΁��)8���Q��g��u�H�z��lu�l�f��tQ�Pj8�(����տ�����x���2�<1��dä�2xT��?��ܥ�E<Z�q�+���/�q/Y�
���������,	������+�W5��   �   +����c����ܽ����*Ҙ��i���(�D�����x3ۼ��,��t��u��V�; ���Z���W9�\���z��rݿ
;	��%�A�D]���t�qj���E���d��l�t�Dt]��OB�B&�(O
�D�߿@f��*����<�\����O^��a	�
��H��	� ���&'�aaC�5g��DK��$zƽ�����x3��   �   ��p车�ؽ�Y�����׋����E�z������ ���3ļ
�&��������Y��������g<��/��?3������X���'�R�D�>-a��y�f����[ ���y���a���E�t�(�$���/�WD��H񄿸S?�}=��𯾏ja�K�
�~ꤽGB�,����.ּ ���a&���^�G쎽�⭽�?ɽef޽qT��   �   +����c����ܽ���&Ҙ��i�}�(�̟� ���2ۼ��,��s��pt��V�|����Y��4W9����%z��)qݿ�:	�4%��A�>]���t��i��'E��d��,�t�4s]� OB��&��N
�Z�߿�e������!<������C^�Ka	�2	���H��	�����&�aC�g��4K��zƽ
�����y3��   �   T
8���3�{�(�Ҁ���?Fڽ�髽DB���>���q��N@���������Z�M�H����n0���u�ƈ���wӿ�����r(8���Q�Pg�t�u���z�ju�(�f��rQ��h8������cտ<����x��2�/������9vT�R>��ڥ��9Z��+���/��.Y�ƕ��ܯ���潺,	������+�!W5��   �   \��u����y�~�b�gQF�Zr&�f��u#Ͻ�国Z�n�ϕN�;�b�5ݜ����@��蔾�߾�"�Y�b�r��ɼÿ{��ȴ���)��+@���R�>J_�
�c�F�^�3R��?�$|)���me�E�Ŀ�����d�9O$��A�0���j�E�Y�������>{���g������D����ܽ���0�,���K��g��6}�X���   �   �Fɾ�,žDW���ԩ��/���r|���M�pS!������$�����������~ 轊r/�h�����Ǿ����ZJ��퇿�x���ڿ~������'+���:���D��]H��oD�$�9�`;*��8��`���ٿ�����[��3tK�)��<ʾf���<4�N��vv�����0ܠ���ƽ*{��7(�C�T�����_�������R���:ƾ�   �   ������D�j����-۾�*���u����p�bl8�Ԣ
�7ԽQ0�������[߽��fj���������~�.��k��.��Q���i��p�XN�/!�^k)�8,���(�*3 �x5�b�<C����TЗ�,�j���.�����0h��0Pm�M�!�9�<����ϻ�@�޽����>�fx�:I��S�� �޾����~	�Q���   �   z�O�~�K��%A�T�0�t������پK¬�,v���F�������x�˽�۽v��W�H��}����о ���cD�J�&`���Կ��޿g�������*�LC�ڟ�ȓ�Q���'�ܿ�)��H1��˔}��C�"U��о��"[J���1��"qҽ/���=��K�4���Z���>޾� ��)���2���B���L��   �   �ύ�Y#������c�q���U���6��I������\a����G��f����
�߽�: �ƙ)��n�'����n~��NN��Q��u �������̿�Nݿ迡y�40��ۿ�ʿཱི��r��_��rL�D�h��g<��.n���)�z3���:���m�ɳK��ኾLE����3���:9�$�X��\t�-��������   �   +��H����s���?��EF����q��G��	�C8���v������ǟ=�Ѿ�D�콊V�����?���������	&��f!�NYJ��u���ݠ�{���-f��)��Q���	q���<���C����q���G����3��Us��������=����̤�W�����?���������*��!��\J��u��􎿢ߠ�I���i���   �   �|�q3��ۿ�ʿ}���Au��P��/uL�{F���?���n���)��4���,���k�b�K�}ߊ��A��q��^�� 79�!�X�zXt����͍�� ��KŽq�s�U� �6��F���R���^����G� d����(�߽r; �j�)���n�j���뾦���QN��S���"������̿RݿG��   �   E����j��W����ܿE,��R3��&�}���C� W���о����]J������oҽ���4;��K�m�������r9޾���l&�ڪ2���B���L��O�.�K��!A���0���4����پj���,s��7F�y�����P�˽��۽:��+�H�f�� �о֠��eD�G��a��*׿���޿M�������,��   �   ,���(��4 ��6����E�
��� җ���j���.�����1j���Rm���!�:�u���^ͻ��޽��N�>��x��E�������޾.��h{	����-��3�jA������(۾P&���q����p��g8�X�
�"2Խ0-���󳽤[߽��Gj�d������,�.��k�"0�������㿰��O��0!�m)��   �   r_H�tqD���9��<*� :��a���ٿ%���-]��vK����>ʾ���1>4�q��"v��/��٠���ƽ�w��3(��T�Ԧ���[��_���N���5ƾ�Aɾ�'ž�R��9Щ��+��l|�#�M��N!����������0������ �hs/�H����Ǿ���\J��(z���	ڿt�����P)+��:���D��   �   ��c���^��4R�p�?�F})���g󿙝Ŀ� ����d�rP$�qC�K�����E���������%{�U�g�e���<@����ܽ؏���,�e�K�4�g�/0}��T���X���q��!�y���b�LF��m&����*Ͻ������n���N���b��ܜ�1�{@��锾=�߾��"���b�A��ӽÿ��򿔵���)��,@���R��K_��   �    �z�dku�X�f��sQ��i8���X��cտ��ɺx��2�c0���¤�NwT��>�ۥ��8Z�V�+�w�/��(Y����>���8�~)	�S����+��R5�8���3�v�(�}����k@ڽ�䫽>>���>�N�����#@�X������жM������+o0���u�P���5xӿ���&)8���Q�`g���u��   �   �E��vd����t��s]��OB��&��N
��߿f�������<�4�h���^��a	�w	���H��	�\���"$��]C��d���H��wƽ���1���1�)���"`���ܽ=���PϘ�0�i�s�(�H��D���t.ۼ��,�Ts��et��V�����Z��jW9����\z��tqݿ�:	�v%�D�A��]�L�t�j���   �   ��`���\�T&P���=�� (���lQ��¿s���+�b���"�?O����I�@�X]����ԕ$��vӼ,S��|�м>4��v<�n�q������驽<m����ŽȽ����*b��X5����)9N��U������k�@�-�0�o��	��Jn��ؽ׌6�����_�۾���&|_��ϕ�9����S����U'�zx=�P��\��   �   �\��pX�fgL�j�:�:%��.��z�	ɿ�z1��:_��6 �;�ݾa���h�=��꽝����d)����AмJ���x%���[��Y��57��K���r�Խy��c:㽃{ܽ��̽T׵��<��7s�o�3�b���\B����i� <����Go�T�ֽ$�3�X���_Mؾ�]�5�[��t�����޳뿮k�D�$�PR:��[L��yX��   �   ��P�r�L���A��>1��B�$}��X�&���N����T��?�q�Ҿn����^5�6I㽬����8���&g��g8�o�r��j��*ĽB��RA�<��ޮ������X��Ԥ���~ڽR`��ƹ���H�ڴ���м`�ʼP���<r��lн�J,����'�;���nQ�}����O���!�(����M1���A�ZM��   �   FK?���;�v�1�8#���8��-�п�p��ஂ���B����U���抁���(�V�ؽ�ꎽoT�� D�Pa�oV���}��xM�@��v.�\cE��W���b���e�V|`�<S��B?��[&�8�
��ܽ����v���7�J����-�m�y�m�ǽ� ��x{�������	�vA�ǁ�4����yп�(��fD�܇#�zU2�<��   �   *���&��}����`��v�߿yҺ�F��9�h��2-�e��S����g�.N��ͽO7��t�~��I���$���4ݽ}���5�
�]�k��M���[���������Lk������Ǐ�|�a�T��,,�����ɽB���Dl���\�x���
Ҿ������a�]`��R����,�
�g����������Y��h��/�f'��   �   �/�����V	�����L>Ὶ+¿��������%H�B��6Xվ�N����I��	��Ný%���:���4��Eu��r!#���S��u���)��!��b�־��o/��R���s����j�*Ӿ�����r�����yJ�u�RQ�	X���/��0��� ��7&�k�E������Ծ�i�L9H������[��7_ÿ"��R��� 
�.���   �   �����B�4��Կ�T���ע�� ���X�A^&�����P��M�w�r|+��2�f������.ɽ�c�͖-�,�g�r����z�������u-���%��a.��1��-�$>$�X��H���ྚ�������37_��&�z��㝽�wO��ε������@)��v��;��ۙ��&&'��zY�n6���R������ֿ&�迈&���   �   �*ʿ�uƿ���r.���˙��߃��Z���-����R4ƾ�����I�IQ�N
ٽr���̽�3 ��5-���l�񾞾��ξ��!����8�dcP�Q�b��vn�-r�>km�&�`�7�M�_�5��T���}=ʾ���Gf�L�'����.�Ž|ܹ��`ֽ���3@J�����j�ǾO����/�%�\��l��҈��X䮿�⽿?=ǿ�   �   �]���`��;[��Q��.�p���M���)����aϾa���ms^����:��ʘŽj�ƽ*���H"�`%b�B?��=jҾ�	�f,��P�]$t�����#������K`��lc���]���
�� �p��M���)����Ͼ齙��v^�K�����|�ŽT�ƽ4��LF"�|!b��<���fҾ~	�c,�h�P�7 t�e����������   �   �r��fm���`�\�M���5�#������9ʾ��Cf�I�'�I���=�ŽEܹ�3bֽ���#CJ�ɥ����Ǿg��[�/�~�\��n������殿�彿@ǿ�-ʿ�xƿN����0���͙��ჿ�!Z�;�-����$7ƾ������I��R�mٽoq���̽�1 �z2-��l�˻����ξ<��� �8�d_P��b�prn��   �   =1�c�-��:$�/
��E���ྯ�������g2_�&�$u������N���������B)�T�v�>��1���c('��}Y�/8���T�������ֿ���w)�������E�n7� �Կ8W���٢��"���X�G`&�����R���w�~+�4�B���b��8+ɽa��-��g�!���kv���
���1*�q�%�:^.��   �   ��������8e�CӾb���?o��ᝀ�uJ�����K�6T��n-��\��0��T'�~�E�[���.Ծ�k��;H������]��?aÿu������!
����@1�b���W	�T���{@�{-¿D���e����'H����OZվ9P��_�I�w	��Ný���������/��Zo��t#���S��r���%��� ��S�־꾯)���   �   ���g�����Gď���{��zT�?(,� �ޖɽ��?l���\�����Ҿ������a��a�������,� �g�<���������Z�j��0�xg'�|*��&�:�®�`��-�߿�Ӻ�)G���h�+4-��f�����!�g�O�&ͽ�6����~��F�� ���.ݽ���R�5�P}]�����
���W��{����   �   ��e��v`��6S��=?�\W&�h�
���ܽ����v���7�\����-�A�y�X�ǽ� �`z{�������	��A��ǁ�R���{п�*��RE��#��V2�B<��L?��;���1�0#���2:��W�п~q��������B����]�������=�(���ؽ|ꎽ�T���C��a�*R��<x���F�B~���-�9^E�V�W�ïb��   �   ��Y���������Jyڽ�[��������H�ӯ���м��ʼ,���<r��mн�K,�L��>�;����oQ�*����P���"���B�\N1���A�LM���P�\�L���A��?1�DC��}��Y�ɯ�������T� @� �Ҿل���^5�zI�V���3�8����b�Db8�l�r�Zf��Ľx��>����>���   �   �6�xܽ^�̽ZԵ�:��}2s���3�$����=���i��9��h���o���ֽ��3�ϰ��Nؾ!^���[�<u������u��l���$��R:�4\L�*zX���\�qX��gL�ƕ:�R:%��.�{�Nɿ��1���_��6 �z�ݾ������=���V����c)�ȋ漜=м�D��Gu%�t�[�jW��_4��,����Խ����   �   Ƚ����8b��d5�� ��Q9N��U�`�����k��-�|�o��
�rKn�x�ؽ�6�������۾���X|_��ϕ�Y����S�*���U'��x=�P��\���`���\�H&P���=�� (���LQ��¿W�����b���"�Oᾷ���@��\�P���t�$��uӼ�R����м�3�Bv<�6�q������驽0m����Ž�   �   �6�xܽb�̽WԵ�:��2s���3���� =��|�i��8��l��:o�׋ֽ��3�,���Mؾt]���[��t���������xk� �$��Q:�J[L�(yX���\�pX��fL���:��9%�@.�'z�ȿ�1���_�(6 �~�ݾڤ����=�ڵ꽊����b)�0�漈<м�C���t%�6�[�TW��N4��"����Խ����   �   ��Y���������Fyڽ�[������J�H�a��0�мX�ʼ_���9r��kнJ,���o�;����mQ����SO��!ῲ����L1��A�rM���P�~�L��A��=1��A��|��W�G��������T��>�D�Ҿ����=]5�*G������8�����a�oa8���r�f���ĽT��>����;���   �   ��e��v`��6S��=?�]W&�^�
���ܽk����v���7�����-�N�y�X�ǽ�� ��v{�f���+�	�dA�ZƁ�L����xп�'���C��#�dT2��<�J?�p�;�L�1�(#�
�)7����пfo�������B����ˀ��ȉ��ۯ(�{�ؽL莽�T�c�C�ia��Q���w��lF�~���-�'^E�N�W���b��   �   ��� g�����Jď���{��zT�4(,� ���ɽ���$=l���\�����LϾ�&����a��^��c����,�D�g����������X��g�F.��d'��*�F�&��|�f��J����߿�к��D���h�,1-��b������g�'L�Lͽ�3���~��E��2��I.ݽb��!�5�*}]�����
���W��{����   �   ��������>e�HӾc���=o��۝���tJ����.K�1S���+�����@���]$��E�$����Ծxh�T7H�G���oZ��\]ÿ��������
����J.�z��4U	�J����;῍)¿񜡿�����#H�����Uվ�L��֮I�]	��Jý��������.��^n��#�^�S��r���%��� ��I�־꾯)���   �   >1�e�-��:$�1
��E� �ྪ���}���?2_��&�t��2���~K�������콂>)�حv�9��Ж�� $'�-xY��4���P��S����ֿl�迨#������?��1��Կ�R���բ�3��X��[&�����0N��z�w��y+��-�����r��8)ɽf`���-���g�����Ov��o
���,*�p�%�9^.��   �   �r��fm���`�`�M���5�$������9ʾ�<Cf���'�������Žhع�`\ֽH���<J�l���}�Ǿ]��#�/��\��j�������ᮿ7ཿy:ǿ
(ʿ,sƿ}���+��]ə��݃�^Z��-����1ƾ@���l�I�kN�dٽLm���̽�0 ��1-���l�����b�ξ/�����8�`_P��b�orn��   �   �]���`��=[��S��2�p���M���)����RϾC���s^�G�����=�Ž�ƽZ��AC"�{b��9���bҾ5	�B`,���P�8t�(���9������[��O^���X�����p�$�M���)�Z���Ͼx���o^������Ž��ƽ���mE"�� b�M<��`fҾp	�c,�_�P�0 t�d����������   �   �*ʿ�uƿ���u.���˙��߃��Z���-����94ƾ����y�I�KP�2ٽTm��̽/ ��.-�_�l�������ξ� �����8��[P���b��mn�
r�Vbm���`�i�M�m�5��h����5ʾ뚾�>f�t�'�;���/�Ž�׹�L]ֽ���s?J�V���@�Ǿ?����/��\��l��Ј��W䮿�⽿?=ǿ�   �   �����B�4翃�Կ U���ע�� ���X�=^&�����P����w��{+��/�t���N��f&ɽ^��-���g�唖�cr����?���&���%��Z.�~ 1���-�.7$���C��ྉ���,���-_��&��n�������I���������@)���v��;������&'��zY�j6���R������ֿ'�迊&���   �   �/����V	�����O>῜+¿��������%H�>��Xվ�N���I��	�lKýv󞽔����*���h��e#���S��o��"��7���Z�־�	��#����������_�@Ӿ饹�dk�������oJ����"E��N��)��k��>���%���E�v����Ծ�i�A9H������[��6_ÿ!��P��� 
�0���   �   *���&��}����b��x�߿yҺ�F��9�h��2-��d��2���g�dM�Tͽ�3��.�~��B��*���(ݽ�����5��w]���������S��K���B
���b�����������{�2uT�p#,�&��r�ɽ����6l���\�ʉ���Ͼ�����a�.`��5����,��g����������Y��h��/�f'��   �   FK?���;�x�1�8#���8��-�п�p��ஂ���B����=������� �(���ؽZ莽� T���C��a��M���r��@�Rz�T�-�%YE��|W���b���e��p`�1S��8?��R&�h�
���ܽ�����v�&�7�(��2�-��y���ǽi� �,x{�`�����	�nA�ǁ�3����yп�(��fD�܇#�zU2�<��   �   ��P�r�L���A��>1��B�&}��X�(���O����T��?�d�ҾU���,^5�H�����/�8�h��d^��\8�i�r�$b��$�ý�{��:�W�����Y��������0���sڽwV��i���J�H�ة�Ƚм8�ʼq��&9r��kнfJ,�s���;����nQ�{����O���!�*����M1���A�ZM��   �   �\��pX�fgL�l�:�:%��.��z�	ɿ�z1��:_��6 �6�ݾV���@�=����Ȓ��Ub)�t��t9м4?���q%�}�[�U���1��$�����Խ���d3㽡tܽ�̽@ѵ�A7���-s�L�3�����7����i��5��H���o�Ëֽ��3�I���UMؾ�]�3�[��t�����߳뿮k�D�$�PR:��[L��yX��   �   ��6�^�3�:t*��z�B>�o9�Ņȿ񅡿��z�8�:��/���-�x�� ���ǽ�.p�9�ͥ�h߽�L~��p8"�yCL���t����x!��dI������,����=�s��-E��x�0����L�`S��`���p����!��Q+��6��FN��k�ࣳ�r���7��Kw�_ꟿKǿ���8�
��7�\*���3��   �   ��3�@�0���'�H���	��i�cPſ�䞿ZZv���7�����϶���t��<�jlŽ��o�$���ϼtN��8@޼ʤ��<���j�v(��!Ο��y��\����m���y���2��죍���h�t�1�*�������� c��`�߻(���=6,�ww���%��g�\����� ��4�^Zs�k����ÿN�h��J��К'��0��   �   �	+�f(�X��������Z�w����@��bJj�
�.�����Y�����h��
�����o�@;�������b� �f�P�h���֑��Zy½*�ܽL2��������ǆ��#�A�ʽ�`��Jʈ�O�K�ְ��İ�p�e��o\�x��-{/�����	�]��C��I��,�0�g�L"��.��µ��w������#(��   �   R�����"��\�>�qп�d���L���sW��b ��.����+aV�Q�!Ҵ�.fp�F4��(��(A��Pv�����Jʽ���p���`#�}�1��W:�N<��X7���+����R|���۽����~�U�2������3̼֭���6�r���s� ��DL�����⾭���U�z���g���пp��ʫ��y�D��   �   ����z
�t��sW�I�׿���Ě��%x��?�'h�CQ̾#ҍ�^?�ը�������v���U�W�e�濎�mF��n\�"��D8�t�W�Ks�4��^���M~��>���A��u�j�̲L�#�+���	�2�ӽҲ����`��T+�.+��JE��0����꽔b7�Yz��͏ɾ�R���>���w��������ؿ�h�%�^�
��   �   C����k𿹍俁Iҿ�*��w���C���w�U���$�ik���X����s�X�%�e὜���=��������$�ͽ�4�7�0���]��N��������q���btʾ�G;b�Ⱦ����r¬�=���h9��r�P�=#�'T��~����턽��Y�Y�]��\��/5ӽ�b ���o�����.�$�}@V��4��5񡿉j��O�ӿ���A��   �   wο�Kʿ�0��X���L蜿�����^���1�F��[�ʾ�����bK�:_�gtƽ$���ݐ����^bֽ&$��C@���y�M����ݽ�n޾w����p�.j�^��������&���ؾ0�#���um�o�4�x(��N½w�b���*l���L��GO	�	�I�fv���k˾�i	� 3�F�`��ڇ��Y��W��.b����ʿ�   �   j�������f5���N��/~��OY��R3����[۾�j��P�i��y$�����]��ߙ�f���iҽy�� �C� 7������U_־���
���+���:�HoD��eG�0{C��9�"+)�1@����æо�A��5�|��:��^���Žr6��]���={��Y��W�%�Fl��j���ݾ�����5��\����Ṑ�_U��R8���   �   y����3��c�t�H`��LF�<3)�bE�m)ݾ�x��f){�G5�6>�ܶ���蝽�l��U5ý���F%:��̀��f��[�����9,��8I�0�b�|�v�(������5��n�t��K`�'PF�6)��G�"-ݾi{���-{�>5�(@����W靽l���2ý���":�zʀ�{c��h��~��?,��5I�W�b�V�v������   �   bG�wC�p9��')�_=����̢оf>��[�|�l�:�<\�8�Ž�4�����~|��9�罾�%��l�.m��q�ݾ��J�5�\�ց�������W���:��̶������7���P���~�SY�QU3�����۾�l����i��{$�"���^���ޙ����fҽ���2�C��4��h���#[־�����B�+�;�:��kD��   �   I�����������x�ؾD﷾犖��om�q�4��%��J½�*���Pl���N���P	���I�Wx���n˾�k	�]3�2�`�x܇��[������d��!�ʿ�ο.Nʿ�2��u���-ꜿ@�����^��1���Ӹʾ@���/eK��`��uƽ����ې�<���^ֽ!��?@��y�騜��ٽ��޾����m�!g��   �   �B;��Ⱦ���h�������Z6��c�P�.	#��M��Ԛ��Bꄽ��Y���]��\�� 7ӽ�d ���o���������$��BV�O6����|l��x�ӿϹ忬����n���俏Kҿ�,�����������U�)�$��m��HZ��,t���%��f�����Z��x�������H�ͽ�1���0�o�]��K��l����������oʾ�   �   �z���:��P>��y�j��L���+� �	�ӽ���x�`�P+�g(��IE��1��r��6d7��{����ɾGT�q�>���w�E������ؿ�j�&�~�
����|
�~��UY���׿����Ś��'x���?�Ei��R̾3Ӎ�m_?�D���&����v���U�Q�e�:���~A��V�3��b?8���W�,s��0��亊��   �   3I<��S7�]�+�����x���۽����~���2�x���-̼&�뼼�6�,���O� �AFL���2!�Ѝ���U�k�������	п��񿢬��z�<�J�����#�Z]�?�п�e��WM���tW�pc ��/�^���EbV����Ҵ��ep��C4�((�`#A��Iv�B����ʽN�������\#��1��R:��   �   �~��̀�����ʽ/\��Bƈ���K�_��\���Ľe��g\�$v��M{/�����H�	�8]��D�������,�P�g�#�������fx��������$(��
+�(����4������[�"����A��3Kj���.�ҫ��췭�]�h��۞���o��9��������ߞ ���P�ހ�������t½�zܽ�,�ܗ���   �   k��w���/��h���]�h���1��#��^����(W���߻�󖼏6,��w��&���g�칰�
� ���4�[s�uk��}�ÿ�N뿺�����0�'�|�0��3���0���'����*	�9j쿱Pſ0垿�Zv���7����ж��t��<�plŽ5�o�`���ϼ�J���;޼��Z�;���j�&���˟�w��p����   �   ����.����X�s��-E�y�|��d�L�U��@��������"��tQ+��6��|N�c�k������ٵ7��Kw�zꟿfǿ���D�
��7�\*���3� �6�Z�3�2t*��z�6>�S9𿩅ȿ؅��d�z��:��/�����x��� �C�ǽh.p��8����̥��޽��}��88"�KCL�u�t����l!��\I���   �   �j��w���/��d���O�h���1�X#������pT����߻��I5,�w��[%���g�%���|� �ֻ4�Zs��j����ÿ�M�0������'���0�H�3�ܨ0�F�'�����	�Ci��Oſ�䞿�Yv�*�7�>��M϶���t�<�XkŽ��o�:���ϼ�I���:޼t���;�6�j��%��l˟�w��f����   �   �~��À�����ʽ'\��0ƈ�U�K�������,�e��c\�s���x/�ȣ����	�- ]�C��o~��z,�e�g��!��������^w�v��N��.#(�*	+��(���� ��v���YῘ���<@��6Ij�%�.�����^���7�h��	�ʜ���o��7��������ݝ �͏P�����\���Ot½�zܽk,�ʗ���   �   )I<��S7�X�+�����x���۽�����~��2�����(*̼��`�6���d� �mCL����D�ɋ���U�����u��qп�����x�V�\��&���!��[��<�п�c���K��1rW�Za ��,�9���I_V����ϴ�rap�
A4��(��!A�nHv�����Iʽ����|��x\#�ѷ1��R:��   �   �z���:��P>��z�j�|�L���+���	��~ӽ����r�`�qN+��%��EE�r.������`7�-y��1�ɾ�Q�:�>���w��횿$����ؿ�f�z$�F�
�����y
�b��rU�y�׿~��5Ú�z#x�E�?��f�>O̾�Ѝ��[?�S��������v�P�U���e�>����@��kU����)?8�ԂW�s��0��޺���   �   �B;��Ⱦ���h�������V6��Q�P�	#��M��A���V鄽ϚY�a�]��Y���1ӽ�` �G�o��|�󾊥$�a>V��3����h��D�ӿC��������Ri�h��WGҿ�(������˓���U���$��h��eV����s���%�(a��������������4�ͽ1���0�&�]��K��T����������oʾ�   �   H�����������x�ؾB﷾⊖��om�G�4�:%��I½f퓽纁��h��dI��$M	�@�I��t��li˾!h	��3���`�ه��W��;���_��C�ʿ�οPIʿL.��'���P朿㙆�$�^�S�1�a��z�ʾ[����_K��\�=pƽD���ِ�J����\ֽ� �$?@���y�Ĩ��yٽ��޾
����m�g��   �   bG��wC�q9��')�`=����Ƣо\>��4�|�+�:��[���Ž�2���񒽂w����罗%��	l�0h����ݾ����5��\�~��շ��'S���5�����^���$3���L��d~��LY��O3�J���۾�g��=�i��v$���轑Y���ڙ��
��9dҽ����C�\4��=��� [־�����<�+�8�:��kD��   �   z����3��f�t�H`��LF�<3)�aE�f)ݾ�x��.){��5��=�޴���坽Nh���.ý����:�<Ȁ��`�����!��e,�52I���b�D�v�ڽ��K����1��D�t�>D`�oIF�F0)��B�f%ݾfu���${��5�P;�"���u䝽�h���0ý���|!:�@ʀ�Oc��C��o��4,��5I�R�b�T�v������   �   k�������h5���N��2~��OY��R3����N۾�j����i�,y$�Կ�([���ڙ��	��Qaҽ���>�C��1��"���W־������+���:��gD�T^G��sC��
9��$)�q:������о�:���|�<�:��X��Žb0���:x��>�罙�%��l�qj����ݾ���x�5��\����߹��_U��Q8���   �   wο�Kʿ�0��\���N蜿�����^���1�A��I�ʾa���ibK��^�&rƽ����'ؐ�����Xֽ��I;@���y������ս��޾ш��k�d�2�������������ؾ(뷾y���Sjm���4�"�:E½Uꓽ<����h��dJ��dN	�k�I�0v���k˾�i	��3�<�`��ڇ��Y��W��-b����ʿ�   �   E����k𿼍促Iҿ�*��w���C���w�U��$�]k��wX����s���%�Bc�ݖ��:��扃�%�����ͽ.���0�'�]��H������y
��w����jʾ4>;��Ⱦ����C�������)3���P��#��F��%����儽�Y���]��Y��3ӽb �p�o���ӽ�"�$�t@V��4��2񡿇j��N�ӿ���B��   �   ����z
�v��vW�K�׿���Ě��%x��?�$h�6Q̾ҍ��]?�x��������v��U�g�e�𷎽)<��{O�5���:8��}W�s�h-��m���@w��(7�� ;��[{j��L�Њ+���	�bxӽ������`��H+�<"�DE��.�� ��b7�(z����ɾ�R���>���w��������ؿ�h�%�^�
��   �   T�����"��\� >�qп�d���L���sW��b ��.�k����`V����д��ap��?4�(�A�Bv�����
ʽ�{��П�UX#�O�1�N:�QD<��N7���+�S���t���۽	��vy~���2�����@"̼Ơ�>�6���� �bDL����v⾤���U�x���e���пo��ʫ��y�F��   �   �	+�h(�Z�����
���Z�x����@��`Jj�
�.����N���z�h�Q
�����(o�7�\������ٙ ���P�B}��i����o½vuܽ�&�֑��wx���z��佦�ʽMW������/�K���𱰼��e� Y\��o��x/�࣡�:�	�� ]��C��9��,�,�g�K"��+������w������#(��   �   ��3�B�0���'�J���	��i�ePſ�䞿[Zv���7�����϶���t��<��kŽ+�o�*��tϼ4G���6޼�����;�|�j��#���ȟ�Rt������h��t���,��ʞ����h�[�1�8����t���E����߻��4,��v��l%���g�R����� ��4�]Zs�
k����ÿN�h��J��Қ'��0��   �   >P�������G����P��N���䠿R ����G���k־�����J��n��j���4Z�A���ּ(t¼�kԼ<Y���x��}7���R�_0i��Kx��~��py�5�i��P��m-��O������1�� ú��;�<� �;+��`dӼr���޽x�7��q��wSϾܵ�w�D�ʯ�eǟ�?j���߿7t��^��~���   �   ��F��Ξ����o�ܿ77��VH���}��VD��V�9�Ҿv�� <G��?����|
Y�4��l��|�ӼDC�u}���.�_�O�=o��s���[���'��>+��\4��Fs��M��!�ަ������q»���:��;p�\;@�лfռ��o��x۽��4�*��B�˾[X���A�"�{�G���p���AܿÒ��L�����   �   �@	�����R ��8�jҿ9��}���L�q���:��	��9Ⱦ�����Q=����I���0V����f� ����~���pA��7m�fh�����%���<½��ȽB�ǽ�4��%,���Ϙ�K�{���@�՟��u��t
��n0� ��L��"mܼ��h�z�ѽ�O,�����K1¾�y�#r8���o�����Ĵ��<ҿ�I�|k ����   �   ���cF��%�R*ڿ�<¿�"���͊�$@^�~+�X��B̷�"<��?�-�$��5��S��(&�)���4���^���������xν���AH�����o�nu��K��g�Z�˽�_��-#y�M�.���"R�� XE�q|����)!_��ý�?��ot����z����)��/]�8���B���y¿��ڿp��u����   �   2#��0߿�0Կ�,ÿ����'���Ow�T�E�8P�ӗ�����c�A��ȺϽ�&���`T�ۧ<�I�K�,>z��G�� ̽�������!~/��aD�XJT���]�a~_��qY�x�K��8�;u�F��&ѽග���]�u:�b�׼��ż���-0V��n�����!cZ�ӡ��;�w���mE�}�w�w����:����ÿ��Կ2�߿�   �   ~ſ����_�����r���c�T���)���ML¾d���	%C��t�a˶��"���[�t_�t�� ����?㽎��@R5�$ Z��?}�l�����`���:��,e���+���d��l�n��H�>�!� C��ȸ�}��ć;�vD�X0���P����$&��vP=���ӎ������z*�4V��{��		��
����¸��¿�   �   �w��[r��|2��-z����z�0�V�/'1�����ؾg꠾�Jg���!��߽꿞�p�y�q�l�Ű�����K�U�1�J�E?}� ���ܱ�.Ⱦ�wپ8��J�PS⾟�վ��¾�+��?����ml��g9�J���
˽%���W��;��dR�X��zwֽI��4Cg�"ࡾڤھ�m���2�ϽX� "}� ���������   �   0��ݩ����y�K�d��KJ��,��E�T'��{�������8����>����ɉ�ƀs����1������� T��Y���䫾��ϾK�򾶳����TI���Z�t���*��j��Ⱦ����R��F�8���nн��aBj��C]�Ү���ĵ��b��_<��Q��6���e����S/���L��g��}{�>(���   �   � R���M�0C��V2��o�� ���ܾ'ܮ�Kȅ���E�O��7�Ƚg�����r�~�w��9���wԽ���`�N�^������n��)	�OM �J�4���D��N� R��M�sC��Y2��r��"�L�ܾ߮��ʅ�e�E����|�ȽJ���V�r�h�w��7��}tԽ����N����ؕ����⾪&	��J �5�4���D���N��   �   ��#W����(�@f�3�Ⱦ�������)F�G���jнI��i?j��B]������Ƶ�fd�Xb<��S�����i�6��7V/���L�Dg�x�{�+*��2��ī��<�y���d��NJ�o�,��G��*�n~������ʫ8�j��v����ʉ�k�s�@��d.�������T�<W��`᫾��Ͼ��������YF��   �   �E羅N��վ��¾(������hl�sc9�
��˽�����W�V�;��dR�QY���yֽT��?Fg�H⡾��ھ�o�I�2���X�Z%}�Ꚏ���������y��Ut��]4���{����z�ЛV�\)1�\�i�ؾd젾lMg���!���߽"�����y���l��������=F�fR���J��9}�ȫ��Oر��Ⱦ
sپA3��   �   �6��ua��9(���a����n��H�'�!��<���¸�:y��>�;�A��.���P�s����(���R=��������J��{|*��V�}���
�������ĸ��¿{ſ���������������T�b�)�b��DN¾ʹ���&C�(v��̶�C#���[� q_��
��`���}:�>��N5�'�Y��9}�&��h��B\���   �   �x_� lY�>�K��7��p�PB�v ѽԱ���]��4��׼��ż���1V�p�����(eZ�N��� =�ٜ��oE���w�����1<��H�ÿ��Կ�߿%㿊2߿�2Կ
.ÿj����(���Qw��E�lQ����U	��M�c�b���Ͻd'��r`T���<���K��8z��C���˽u����}��y/��\D�ET�'�]��   �   �k��q��G� a�V�˽�Z��Yy��.��|༸I��lLE��j|���<"_�^�ý�@��qt�󲾥|��� *�w1]�%���W��;{¿�ڿ����������G����+ڿ�=¿�#��sΊ�kA^�+��Y��Mͷ��<��.�-�8 罨M�S�"'&�����4���^���F����sν}{�M��D�����   �   P�ǽ�/���'���˘���{�P�@�(���l�����`C0�������0mܼ��h���ѽ{P,�6���K2¾Nz�s8��o�����uŴ��=ҿ�J�l �,��A	���JS ��9��jҿ�9��	���-�q�A�:�v
�`:Ⱦ(���rR=�n������0V������ ������8lA� 2m�e���颽M!��X8½��Ƚ�   �   �(��2���s���M�\�!����p���H`»��: ��; �\;�л�fռg�o��y۽c�4�t*����˾�X��A�ϟ{�yG��\q��BBܿS������j��b�������������ܿ�7���H��o�}� WD��V�}�Ҿ���X<G��?����\
Y���������Ӽ�?�){�1�.��O�vo��q���Y��&%���   �   �py�4�i��P��m-��O���$�1� ú���;,<��;P-�� eӼ�r���޽��7��q���SϾ�����D����{ǟ�Uj�� �߿Kt��d�����>P�������7����P��N���䠿< ��ͮG�����j־����کJ�`n�Tj��Z4Z����4ּ�s¼`kԼ�X���x��}7���R�B0i��Kx��~��   �   �(���1���s���M�L�!�P��>����^»��:p��;�];8�л�dռЂo�nx۽��4��)����˾+X�G�A�Ǟ{��F���p��cAܿY�����֔����������������ܿ�6���G��[�}�(VD�,V���Ҿ���f;G�@?�����Y����Ȭ�`�Ӽ`>�z���.���O�o�qq��pY��%���   �   3�ǽ�/��v'��|˘���{�'�@����0l��d���90����h��$iܼ��h�R�ѽ�N,�����0¾#y�~q8��o�����Ĵ�<ҿI� k ��n@	���@R ��7�)iҿE8��ǯ�� �q���:�@	��8Ⱦ䱋��P=������}���-V�|���� ����ɬ�kA� 1m��d���颽!��$8½��Ƚ�   �   �k��q��G�
a�@�˽�Z��y���.��{�H��tGE�,c|�T}� _�7�ý^>�<nt���hy����)��.]�q���R���x¿m�ڿ�����������D�����(ڿc;¿�!���̊��>^��|+�4V���ʷ�;����-����
혽h�S�$&� ���4���^�A������sν{��rD�����   �   �x_�lY�4�K���7��p�DB�V ѽ����^�]��3�2�׼8�żK���+V�>l��/��.aZ�����C9�E��?lE���w�P���c9��'�ÿ1�Կr�߿b!��.߿;/Կ�*ÿ�����&���Mw���E��N����k���c�f��̷Ͻ>$���[T��<���K�*6z��B��3�˽�����}��y/��\D��DT��]��   �   �6��ma��4(���a����n��H��!�J<���¸��x����;��>�.+���P�F����"��AN=�x�Ԍ������x*�	V�lz�����`������¿�ſ!����췿�������
����T���)�����I¾����k"C��r�ȶ������[�m_�H	�����\9�����M5���Y�~9}���S��3\���   �   �E�N��վ~�¾(������hl�Yc9����˽����W�~�;��^R�
U���sֽ��@g�ޡ�#�ھ(l���2�.�X�}�h�������𢿊u��[p���0��cx��r�z�\�V��$1�����ؾ蠾Gg���!�ܮ߽Q�����y�U�l���������D��Q�w�J��9}�����-ر��Ⱦ�rپ53��   �   ��"W����(�>f�-�Ⱦ������� F�
���iн
���;j�>=]���������2`��\<��O�����:b���
Q/���L��g�+z{�W&��*.��񧃿�y��d��HJ�B�,�oC��#�y��������8�����>Ɖ��ys����n,��4�}��T� W��-᫾��Ͼ��������SF��   �   � R���M�1C��V2��o�� ���ܾܮ�;ȅ�ɵE�����Ƚ������r���w�@4���oԽ@}�&�N����Ȓ�����^$	��G �2�4�S�D��N��Q�1�M���B�pS2�m�4��|ܾ�خ��Ņ�
�E�@��\�Ƚ_�����r��w��5���rԽj�M�N��������^�⾗&	��J �.�4���D���N��   �   0��ݩ����y�N�d��KJ��,��E�L'��{������ͨ8����򶽨ǉ�zs����;*����Ϊ�fT��T��ޫ���Ͼ�򾀮�ں�_C���&T����r%��a�&�Ⱦ+������F�؅�8eн����7j��;]�����µ��a��^<�RQ����ke����S/���L��g��}{�=(���   �   �w��\r��~2��/z����z�0�V�,'1�����ؾU꠾YJg�:�!�ر߽�����y�8�l���������@��N�~�J��4}������Ա��Ⱦpnپk.��@羨I�t�վ>�¾I$����/cl��^9�f��F ˽����W���;��]R��U���uֽ����Bg��ߡ���ھ�m���2�ŽX�"}����������   �   �ſ����a�����s���d�T���)���@L¾N����$C�st��ɶ�� ��O�[��j_��������4㽨���I5��Y��3}�������~X��3���]���$��k^��ŏn���H���!�K5�����zt���z;��:�
)���P� ����$���O=��󉾬�������z*�*V��{��	������¸��¿�   �   4#��0߿�0Կ�,ÿ����'���Ow�S�E�5P�ʗ����U�c������Ͻ!%���[T���<�j�K�1z�&?����˽չ��z�_u/��WD��?T���]�s_��fY���K��7��l�p>��ѽL�����]�-���׼(�ż̐� ,V�m�����bZ������:�l���mE�v�w�u����:����ÿ��Կ7�߿�   �   ����eF��'�U*ڿ�<¿�"���͊�$@^�~+�X��8̷�<����-�Q���혽ΞS�L#&�
��4�ھ^� �������nν1u�� ��@�����g��m�-D�*Z��˽<U���y��.�|o��>��:E�lZ|�J{�/_��ý?�xot����z����)��/]�6���@���y¿��ڿr��w����   �   �@	�����R ��8�jҿ9��~���N�q���:��	��9Ⱦ�����Q=�0��x~��5.V�(���� �Z�����gA��+m��a���墽����3½��ȽN�ǽ�*���"��ǘ���{�/�@���Lb�����	0��������gܼ��h���ѽPO,�k���81¾�y�r8���o�����Ĵ��<ҿ�I�~k ����   �   ��F��О����o�ܿ97��WH���}��VD��V�7�Ҿp��<G��?�e��T	Y����ث�|�Ӽ�;�x�B�.���O���n�ro��DW���"��o&���/��0	s���M�j�!�v��^�@K»@M�:د�;�];�л�cռ��o��x۽��4��)��8�˾XX���A�"�{�G���p���AܿÒ��L�����   �   @俜s��vտ�ZĿ���������x�<G�v�W{��v�m�c�%�����۞�ad���0�Q��|��mX��Z#��1��|?���J�֕Q�g�R��OM�'@�4,����z�޼0ē�� ��>5:\�<��k<��<��j<��;|[5�T��@�����oZV��8��^!߾��L�D�U*w��g���5���#Ŀ�eտs��   �   !�࿘�ܿ�ҿ�6��-Ы�������t���C�~j�R�⾞����i���"�q�ེe���b���0�H���5�����.���@���Q�y!`���i��lm�.~i�\d]��H�Cp,�9@	���¼l-^�0�o��;h8<<еm<Q<��;\:����ۜ�B����R�ܮ��s�۾l����A�c8s�N��z������ҿG�ܿ�   �   ]/ֿ��ҿ15ȿ������Z~����h��=:����(;׾�g����]��}��~ս9s����[���1��w#��2(�&�9�.wR�\In�ڄ�����B����������n����n��芀�NX�)�$���g��Ⱦû��-; ��;��< �:��I�������c ��I��O��hѾ���5�8�w�g�*������$���Vȿޫҿ�   �   S�ſ�h¿�Ÿ�cΩ�"Җ��_���7V�3++�0$���žL}���^K�=��9Ľ�,����S���5��4���F�z?g�KL����4���XCʽl0۽����2뽒�b�ܽ`�ɽF���%b��*{c��"���ʼpcK��3x� N�� CS��+j�!r�ዽ��ܖ9��ӈ��������)*�ݻU�\������D�����~�¿�   �   �䰿�ɭ�"��ݔ��,|��lf�\�>�t�����4���=~���3�����U宽�W~���L�}h?�P9O��Qu�D蕽ԛ���ڽ����D�����<2(�A�-�+A-�j'�&;���
��/�X+�������U��	��̧�<�H��2�>ꐼ�m������սC2&���t��/��4�����>�>�Yg�T���! �����p���   �   ��Q��B����܂�8�g��YF���#�Z��'#ɾ���WY�����GֽL×���f�ΎI�͂Q��(x���&�Ž9���7����0��fJ���`�	Jq�:�z�}P|��%u�V�e���O��m4��^��}�C������x^/�DI�\���d���B���g��˻�<��&MT�P ����ɾ�:���$��G��oi�����9I�������   �   &��v\{�Q[n��WZ� &A���$�����wؾg�����w��3�K����+����~R���M�8o��昽H�Ƚk���h%��`K��Ur��Ջ�l5���Ѩ�jl��?6���譾�֣�u放�l����[�212�La
�(eͽ�ϑ�[�I���� ��1n�c�S�H���/����-3���z���v�۾��	�M'��CC�Z=\���o�f%|��   �   ��N�� K�fL@���/��\�,t� ھ�/��߄�E�t��(�ǽBލ��Y��<E���[��������6�̮*�}�Z�����Ԓ��i�����ӾM�����8�󾬦��m�M�;UĴ�Q���z�Q%E�N�F�ؽaژ�baX�5�'�>� ���E��&���:ͽV��szM���в�
�߾�Y���`-2�R�A��K��   �   �!��T�%�����`F�H;����@n���K� ��ֽ�ז��\��8�s�@��t��Ω����Xq$��k[�󃍾�x��$�Ծp���F��`��@O�՛!�.W����1��uJ��K;�����p��y�K���� ֽrږ�c�\�o�8��@���t�e̩����n$�>h[������u����ԾB�����Э��L��   �   ���"�i�_�;����N��,�z�Y!E�4���ؽ�֘��\X�y�'�R� ���E�(��4=ͽe��h}M������Ҳ�\�߾�[�0�02�.�A��K�� O��K�4O@�W�/��^�v�8ھ|2������E����3�ǽ9����Y�0=E��[��������4�ի*���Z�6~��ԏ��䭼���Ӿ���0���   �   2��	孾3ӣ�D㔾�i���[�-2�^
��_ͽ�ˑ���I�������m���S�
���-����/3���z�6��K�۾e�	�t'�aFC�'@\���o��(|�����_{�E^n�~ZZ�c(A���$�y��Tzؾy�����w��3�����-��H���~R��M��o�f䘽��Ƚ
���e%��\K�(Qr��ҋ�72��*Ψ��h���   �   �J|��u���e���O�}i4��Z�Yw��=��ʕ��X/�@�x���4a��C���g��ͻ�˴�wOT��!��ʂɾ<���$��G�hri�����J��=�������R������+ނ���g��[F���#����4%ɾ����YY�T���Iֽ�ė���f���I�
�Q�g%x�(�}�ŽW��� ��-�0�bJ�Ɗ`��Dq���z��   �   �<-�,'�7��
��(�%������vU�o��§�`�H���1��萼rn������ս�3&�ît��1��N��*����>�\g�|���i!��n������0氿˭�x�����@}��Xnf��>���`��K6���?~��3������殽�X~�يL�gg?��6O��Mu��啽1���]ڽ����������5.(���-��   �   ~��b�ܽ��ɽ�{��`]���rc�}"���ʼ�PK�P�w� ��,S�4*j��r�⋽���3�9��Ԉ�U���҄�'+*�M�U��\��� ��Y�������¿��ſ�i¿�Ƹ�eϩ�Ӗ�F`���8V�3,+��$�Ցž~��%`K���:Ľ:-���S� �5�74���F��;g��I����H����>ʽ<+۽ݛ��,��   �   �����j��B���<GX��)�����^����û�$.;��;ȭ<@1�:��I����y���d ��I�EP��tѾo���8���g��*��k����$��{Wȿ��ҿ;0ֿ��ҿ�5ȿ���,����~����h��>:����;׾%h����]�.~�Bս�s��!�[�@�1��v#�:1(�ġ9��sR�9En��ׄ������>��(��������   �   �`]�k�H��l,��<	���¼#^� �o�`��;><<��m<�Q<��;�:�|�Pܜ����f�R�T����۾ڮ�Z�A�9s����mz�����Nҿ��ܿ����ܿ_ҿ57��yЫ�癓�R�t���C��j����ְ��Z�i��"�����e���b���0�ҩ��4�����.���@��Q��`�j�i�bim�~zi��   �   @�4,������޼Zē�H!��75:��<l�k<��<(�j<�}�;�\5����`@�����ZV�9���!߾��o�D�z*w��g���5���#Ŀ�eտs�@俗s��vտ|ZĿ���������x��;G�Y�&{�ɋ��>�m�8�%�[�佼۞��`d�Z�0�/��`��PX��Z#���1��|?�x�J���Q�R�R��OM��   �   R`]�=�H��l,��<	���¼�"^���o����;�><<�m<hQ<P�;p:�-�`ۜ���k�R�����(�۾8����A�8s����y��2��wҿ��ܿ����ܿ�ҿk6���ϫ�I���I�t�&�C�j�������G�i�J�"�����d��zb�3�0�����3���!�.�͔@�x�Q�`���i�im�1zi��   �   Y����j�� ���GX��)���R^����û`+.; �;�<�U�:��I�(�����[c �I��N���Ѿ;����8���g��)�����i#���Uȿ�ҿ�.ֿِҿY4ȿG��Ҡ���}����h��<:����:׾�f����]��|��|ս�q��=�[���1��t#�O/(��9�YrR��Cn��ք����F>��̈�������   �   2��+�ܽ~�ɽ�{��@]���rc�1"�$�ʼ�NK���w����� S�� j�To�~ߋ��~��9��҈�����(�� )*���U�Z[������J�����V�¿#�ſog¿�ĸ�Nͩ�$і��^��&6V��)+�9#�8�ž.|��K]K����6Ľ�*���S���5�84�P�F�E9g��H���j���>ʽ�*۽b��n,��   �   �<-�'��6�У
��(�[%��v���
U���(���P�H�d�1��␼Fj����*�ս�0&�f�t��.��S�辘����>��g�C������������P㰿Dȭ�������� {��rjf���>�	�C��/3���:~���3������⮽�R~��L�Rc?�l3O��Ju�䕽営�6ڽ�������{���-(�ɉ-��   �   �J|��u���e�|�O�ii4��Z�$wｍ=��v���*W/�2=�@��Z��q>���g��Ȼ�b���JT����{~ɾ@9�4�$��G��mi�^����G��%������vO��ª��pۂ���g�eWF��#�؇�� ɾ;
���TY����(Dֽa���&�f�5�I��|Q�t!x�g�Ž���~����0��aJ�e�`�SDq�H�z��   �   l2���䭾)ӣ�;㔾�i����[�-2��]
��_ͽ`ˑ�%�I���\���i��S����8���-+3�7�z������۾��	�>'�yAC��:\���o�G"|����KY{�IXn��TZ�w#A���$�����tؾ
���/�w��3�����'�����xR���M�o�j☽�Ƚ@��%e%��[K��Pr��ҋ�2��Ψ��h���   �   ����i�X�;����N���z�=!E�
��ؽ@֘��ZX�^�'��� ���E�I#���6ͽΞ�2wM���sͲ���߾�W��	��*2�}�A��K���N���J��I@��/�"Z�r���پ-���܄��
E�¦�؉ǽ�ڍ���Y��6E�ɭ[�������3��*��Z��}������������Ӿ׹����   �   �!��T�$�����\F�zH;����3n����K���>ֽ�֖�)�\���8�6�@�3�t�{ȩ�3�k$�\d[�2���r����Ծ����}�B���I�\�!��Q����}��B��D;�����k��ڴK�����ֽ�Ӗ��\���8���@�Њt�Vʩ�O��n$��g[�T����u��Z�Ծ�����ĭ��L��   �   ��N�� K�dL@���/��\�)t���پ�/���ބ��E�2��S�ǽݍ�[�Y�p7E�ج[�I���
��
2�_�*�O�Z��{������O�����Ӿ��徔����󾂝�:e�N};:����J����z��E�����ؽrҘ�LUX��'�1� ��E�h$���8ͽ����yM����ϲ���߾�Y���S-2�I�A��K��   �   %��v\{�R[n��WZ�&A���$�����wؾX�����w�a3������*��|��syR�>�M��
o�n�����Ƚ��5b%�AXK�Lr��ϋ��.���ʨ��d���.��D᭾�ϣ��ߔ��f����[��(2�eZ
�ZͽǑ�،I����$���#h���S�p�������-3���z����A�۾��	�<'��CC�Q=\���o�d%|��   �   ��Q��C����܂�8�g��YF���#�X��#ɾ��nWY�|���Fֽ�ۂf�d�I�@{Q��x�웽��Žh�������0�j]J���`��>q���z��D|��u�K�e�_�O��d4��V�jp��7�����GP/�3�X꯼W���=���g�Fʻ�����LT� ��d�ɾ�:���$�޽G��oi�����8I�������   �   �䰿�ɭ�%��ޔ��-|���lf�]�>�s�z���4��q=~�x�3����_䮽�T~���L��b?�l1O�+Gu��ᕽ�����ڽ����j������)(���-�\8-��'��2���
��!�O��\�����T����������H���1����j����}�ս�1&�#�t��/�������4�>�Qg�Q��� �����q���   �   T�ſ�h¿�Ÿ�eΩ�#Җ��_���7V�3++�.$���žB}���^K���_8Ľ�+����S�e�5�4��F��5g�OF���잽�����9ʽ�%۽ݕ潐&�-��*�ܽ��ɽhv��TX���ic���!���ʼ;K�`�w� J~� �R��j�So��ߋ����9��ӈ�����߃��)*�ջU�\������D�������¿�   �   _/ֿ��ҿ25ȿ������Y~����h��=:����%;׾�g����]��}�~ս�r����[���1�-t#��-(��9�roR�@n��Ԅ�I���;��P����񟽊����f��v��� @X��)����T��p~û _.;@�;��<�}�:8�I�������c ��I�lO��TѾ���0�8�t�g�*������$���Vȿ�ҿ�   �   #�࿘�ܿ�ҿ�6��-Ы�������t���C�~j�P�⾜����i���"�:��le���b�\�0�p��>3�����.��@�D�Q�b`���i��em��vi��\]���H��h,�q9	�V�¼�^� �o���;hE<<(�m<,Q<��;�:���iۜ�����R�Ю��j�۾j����A�a8s�M��z������ҿG�ܿ�   �   O�����ӭ�������䂿�Y`���9�����P��+��2)����?�
��^vֽPȩ��0��P���Tw��Bu�\�v�5bx�CEw�S�r�1�i��"]�KL��a7�O��/��
üz�(ѻ0�;e+<���<Z�<���<p̴<�8v< `�:�1��U�P�0��*����h����l�T��8�TG_�蔂� e���������   �   �B��Lb��m��~"��ƽ���\�{�6�ES�Zf��0������L<�l1��ҽ�ꦽ.���,����v���v�E�z���~� I��Ь~�I�x��zn�:�_��<L�.4�����M�<ڤ��1� �ѺH�;��k<"ҡ<��<�ԩ<�Ph<��:�䠼Q�M��(���x��Xe��v���ܾ���#5��[�,}���	����Vg���   �   �;��v��.����#����t���Q���-����
ؾ����G�r�F�2�����ǽ~���2���*;z��]v�1�|�P̃� ���t�������@��~㑽������uwv��Y� '7��1��ȼ�`�`6`���;ܵN<n^�<n��<�=< ��8n��Y�E�˺������Z��难$%Ҿ#'	�m�,��AQ�k�t��.��W���u����   �   ����|������=g~�]pa���@�����v���Wƾ�	��}�^��g#��� ���Ze��)�~�]r��w��1������3-���K��
���JP���f���h���������d����J��0�w��C�^����������� :�}�;,.<x �; ���{��3�9�H���ٍJ�T6���¾����7�@�V�a�
�~��势�2���   �   s���?���+w�{�b�X�H���+�A�����J쯾u脾��D�n�1Խ&U��u����l���k�~�~ǎ����j���%Ͻ�}�f9��=��T9�N�\��>m���I�B�Ƚ�j���̃��|@�����<֊��ӻ ݹ 59l���ꟼPP,��{��3,���=6�銀��Э�lV⾤%�mJ,��I�U�c���w��v���   �   ��d�ԧ`��U��C�r�,�p�u�|¾�����c��'��A������r䉽׃g���[��j�����V���.�����V��T���,%� �2�`<���@�]`?���7�H�*��o�:���gֽ�¦���s�O$���ɼ�f�8���:������� �Zo���lؽ%����`��M���yľF���
��..�<�D�9V�u?a��   �   ��>��Q;�u1�]"�u�����J�ɾ����=�x���:�y��ƽ.���d�>=J�t�O�Tp��������>��5����'�j�B��/\��r��0������.��/򁾟ss�%\��~?�N* �AQ ��Ľ�����B��` ��%��,���� ƼR��O�u��>���^	��?�Q^�����9Ͼ/$��(���c$��2�<��   �   �"�9�;��+��mf澔Iľʀ���e��[sE�
!���ս�@�c�Vg9��:2�.K�T���FϨ���ܽ���_�0�D�V�A}�����+�����Qٴ��[��3ű��j��F4��4z��y�a��x7�hT�%�ֽ�(����V�{��4�������e^�0 ��齓� �)6U�n͈�rة�4̾�1�XJ�z�����   �   ��W��q޾��ʾ����=���W�x���D�W���EܽL{��kT`��)�ky���!���O��莽FŽ�%��_.��N]��%��od��������Ѿ�R㾿����K�뾬u޾��ʾ��������x�	�D� ��8Jܽ�~��2Y`��)�O{���!��O�R玽�CŽB$�n].�sK]��#���a������{�ѾO�����   �   �X������og��X1���w����a��t7�\Q�J�ֽ�$���{V�V��ʜ�����Jg^��!���齔� ��8U�Lψ��ک�̾65�JL����U���$�r�V�����i�{Lľ2����g��evE�_#�$�ս������c��i9��;2��K�~����ͨ���ܽ�����0�ϟV��<}�a���(������մ��   �   k��wlns�\�[�:z?��& �!N �lĽ�
��>�B��[ �,������B�ż���]�u��@��`	�I�?��_���量�<ϾR'�� ���e$�Q�2�b<�6�>��S;�?w1�_"��v�������ɾ� ��h�x��:�S��ԁƽ(����d��>J�םO�.Sp����p���0����њ'���B��+\�Hr�.��䰅��   �   \?���7�6�*�(l�����aֽ����o{s�hH$�$�ɼ��e�����:�䀬��� ��p���nؽ����`�xO���{ľ�H��U�b0.�R�D�V��Aa�d�d�+�`�*U��C�8�,��q��w�~¾����	 c�ڃ'�yD�������剽��g�ʮ[�Aj������������|��<������)%�k�2�\<���@��   �   $���f��zC彊�Ƚ�e��Xȃ�u@�$y���ˊ��qӻ ܹ .9d���ꟼvQ,��|��@.���?6����vҭ�hX��&��K,�҇I�H�c���w�x������1@���-w�W�b���H�`�+�f��[�⾴��鄾[�D���Խ�V���u����l���k�X~��Ǝ�z��� ����!Ͻ�y佾4�����c6�*��   �   ����}��wF��	�w��xC�����D�� �:0��;`6<�;0��R|��a�9�n��7�J�O7��8¾������@���a���~��抿�3��w���b��\����h~��qa�$�@����x���Xƾl
��̓^��h#�B� ���"f��*�~�u]r���w��0�������+���I��[���M��<c���d�������   �   �qv�J�Y�l!7��,��Ǽ@`���_����;4�N<$b�<��<��=< ��8,��g�E�����ƅ���Z�vꚾ*&Ҿ�'	�=�,��BQ���t�S/������ ���,<���v��ɂ��{$��r�t���Q���-��zؾ6���+�r��2����Y�ǽ��������;z��]v���|��˃�������G���>��ᑽu�������   �   -+4���H�դ�̋1� qѺ�;P�k<lԡ<��<�թ<$Rh<@�:�堼�M�t)��/y�JYe�bw����ܾ����#5���[�|}��+
��u���g���B���b������"�� ���{�\�Ĭ6�~S��f� 1�����M<��1�h�ҽ립I.���,����v���v���z���~�pH���~�;�x�xxn���_��9L��   �   =��)��üz�hѻ �;�d+<x��<"�<���<8̴<8v<@[�:<2����P�v��Z����h�����!T��8�qG_�����e��������P�����˭�������䂿~Y`���9�����P��+��)��_�?���<vֽ;ȩ��0��P���Tw��Bu�@�v�bx�#Ew�.�r��i��"]��JL�wa7��   �   �*4�����G�Ԥ�4�1��mѺP�;�k<�ԡ<�<�֩<Th<� �:�㠼��M�d(��rx�CXe��v��ƂܾL���"5���[��|���	�����g��CB���a����&"��u�����\���6��R��e�=0�����0L<��0�C�ҽꦽr-��,���v�I�v�a�z���~��G���~�X�x��wn��_�]9L��   �   �pv���Y�� 7�:,���Ǽ `���_����;��N<c�<d��<��=< ��8<����E�����X����Z�难\$Ҿ�&	�Ȇ,��@Q�}�t�/.������Ӈ���:��bu������R#��`�t���Q�'�-����	ؾĈ����r�=�2�<��.�ǽ@�������8z� [v��|�rʃ�ݴ�����Q
��>��j���唍�m���   �   ����~}��*F����w�;xC�v���쭼h����:���;<:<��;0���v��Y~9��먽��v�J�n5���¾������@���a���~��䊿2��������������e~��na���@�����t��VVƾj����^��f#�� �����c����~�0Yr���w�/������*��H������K��Hb���c�������   �   ���pf��*C�L�Ƚie�� ȃ��t@�$x���ʊ��kӻ�w۹ �9�Q��$䟼�L,�|y��y)��1<6�ǉ��ϭ��T�~$�I,�s�I�~~c���w��u��Y���>��m)w���b���H�m�+����f�⾙꯾$焾��D����Խ�R���r���l���k��~�NĎ�]���'���& Ͻ#x�c3�����5����   �   �[?���7��*�l�����aֽ@����zs��G$�`�ɼ�e�h��̃:�hy��8� ��l���iؽ%��)�`�AL���wľ�C��3	��,.�5�D�V�=a���d�s�`��U�sC���,�jn�9r�?z¾%����c��'�<>�������ች�~g���[��j�X���r����
��e��F�����)%���2��[<�h�@��   �   G��Z@ns�;�[�z?��& �N �(ĽN
��c�B��Z �����򛼜�żX����u�|;��r\	�\�?��\��c륾Q7Ͼ!��U���a$���2��<�a�>�O;��r1��Z"�s�T�����ɾ������x�ּ:�9��k{ƽ	��j�d��7J���O�zMp���𖹽غ���ؙ'�$�B��*\��r��-�������   �   aX������\g��I1���w���a��t7�<Q���ֽ�$���zV�������\Ｇ���_^������݄ ��2U�Zˈ��թ�,̾I.�bH�W�����e ������)���b�wFľ,~���c���oE�J�5�սP����c��a9��42��K������ʨ���ܽv����0��V�	<}����(������մ��   �   ���B��q޾w�ʾ����2���?�x�h�D�4���Eܽ�z���R`�W)��u���!��O��㎽�?Ž�!�?Z.��G]�s!��_��b�����Ѿ5K㾷�����@{�n޾��ʾr���u�����x���D�6���@ܽ2w���M`���(��s��!�m�O��䎽nAŽ*#�j\.��J]�`#���a��D���?�Ѿ�N㾤���   �   �"�2�6��'��gf澊Iľ�����e��;sE�� � �ս9���3�c�Pd9�j62�K�����ɨ�#�ܽ���3�0���V�8}��	���%���|��|Ҵ��T��]���d��H.���t��9�a��p7��M�Ʀֽy ��|tV���|����2���`^���� 齟� �I5U�
͈�ة��̾�1�?J�i�����   �   ��>�|Q;�u1�]"��t�����A�ɾ����!�x���:�H��~~ƽU����d��9J�A�O��Lp����������D�'��B��&\�.
r�E+��	��������쁾�hs�W�[��u?��" ��J ��Ľ�����B�rU � ���훼�żY���u�=���]	�D�?��]��2��9Ͼ�#�����c$� �2��<��   �   ��d�ӧ`��U��C�o�,�p��t�||¾꧖��c��'�RA��햳�l㉽؀g���[��j�ď��,������o��O��]��&%�V�2��W<�E�@�~W?�<�7��*�,h�B���[ֽ���7rs��@$�P�ɼ,�e�l��|:��w���� ��m�� kؽr���`��M���yľ�E���
�v..�0�D�3V�q?a��   �   t���?���+w�}�b�X�H���+�?�����B쯾j脾��D�B��ԽdT���s��R�l���k� ~��Î�󫢽���JϽt��.��n��3������`���<�~�Ƚ&`��xÃ��l@��j��ڿ��0Iӻ �ٹ 9hF��*㟼M,�Lz���*��d=6������Э�?V⾑%�]J,�	�I�N�c���w��v���   �   ����}������?g~�\pa���@�����v���Wƾ�	��f�^��g#�_�m����d����~��Yr���w��.������(��F�����H���^���_������#����x���A��P�w��pC�М�P᭼����:x��;�C< #�;���Fv���~9�H쨽���s�J�)6���¾�����-�@�O�a��~��势�2���   �   �;��v��/����#����t���Q���-����
ؾ����9�r�0�2����6�ǽ����v���9z�[v�x�|��Ƀ����ֱ�����.<��-ޑ�Y������Ckv��Y�g7��&���Ǽ��_�p�_���;8�N< g�<t��<�=< �8���؍E�$������Z��难%Ҿ'	�e�,��AQ�h�t��.��W���w����   �   �B��Lb��n��~"��ƽ���\�{�6�ES�Yf㾾0������L<�Z1�ާҽ�ꦽ�-��>,���v��v���z���~�VG����~���x��un���_��6L�(4���,B�Ϥ���1��(Ѻ8,�;<�k<rס<��<Bة<�Vh<@�:㠼��M�(���x�|Xe��v���ܾ��#5��[�,}���	����Wg���   �   *<y���t��h��5U���<�-�!��t��پ�R��\��)jO��#��X�oE��սn�ͽ�OͽPiϽF�н�AϽ�yɽ�;�����矽𝌽�(p�A�E����"��B������� k�:��)< K�<���<W�<���<�%�<v��<@><P��z���$���ؽ�`%�~Gl��Π��/ҾST��� �@R<��T��qh�<�t��   �   v(u���p���d�-�Q�R�9��5�r1��hվQi��\��&�K��	!����b!��qѽʆʽ�ʽ�5ͽV]Ͻ|�ν,�ɽF���s
��x��������|�@#T��*��� ��X��xC8��gҺ�V�;y<B
�<���<j�<̦�<0�<�v6<�̬����w�{���ս�#�1�h��[����ξ�:��!��G9�3�Q���d��p��   �   �Pi�|:e��Y��gG�̣0��V�C����ʾ ���g�x��UA�v�������ؽ�ƽ{.���½�ǽt˽��ͽ�̽)�ƽm���;��ޑ���������Y�qr0�#�4 ��A�����s�;�pq<��<~z�<X̾<�f�<��<@����缦�r�fEͽJ:�a�^�tK��}pžR�����%x0�C~G���Y��Xe��   �   F�V�(�R��"H�;c7��b"���\��@0��Zɒ�d�i�0�z`�L��tOŽP~��4��H㶽YR���pƽSͽ��н̀ѽf�ν��Ƚk���U���󥽄d���/W��:(��S��_��(0ֻЖI;ئ/<��<�H�<4�n<���;������e�"������!SO�Gn��$ֶ����1���"���7�X�H�9<S��   �   �Y?��;�2��#�nU������̾b+������I�h�����U�ǽ�����3��P���XS������k½��Ͻ��ڽ�<꽉>�����b�޽h�н��a�����Fa_��i$���ּ��_���N��q�;�2
<X�<P�;@��4޼��W�0ѱ��o��Z<���}������ξ3���}�(*$���2��E<��   �   ��$�l�!��>��?�r���&Ծ	ï�Ns���1^��+���eGν�����������
���`������Y׽	���h ��_	�6��z��Z�����M�����������ؽjf���.����V�z���Z���+��\������}�cN����I�K��͢�ni�)�'�rm`����E�����ؾ�c��������r"��   �   M�	����h"���=龧ξw������K�i�h�6���±ս:��������o�Hl�z~��������еƽ���cO��J�͓%��)4���?���G��^J�,sG�A�>�
f0����|\�$߽�V��4���3�6�������0�L�BI��#��8%�� E��ϕ��y׽&���%C���x�$���iķ�X�Ծ��������   �   �޾��پ�;����{M��Ќ���g��9����U�ٽN£��&{��eM�<�O7D���b��I��-M���ҽ�����N�6�1���J��<b��v��C�����Խ���L��R�q���Z�dp>����s� �+�ǽ����S��Y�:�ټȞ���fϼ�_
�J�E�����ߛ½��@X(�TS�zӀ�����GT���bþ��ҾF`ܾ�   �   T����F���<��ʳ������X��_1�
��սhܞ�BQi��0�l�����'#��wO�̰��⚳�g����R�2�a�U���y�x���eY���|��4�/����I���?��C���'����X�c1���U�ս�ߞ��Vi�]0����Y��)#��xO����������罒��U�2���U�%�y�m���W��Pz��k��   �   l����J����q�^}Z��l>������ ���ǽ����~S��T�`�ټ옻��bϼ�^
��E�8���,�½���Y(�gVS�
Հ������V���eþ��ҾocܾQ�޾��پ�;�����O��.Ҍ��h�� 9����ٽMţ�u+{��iM�<��9D�[�b�"J���L����ҽ����IM��1��J�v9b��v�TA��u����   �   FoG�b�>�Ob0��XY��߽3R��F�����6�H����X�L�|8I�� ��$��� E��Е�y{׽z���'C�-�x�ߟ���Ʒ���Ծ��� ��p���	�9���%���@�>
ξ��������N�i�Ց6���޴ս��������e�o��l��{~���Đ��2�ƽz��>N�I���%�G'4�h�?�"�G�$[J��   �   B���������@�ؽla���*��0�V���P���+� I\��{�p�}��^N�j��*�K�Ϣ�Nk��'�~o`��������̻ؾFf��%�����t"�F�$��!�z@�A����(Ծ�į��t���3^���+�B��Iν������j������
��6a�������X׽��콢g �^	�7�����������   �   ��н�������}���Y_��b$���ּЯ_��N���;=
<�<�	;���޼�W�Zұ��p�/\<���}�蠤��ξP���~��+$�K�2�,G<�8[?���;��2�I#��V����I�̾�,�������I����E���-�ǽK����4��r���6T��^��l½6�Ͻ��ڽx��9꽢;�@�����޽�   �   L씽�`���)W��4(��H��U���ֻ�I;ز/<Ȧ�<nL�<��n<h��;ȱ໦ ��e�A������lTO�*o��U׶������"���7���H��=S���V�z�R�$H�\d7��c"�|����\1��:ʒ��d���0�ba�����PŽ{��7�� 䶽�R��qƽ<ͽt�н�ѽ�ν��Ƚ����UR�����   �   yY�<n0��^����	A��+񺀊�;�yq<��<�}�<�ξ<8h�<X�<8�������r�SFͽ ;�d�^�&L��dqž6S��p���x0�&G���Y��Ye��Qi�o;e���Y�fhG��0�7W��C����ʾ����\�x��VA��������ؽ��ƽH/����½ǽdt˽��ͽp̽��ƽ*l��\:��U�������3���   �   ̯*��� ��T���;8��.Һ8c�;l!y<��<���<��<��<��<�v6<�ͬ����9�{�^�սh#���h��[��:�ξ�:��!�.H9���Q�
�d���p��(u�D�p���d���Q���9��5��1��hվ�i�����|�K��	!�����!�4rѽ:�ʽo�ʽ�5ͽ�]Ͻ��ν�ɽ�����	����������|�N!T��   �   �����$�������`k�:��)<�J�< ��<�V�<v��<�%�<B��<�><���"��3%���ؽ�`%��Gl�Ϡ��/ҾgT��� �RR<�%�T��qh�B�t�,<y���t���h��5U���<��!��t��پoR�� \��jO��#��X�fE��սv�ͽ�OͽXiϽH�н�AϽzyɽ~;������柽ܝ���(p��E��   �   7�*�m� �T���:8�`'Һ�d�;8"y<��<2��<t�<���<��<Dy6<0Ǭ�Z���{�@�ս�#���h�M[��X�ξJ:�=!�eG9�ҁQ��d���p��'u�A�p���d���Q���9�65�1��gվ�h�������K�!	!�0��� �qѽ(�ʽX�ʽ�4ͽ\Ͻ��ν�ɽ!���7	��0��������|�� T��   �   SY�\m0�X�L����A�@���;l{q<f�<r~�<�Ͼ<�i�<��<���&�缬�r�*Dͽ�9�j�^��J���ožQ��+��vw0�|}G�ʰY��We��Oi�9e��Y��fG���0��U��A����ʾP����x��TA�������bؽ��ƽ3-��z�½ǽlr˽ȇͽ�̽��ƽ�j��9��A������Ƹ��   �   �딽,`���(W�%4(�lG��T���	ֻ��I;�/<��<N�<Шn<���;h��t���e�?�������QO�\m��ն���V���"���7��H��:S���V���R��!H�b7��a"�������.��DȒ�gd��0�V_�J�㽟MŽ||��R��Dᶽ%P��Xnƽ�ͽ��н�}ѽݸν��Ƚ����Q���諒�   �   ��н���`��n}���X_�b$���ּ��_�ЫN����;�@
<\<`';p��2 ޼��W��α�wn��X<�f�}�!���&ξ��T|��($�H�2��C<��W?�y�;��2�~#�!T������̾�)���
���I����L�����ǽr���I1�������P�������h½�Ͻ��ڽ� �d7꽊9�z�콛��ݱ޽�   �   ƀ�<�� ���Ͷؽa��@*����V�e���N���+��7\�@��e}�DSN���n�K�ˢ��e�	�'��j`�����Q���F�ؾ a��*�U��(q"���$���!�4=�>����_$Ծ�����q���.^���+���XDν<��X��t��������]��R���kU׽K��(f ��\	���"��������   �   �nG���>�b0��~�,Y�T߽�Q����6����z���8�L�0I����~����D��̕��u׽���#C�&�x� ���
·���Ծ����~� ����	�������:��ξ����}���|i���6����ս��������o��l�t~����������ƽ��潝L��G�P�%�&&4�r�?�[�G��ZJ��   �   2���[J���q�*}Z�pl>�Z���� �>�ǽ���~S��S�r�ټʔ���\ϼ�Z
�[�E�L����½z�nU(��PS�|р�a����Q���_þ��Ҿ�\ܾ��޾6�پ�;
����J���͌��g��9�����ٽ����K {�%`M�k<��1D���b�dF��"I��c�ҽd����K���1���J�c8b��v��@��+����   �   #����F���<�����������X��_1��	���սܞ�KPi�� 0������##��rO�)�������~�ӣ��2���U�څy����^T��rw��l�L��C��:��*�������X�\\1� ��սZ؞�^Ji���/����@��!#�zqO�,�������r�����2�m�U��y������V�� z��,��   �   �޾l�پ��;愻�kM��Ќ���g��9������ٽ����p%{�;dM��	<��3D�I�b��F���H��m�ҽ����PJ���1�E�J�+5b�v��>������͸���G����q��xZ��h>������ �S�ǽ����wS�ON�>}ټx���XϼY
��E������½m��V(��RS��Ҁ�3����S���bþ��Ҿ`ܾ�   �   @�	�|��Y"���=龜ξk������3�i�J�6���j�ս����D����o�rl�v~�@������ƽ��潖K�F�O�%��#4�p�?��G��VJ��jG��>�@^0�N{��U��	߽M��Ӏ��;�6������|�L��%I��������D�@͕�Nw׽����$C���x�����ķ��Ծ���l������   �   ��$�f�!��>��?�j���&Ծ ï�Ds��x1^� +����Fνg�������������]��<����T׽��e �L[	�-��ڸ�B��&���}�2��4���5�ؽ�[���%����V�Ʋ��C��l�*���[�@k~�0E}�NN� ����K��ˢ�hg�7�'��l`���������G�ؾlc�������r"��   �   �Y?��;�2��#�kU������̾]+�����ڪI�M��������ǽ����2������Q��� ���h½ʆϽ��ڽZ��\5��6�'����罢�޽y�нE�����0y��Q_�"[$���ּȘ_� hN����;L
<�<�?;�����ݼe�W��ϱ�,o�Z<��}�A����ξ���t}�*$���2��E<��   �   E�V�&�R��"H�:c7��b"���Y��<0��Sɒ�d�U�0�_`����OŽ�}��Q��ⶽ�P���nƽ�ͽ��н�|ѽ��ν�Ƚ?���tN���쥽f蔽�\��M"W�.(�0<��J����ջPJ;p�/<*��<R�<�n<P��;���T�h�e����h���RO�n���ն�Y�����"���7�S�H�6<S��   �   �Pi�|:e��Y��gG�ͣ0��V�C����ʾ���a�x��UA�e��T���gؽ��ƽ�-�� �½�ǽ�r˽�ͽ{̽��ƽ�i��8������\�����iY�Ri0�S��ﵼl�@���𺐣�;(�q<h�<Ё�<zҾ<�k�<��<��������r��Dͽ�9��^�PK��]pž�Q�����x0�>~G���Y��Xe��   �   u(u���p���d�.�Q�R�9��5�r1��hվOi��Y���K��	!����6!低qѽ��ʽ��ʽ5ͽ�\Ͻ��ν�ɽ��������������d�|��T�^�*�{� �*P��38���Ѻ�q�;�'y<V�<L��<�<֩�<��<�z6< Ŭ����{�\�ս�#��h�}[����ξz:�|!��G9�0�Q���d��p��   �   [�-�+�*�9�!�l��v��39㾮�������8����R��2�q��h����W��M��%�(�*�� -���*�J�#��y#	�κ�L�ʽꦥ�|���r�?��D��$���_���0�;�s<t�<��<a=�=��=���<fB�<�2�;�RU��<�5�������#��'`���Z���߾u�`6���!��*��   �   ��*���'�I4������g߾v~��
^���|��<O�X�.�/������?��t����v"��l(���*���(�H"�AN�8��A���̽�̨�����d�H��U���Q ��aO;��N<J�<
��<,��<fS=�;�<t��<Tؒ<p�;��X�x���n��B,�	"��2]�-y������Kܾ�� �����3�N�'��   �   �p"���4f��
������TԾ�)��F����Po��D���%�ʊ��4	�}����H�] �2w!��$���#����4����U��q�ӽ�����(���e��K*���\�}��L�����;��j<��<f�<4��<���<I�<�́<�i;X e�S���K����ٽRd���T�����ǭ��iҾ�����
�������   �   h����'?��R���Tþ��������b[���3�������_����{��N� ���������_�5>��B����3	������ཤ�Ľ�|������V`���)�d��4��PY��hք;sD<|m�<ƪ�<��<�:�<vF<@ R:��~���?����Ͻ��M�G�e��y����4þw�㾄^ �����%��   �   dP��������V㾆Vɾ�9��`&���pn�N�A�ղ��J�����ܽ��ڽ��㽖�F4��H
�hn��������0�����Q�FZ����ὤ�ʽ�1��N_��{��iD�K[������/� �w�P��;�@<�`<T�E<X��;�6i�HƖ�
���у��}ŽM
���8���l��풾�T����̾_*�����Y��   �   EW澇zᾲ^վfBþ/������� �x�	�K��%��a�ۭ�vbŽ�1��(���F�ýr�ӽb�潆��(~���LT�P������"��`���A���d���Ͻ�������}.r�b�5� ���������� �o��X:;��7; ����~!����Gj'�8������� ��(��zU�O傾ಛ�:���L�ȾQAپ|��   �   �(��Ё��#�}��O��� 'v��!M��,'�7��Vٽ�H���ŝ�������Y���>���ʽLW�V=������������ܿ!��}#�(�"��s����R���=�ܽ.޸�|:���a��!�^ټ.L����0������;�Ra��ڽ�i9�����[����@7�z?��hf��/���C�������ҷ�A����   �   ƚ������Տ�jЂ��Af��LD��y"�D.�>�н>��b���ʾl��0a���j��ׂ�~7��v����ͽ�3�F��Z���p"�1�/�;��C�(zH���H��D�b6:�Y�+�)�����`/ڽ��������F����3޼x���ļ.�w�"�U��܍��Ʒ���1��"�+�vRJ���h�ﮂ�����(��Z@���   �   �{���q�D�a�Z�K��1����M��p�½�U��;�j��;�IH"�u��N-���M�l�|��.���̌彤��;J�\3�8�H�d\�8�l���w��}��{�d�q���a�ʠK�2�1���ZR��x�½0Y���j�)�;��L"����-�>�M�F�|��/����Ќ�D��fI��Z3�O�H��a\�A�l�r�w�}��   �   �D�'3:�3�+�4�����*ڽ���&���t�F����*޼z�����ü��gt�
�U��ۍ��Ʒ�������O�+�3TJ��h�d��������*��uB������
	���׏�T҂�fEf��OD�;|"�p0��нb�������l�-5a�Ŭj��ق�99����ͽ4�3������o"���/�%;���C�cwH���H��   �   $�<P����X�ܽ�ٸ�y6����a� �!��ټ2C���0�����;�T\����?h9�Ԟ��\����-8��?��jf�
1��aE������շ�����+��"���X�����!���D*v�Z$M�
/'���HYٽfK��tȝ�P�����[���@���ʽ�X�R>��ũ���������p�!�&|#� �"�5q��   �   �`���Ͻ�󴽺���G'r��z5�z����p��@�n�Ћ:;�8; ���<w!����i'�J��������� ��(��|U�h悾E���횳�C�Ⱦ�CپV~㾥Y��|��`վnDþ����2�����x�:�K��%�|c�����dŽ,4��b���k�ý��ӽJ��2���~�L�hT��O�!����з�à��=���   �   �.��<\���{��cD��U�����/�@�v�(�;��@<��`<��E<���; "i��Ė�����у�g~Ž�M
�Ô8�0�l��V����̾@,�����Z��Q��������8�0Xɾm;���'���rn���A�?���K�8��ܽ��ڽ�㽙�95�~I
�o�+�����0�R��Q�sX�����ʽ�   �   ����R`�L�)����4��H<�����;4~D<Xr�<���<��<�=�<�zF<@UR:H�~�'�7@����Ͻ`	�Z�G�!���n����5þ��T_ �i���&�Z�� ��@��T��%�⾄þ���]����c[���3�������%����}��,� �����������_��>��B����z3	���ȿ��Ľ�z���   �   A�e�I*�X��8�}�P7�����;�j<��<��<���<���<�J�<ρ< i;��d����<L����ٽ�d�]�T������ȭ��jҾ���G�
�T�����jq"�����f���
������UԾ`*��أ���Qo�ҠD�z�%�t��$5	�"��W��H� !��w!���$���#�V���4������󽺹ӽ����'���   �   �H�T��를�K �vO;��N<��<��<���<T=�<�<8��<�ؒ<�;d�X�Ż��n���,�i"�#3]��y��t���*Lܾ:� �����3���'��*���'��4���"��Jh߾�~��L^��2|�\=O���.����D���?��t�_��pv"�Am(�0�*���(�5H"�ON�4����7�̽̨�����   �   L�?�}D��$��P_��H1�;s<&t�<��<V=�=��=���<JB�<�1�;�SU��<�d���̍⽥�#�(`����[��6�߾��k6���!��*�[�-�%�*�2�!�b��j��9㾕�������8����R��2�q��h����c��M��%�3�*�� -���*�F�#��m#	����4�ʽԦ��f����   �   �H��S��ꥼPJ ��{O;��N<��<f��<,��<TT=x=�<���<�ْ< �;��X����(n���+཮"�+2]��x������<Kܾ�� �G��L3���'�K�*�G�'��3�I����Qg߾�}���]��|�j<O���.�ɧ����4?�.t�����u"�xl(�g�*��(�~G"��M������Y�̽T˨�t����   �   ��e��G*�L���}��2�����;��j<\�<j�<���<���<<L�<�Ё<�,i;P�d�J���J���ٽ~c���T�y���ǭ��hҾ����
���c��p"�_���e�p�
�|����SԾ�(�������Oo��D���%�	���3	�����
�@G���Nv!��$�x�#����f3��������ӽ�����&���   �   ����P`���)���꼀���6��P��;|�D<�s�<(��<"�<V?�<�F<��R:��~��
�>����Ͻh���G�~~��g���e3þ�㾴] �����$�o����:>�>Q��2���þ������`[�u�3�}�����b���z��B� ����~������]��<��@�ܲ��1	�h������>�Ľ3y���   �   -��#[��<
{�lbD��T�f���4�/� �v�x�;T�@<T�`<�E<���;�i�������Nσ��zŽeK
���8�J�l�c쒾2S��2�̾d(澬���X�;O�v������L㾯Tɾa8��%���nn�a�A�9��"I�m��zܽK�ڽj�����2�G
��l��������.�v���O��U��x}�"�ʽ�   �   b_罖�Ͻ����1&r��y5������|�� �n��:;`+8;@��,n!����Le'�`���Ĉ�� � �ƭ(�KxU��ゾ���@����Ⱦ�>پ�y��T�	x�T\վ4@þ7���靔�*�x���K��%�&`�ªཟ_Ž$/��l���`ýU�ӽ������|��
��Q��M��*��W������;���   �   ^��O������ܽ(ٸ�
6��3�a�J�!�vټ�A���0����x�;��W��v���c9�՛��X������4��?�pef��-���A�������з����0&��O���ﱾ�z��V����#v��M�B*'���gRٽ\E��������얽�V���;��ʽ;S��8����b���������!��z#��"�:p��   �   �D��2:�Á+����Ì�.*ڽ���ʶ����F����(޼������üf�Kq���U��؍��·���罠��>�+�/OJ��h�ꬂ�����|&���=��Z���~��Xӏ�P΂�1>f�_ID��v"��+��н���0��l��*a���j��Ԃ�4������Zͽ�.뽪��|���m"�ͱ/�w;��C�?vH���H��   �   2{��q��a��K���1���MM���½lU����j�.�;� G"����<-��M���|�,���쾽.�彰���F�xW3���H��]\�*�l�$�w��}�f{�8�q�%a���K���1���[H���½�Q��w�j��;��B"�����-�łM���|��*���뾽�����:G��X3���H�)`\� �l�k�w�I}��   �   �������tՏ�KЂ��Af��LD��y"� .���н�������ͽl�d/a�Ҧj��ւ��5��!���{ͽy/뽯�����l"���/��
;�ҙC��sH���H��D�Y/:��~+���� ��@%ڽ?�����m�F�[��޼��~�ü�n���U�8؍��·����&��?�+��PJ�5�h�I���{���a(��@���   �   �(��������|��=����&v��!M��,'����UٽBH���ŝ�n����X��|=���ʽ�T��9��d��O��7����Z�!��x#��}"��m��	�M�����}ܽ�Ը��1����a��!��ټr8��h�0�����;��R��H��Lb9�h���(X�����5��?�;gf�/��8C��b����ҷ������   �    W�jzᾞ^վVBþ"��������x��K��%��a����bŽn1������p�ýL�ӽ���l���|� �R�\M���L������d8���[罇�Ͻﴽ ����r�js5�L���T䓼����m���:; X8;`2��4f!��
��Od'�6������|� ���(��yU��䂾`���ј����ȾAپ�{��   �   XP��������M�|Vɾ�9��X&���pn�9�A����pJ���꽐ܽF�ڽT�㽴�3��G
�Zm�P��(���.�@���N�T��R{὘�ʽ�*��$X��,{��\D�<O�>����/�@�u��1�;�@<0�`<�F<��;��h�ȼ��Q��Rσ�M{Ž�K
���8���l�N풾bT����̾"*澤���Y��   �   `����#?��R�����Mþ�������|b[���3�����������{��� ����D��Z��X^�>=�YA�
���1	����������Ľ}w������L`���)�^�꼆��X��H�;��D<px�<h��<��<tB�<��F<�S:�~��
�">��"�Ͻ����G���,���e4þB��o^ �w���%��   �   �p"���3f��
������TԾ�)��C����Po���D���%����j4	�^�����G� ��v!���$���#�I���3������󽒷ӽݺ���%��/�e�1E*����x�}�@����;4�j<�<��<t��<:��<4N�<�ҁ<�6i;T�d����J���ٽ�c��T�މ���ǭ��iҾ�����
����
���   �   ��*���'�I4������g߾s~��^���|��<O�R�.�'������?�wt����u"��l(���*�<�(��G"��M�������)�̽ ˨�����H��R�L襼0E ���O;d�N<��<(��<���<U=�>�<���<�ڒ<(�;��X�Z��!n���+��"�`2]�y��렵��Kܾ�� �����3�L�'��   �   zr龝w�nھ��Ⱦʪ��v���v����g��J�5�6�D�-��!/�H]9�J�8v^��0s�J���Θ���Ȋ�����,��O�o�\�U�<8��y��c��m��������7���м@/����;��{<�3�<<��<��=��=��=\c�<��<C<���H��Z7��8��\�޽1����G�)�z�ƍ�������Ǿi�پ�w��   �   h�徍���־�}žF���W��gʄ�Z�c�r�F��S3�g�*��,��*6���F�{�Z��/o��j���s��f�������<]����l���S�T�6����IX��.{��������<�D�ܼ(�.���<;hOb</�<Bj�<q�=f=
_=�$�<Х�<�M4< 1P��ޱ���8�����Yݽ���q�E���w�g�������ľ�}־���   �   ��ھ��־�̾%һ�u�������L|��iX��s<��*���!�4#�%�,���<���O�>�c���t�<H��8���@����v���d���M�y3�	�����/$½Zґ�
M�L�~�����<ё<N��<xu�<>��<��<���<n�<�<(��.����F=�����4ڽ���ݪ?���n�п���C��-5��?�̾E׾�   �   s�ɾ�žT໾AŬ��d��K���d�g��_F�>�,���R���>�.E��-�@	?�-�Q���a���m�4s��.q��4h���X���D��-�TJ�\8����ɽ؁���Lj�~�!���ü��)����:��'<Ά�<z��<@��<�ѽ<>��<��X<`�_;09#���޼�F��4���{ֽ�	���6�:�a�����V.��������Ǿ�   �   ����Hа�wx��%Ù��6��u!o��M�YW/��%�������Y�&����"�)���:�_J�UV��g\�d�\��V��#K��y;���(���� �<l׽�l������>GS�6���c��X�.�@6�a�;�J<�v<�0u<ܼB<X��;@�x����j��E�W�\7���XԽ�
�24-���R�"�x�����A����������   �   L��F��=����t��0�k�t�L��/�z�F� ����<۽žݽ���j����ъ!��`0�?L<���C�3�F��SD���=��3�� &���e7����+�̽�%��B/��t�Z�;� ��$ؼ<z�X�ϻ p 8�9j;�I�;@��:�$��t7`�(�Լ��(���s�`���Oֽ*��
<$�jC��b��)������?���	d���   �   ����r@��f�r��\�+�C��)�
�����.7н,���6ǯ��^���տ�a�ս�^���.�܎"�R�+���1���3�YV2���-�
�&�t������n����4ؽ����P7x�_�=���	�XY����{�`40�`��'B�,ԏ�:�ؼv ��*X�BP��/�����޽�����X6��[N�t�d�WJw�`o��慾�   �   �6^��T�Z�E���2�*��h�e��ʻ�aמ�x���C������w�������*���ݽ>����
��|�����&�F+��h-��H-�9�*�#&�������������ӽ�ᱽ
���xnd��0���	�����\Ӽ��݂�E-���\�芽|���y^̽f�ｊ�	����CM-���=�JtL��
X�Cz_���a��   �   �]6��+��#�����e��ʽ����W���)�_��LA�;�5�<��}S�>y�~���\ ��h�ν��콑��zP����x)���2��9��;>��~?���<�S`6���+�&�����i��ʽ��������_� RA�i�5�4<�ʂS�bCy�0������νL�콈��&Q�/���x)�)�2��9�':>��|?�d�<��   �   &�����i����ӽޱ�����Lhd�i�0�e�	��㼞SӼ~��V~��-�R�\��劽p����\̽��0�	�����M-���=��uL��X��|_�_�a�M9^���T��E��2������1"�Yλ�yڞ�V��sF��x��~z�������-���ݽG�����
�!~���C�&�AF+��h-��G-�%�*��&�S���   �   j���g1ؽM����횽1x���=�Y�	��O��Lz{��#0�`���B��̏���ؼ���-'X��N������Կ޽����Y6��\N�3�d��Lw��p��r煾	����A��R�r��]���C�7)�����V:н���ʯ��a���ؿ�y�ս�a񽼞���v�"���+���1���3��V2���-���&������ϒ��   �   ��̽ #���,��>�Z�D� ��ؼ�z�hmϻ /8`pj;8d�; ��:`���+`���Լ�(���s����Oֽ^���<$�kC���b��*��� �������e���M���G������<v����k���L��/�,��� ��罅?۽��ݽ�����������!��b0��M<�p�C���F��TD���=�+3�� &����6� ���   �   $k��춋�`CS�J��\����.��;5��y�;��J<��v<4;u<��B<ѹ;Ќx�|�������W�7��YԽ	
��4-���R���x�����h������i�������Ѱ��y��ję�8��z#o��M��X/��&�%����	[�}�����)�X�:��`J��V�0i\���\�'�V��$K�;z;���(���� ��j׽�   �   ̀��1Jj���!�<�ü��)����:��'<Z��<���<��<bս<ƿ�<p�X<@�_;�3#�b�޼c�F��4��Y|ֽ#
���6�F�a�����0/��
���'���LǾ��ɾV�ž|ỾRƬ��e�� ���ԉg�aF�c�,���^���?�RF�9-��
?���Q�B�a��m��s�	0q��5h�� Y�: E�e�-�\J��7����ɽ�   �   �ё�bM����~����@&<Lԑ<8��<$x�<ȝ�<��<���<p�<`<�������iF=����"5ڽ���x�?���n�Z����D���5���̾F׾�ھj�־�̾�һ�!��������M|��jX��t<�\*���!��4#���,���<���O�K�c�ët��H���������I�v�T�d��M��3�������#½�   �   >�����<�\�ܼ@�.���<;�Rb<�0�<�k�<"�==�_=�%�<���<\O4<�,P�bޱ���8�����Yݽ��טE��w�����b���u�ľk~־�������n�־R~ž����fW���ʄ���c�ٚF�gT3�Ҩ*�/,�A+6�5�F�
�Z�*0o�"k��t������죆�p]���l�S�p�6����,X���z���   �   ަ��h�7�0�м�.�h��;�{<�3�<j��<��=�=��=bc�<��<�C<`����1[7�9����޽M��հG�N�z�ٍ�������Ǿw�پ�w�}r龚w�cھ��Ⱦ����i���i����g��J�2�6�H�-�"/�[]9�6J�Qv^��0s�T���֘���Ȋ�����*��E�o�N�U�<8��y�zc���l���   �   ������<���ܼ��.�`�<;<Tb<D1�<Bl�<`�=H=�_=L&�<l��<xQ4<�!P��ܱ�p�8�����Xݽ6����E��w����������ľ�}־������ᾀ�־u}ž֩���V��ʄ���c��F��S3��*�b,�h*6�K�F��Z�/o��j��{s�����X����\���l�܏S���6����W��z���   �   eБ�oM��  ~����(<FՑ<*��<y�<|��<��<���<�q�<�<󷻺���D=���"3ڽ���ة?���n�&���&C��Y4��[�̾,D׾�ھ��־�̾Bѻ�����h����K|��hX�s<��*��!�I3#�`�,��<��O�@�c���t��G���������/�v�d�d�N�M�<3�������"½�   �    ��yGj���!�"�üܞ)���:t�'<���<ƫ�<*��<�ֽ<P��<X�X<@�_;�,#���޼3�F��2���yֽ\�K�6�~�a�����=-������»���Ǿ�ɾ��ž߻�Ĭ��c��V�����g�Q^F���,�Ј�?��s=�D��-��?���Q�=�a��m�ks��,q�3h��X���D�W�-��H�*5����ɽ�   �   	i��F����@S�q��RY��t�.�@5���;l�J<|�v<$>u<L�B<hڹ;�tx�J���͖�0�W��4���UԽ�
�:2-�M�R���x�;���̪��&��h��������ΰ��v�������5��1o��M��U/�$�z��H�rX�ʙ�.���)���:�]J�@V�oe\��\���V��!K�ew;�c�(�޸�� �Jh׽�   �   ��̽V!��N+��<�Z��� �ؼz� gϻ 280|j;k�;��:0���$`��Լ��(�u�s�����Kֽ���9$��gC�7�b�(��#�������Db��OJ��_D������Ss��h�k���L��/����� ����9۽׻ݽ����~�5��Ԉ!��^0��I<�]�C���F��PD��=�3���%�G��4�2���   �   ����/ؽ�����욽�/x�j�=�c�	�N��Hw{�� 0����B��ɏ�,�ؼi���#X��L��$���"�޽����V6�tXN�0�d��Fw��m��2䅾�����>���r���\�[�C�{)�՞����3н����&į��[���ҿ���ս�Z������e�"���+���1���3�lS2���-��&������S���   �   ����� ����ӽLݱ����Xgd���0���	�����QӼt��}��-��\�R䊽]����Y̽����	�׳�IJ-���=��pL�2X��v_�7�a�3^�|�T��E���2�p�����!ǻ��Ӟ�N���@�����xt��$����&��٤ݽ������
�2z�H����&��B+��e-�[E-���*��&�����   �   �\6�H�+�	#�5���d�$�ʽ�������x�_��KA�u�5�!<�z|S�<y�p���������νw�����jN�L���u)� �2�ý9��6>�y?���<��Z6�ٚ+�� �ۿ�s`�(�ʽ����������_��FA�u�5�7<��wS�o7y�����^�����ν������M����u)�w�2���9�68>�M{?��<��   �   �5^�H�T���E�'�2���0�ὡʻ�מ�$��TC��H��$w����)��˧ݽ������
�t{�P��]�&�GC+��e-��D-��*��&�@��&������󽋫ӽ�ٱ�����ad���0���	�����HӼ��⼶x��-���\�(⊽N���.X̽ ���	�ų��J-���=�HrL��X��x_���a��   �   3���.@����r���\��C��)���<���6н䕹��Ư�K^��Qտ���ս�]񽍜�����"�#�+�:�1���3�T2�!�-���&���ł���.���i,ؽ�����隽K)x���=��	�bD���e{�|0�����B�����ؼ���� X�K��ަ��B�޽��P���V6��YN�ȋd��Hw��n���兾�   �   �K���E������t���k�M�L��/�\�(� ���}<۽|�ݽj��4�����l�!�B`0��K<���C���F�RD��=��3��%��Y4�����̽����(��&�Z�ǻ ��ؼ��y��Gϻ `@8p�j;P��;�z�:ꔻ�`�H}ԼC�(�-�s���rKֽ��:$�VhC�y�b��(��:���м���c���   �   c���!а�^x��Ù��6��\!o��M�CW/��%����~��Y���{��)�j�:��^J��V��f\�|�\��V��"K�x;���(���� �Jg׽�g������==S�����Q��\�.��14�З�;��J<��v<�Gu<��B<��;�Px��������W�4���UԽ
��2-�/�R���x����ګ��`��û���   �   R�ɾ�ž@໾2Ŭ��d��B���Q�g��_F�-�,���@��n>�E��-�	?���Q���a�H�m��s�..q� 4h���X���D���-��H�5���ɽ(~��GEj�1�!��üT�)�`i�:��'<<䯱<���<8ڽ<�ġ<�X<��_;�&#��޼2�F��2���yֽ����6�I�a�g����-������μ���Ǿ�   �   �ھ{�־�̾һ�p�������L|��iX��s<��*���!��3#��,���<���O��c���t�H��������v��d�םM��3�
������!½�ϑ�0M�����}���\/<Fؑ<���<�{�<��<�< ��<�s�<(<0뷻����C=����23ڽ���4�?��n������C�� 5���̾E׾�   �   _�徆����־�}žC���W��dʄ�V�c�n�F��S3�c�*��,��*6���F�k�Z��/o��j���s��V�������]��o�l�.�S���6�!��;W��
z��n���@�<���ܼ(�.���<;LWb<�2�<�m�<��=�=X`=t'�<���<tS4<�P��۱�
�8�����XݽB�� �E�@�w�G���冮���ľ�}־���   �   �q����J.����Cr�>Z��tE�}�6��0�5��C�*�\�{�}�zG��V���س���aɾ��Ӿ�[׾�ӾɾG��������]��wh��9�,d��Ͻ*v��`�+����� �d�>< �<X��<,=�m=�=��<P��<�d<��*;(<?��5��K�Y����Ͻ���M�'�5�I��*j�zs��8Ď������   �   ?��<���ތ�߂�;n���V�B���3���-���1��{@���X�4�y�ԏ��ԣ�%����ƾ�GоV�Ӿ\eо�ƾ�赾�~��"�����e���7�Bl��#Ͻ�Ǎ���-��E�� Q<��n.<zf�<l-�<�3�<
�=8D�<e�<Tr�<M<@<�:�.V������,P�Ø���Ͻt�(�&�L�G��g�
с��ь��͓��   �   j��2Ό��.���y�̆b���K��G8���*���$�n�(�&�6���M�m�<����ɛ�����<����Rƾ��ɾ��ƾd;���(���������Kz^��3�t�
���ͽg��у4�����x?�����;~n�<J��<T�<V~�<rc�<Fk�<Pa�<��<0�U�Zc���y���]��l��`�ѽ+���$$�0�B�_g`�7Jz��:��ʅ���   �   �$���K����w��ge��CP��";�.�(�*����Q���K'��<��Y��8{�A���៾ʣ��e趾`�����\����N���5����{���S��,��T��c̽�d����A�p�ݼ�Z.�p�; %C<X��<�A�<�ܺ<�&�<�܈<4�"< �9:М2��̼&)��%v�\����ֽ9R��� ���;���U��Al���}�j�   �   ��p�6lj�@�]�:�L��9�C�%��A��	�����J����&���@�: _�,�~��d���ѓ���L��y����잾)��H����i���F� �$�cP��ͽh]��	�W�
�䊔�H����};�z(<\`<8�h<pD<���; ���}&�j^��<����T��d���ε��Nདྷ��Ǳ��q4���I���[��i�map��   �   h?U��M�A�(�0�O�e������X�(�཯�彉	��z��[�$��?�%�Z�H�u����)���
��w���������eq���V� �:��d�2<���ӽ��`�y�12����D������@�� �.;p�9; (��������f���ʼm:��\S�\3��U�����ͽ̟��@=�u�.�)>���J��zS�^-W��   �   �9�h�0�l�#��w���轠�νyP�� ���Y���,ʽ�*罝����v�5��7M�fa��}p��y�;�z�u>u���i�r�Y��FF��	1�*�?���V��(X��Gh�3-���������0�i� '6��:��Qu�Q��7� ���1���i��-��g��y�ѽ���W���C�e� ��,�q[5�<�t]?���>��   �   $� ����$;�pi��ӽ�m��䟽-���襈� ���R������!�ӽF������>&�r8���F�ԥP��U�
YT���N��E���9���+��X��N�������ֽb
��ܦ���as��A����&#�����\A缛E���'��V��+�����Uǽ��潘4��E�T��?#��*���.��1��31�ڮ.�Q)��   �   �����ZL߽���-£�nd��u�g�b�J��n=��?B�{Y�p���*����f��94὜��#^�(�!�l�,���4���8��a9�D-7��u2��+�7�"�Q>���Ծ��FO߽���ţ�<g����g���J�?t=�lEB�܀Y�� ������wj��Z8�Ν�b`�b�!���,�d�4�:�8��b9��-7�5v2�Ŗ+���"�W=��   �   $���ʮֽ���\����\s�$�@�������H�ἤ7�r@�.�'��V��(������ǽ9���2�D��R��>#�*�F�.��1�741�ѯ.�dR)��� �4���<��l���ӽ�p�� 矽 �����������U������ӽDJ����tA&��t8�e�F�G�P�(U��ZT��N�$�E��9���+��X��M��   �   �U�cﹽDV��Ch�-�l�������<�i��6��:� @u��G��� �O�1���i��*��d����ѽF��P��C�� ��,��[5��<��^?��>���9�8�0�;�#��y���4�轞�ν^S��坴�V���/ʽj.罘�#����5�':M��ha�U�p��y���z��@u���i�ʯY�jGF��	1�*����   �   ��ӽ�𥽘�y��-2�H�鼴���@������.;��9; 0K�P����f���ʼ�5�4XS�1��<����ͽv��Q�9=�Ҋ.��>���J�Q|S�/W�6AU�ϥM��A���0�����{���'���བ�彮��6��T�$��?��[��u�%�����M��Ą��%������fq���V�î:��d�<��   �   ��ͽ�\���W��|
�����8�p~;��(<�f`<4�h<�D<��;�a��p&�tW�����0�T�*c��j͵��M�x�����]r4�ӗI�&�[��i�	cp�]�p��mj� �]��L�- 9���%�DC�N�	�'��l����0�&���@�L_�y�~�f����+���%N�������ힾÓ��I����i�j�F���$�tP��   �   �c̽d��a�A�@�ݼ�S.�@�;d,C<���<�E�<d�<�*�<�<d�"< Y::�2���˼�#)��#v������ֽHR�
� �~�;�d�U�Cl��}� ����%��^L���w�ie�+EP�$;�K�(�&+����m��-M'�}�<�x�Y�N:{�
B��㟾줭��鶾����(��R����O��|6����{�Z�S�. ,�U��   �   ��ͽ���4����� 6����;�p�<¹�<�!�<ހ�<f�<n�<dd�<��<��U�x`��>x���]�dl��Q�ѽL��G%$���B�	h`�Kz�d;��Q����j���Ό�=/���y���b���K��H8�P�*���$�B�(��6���M�Gm�巈��ʛ�{�������Sƾp�ɾ��ƾ<���)��i	��\����z^�3���
��   �   �#ϽqǍ�	�-�XD��G<�Lq.<�g�<�.�<D5�<��=�E�<�f�<�s�<�M<�Q�:X,V�b���^,P�Ø���Ͻ"t�a�&���G�S�g�Jс��ь�@Γ��������Wތ�W߂��;n�.�V�tB�7�3�j�-��1�&|@�6�X��y��ԏ�գ�����^ƾHо��Ӿ�eо�ƾ鵾�~��N���2�e���7�Fl��   �   ��Ͻv�� �+������ ���><b�<���<@=�m=�=2��<���< �d<0�*;P<?��5�?�K��Y����Ͻ���f�'�M�I��*j��s��@Ď������q����E.��
��Cr�>Z��tE�|�6��0�15�!�C�K�\���}��G��i���쳹��aɾ�Ӿ�[׾�Ӿɾ>���|���}]���vh���9�d��   �   �"Ͻ�ƍ��-��B��`=<� s.<~h�<:/�<�5�<��=F�<g�<bt�<h!M<�a�:�)V�����B+P�U��Ͻ�s���&���G�W�g��Ё�1ь��͓����⡓��݌��ނ�z:n�5�V��B�d�3���-�N�1�F{@�>�X�ǁy��ӏ�Iԣ�С���ƾ&Gо��Ӿ�dоƾH赾C~������7�e���7��k��   �   ��ͽ���Ԁ4�d����,�� ��;Rr�<ܺ�<�"�<���<�f�<�n�<�e�<`�<p�U�^���v���]�k����ѽ2���#$��B�.f`��Hz�@:�����ri���͌�.���y���b���K��F8���*��$���(�`�6��M�*m�����3ɛ�����r����Qƾ��ɾ�ƾ:��(����@����x^��3�`�
��   �   a̽b��k�A���ݼ\M.���;�/C<���<�F�<��< ,�<R�<��"<��::؍2�d�˼�!)�� v��}��N�ֽ�P�/� �D�;���U�"@l��}�t�#���J��Ȭw��ee�YBP��!;���(��(����C���J'���<���Y��6{�'@����������2綾 ����
������M���4����{�ɂS�,�mS��   �   ��ͽTZ����W�)z
�����嶻�~;��(<�i`<��h<�D< ��; Tk&�rT�������T�aa�� ˵��Jཤ������o4���I���[�7�h�_p�K�p��ij��]�<�L��9���%�j@���	���������&��@�I�^���~��c��D_���MK��򬥾)랾�����G���i�Y�F��$�xN��   �   ��ӽ-��y�+2����^���0��@����.;�9;  ?������f�l�ʼ4��US��/��L���d�ͽJ��S��:��.��>��J�>xS��*W��<U�m�M��A���0�P����9���I�:~����t�����y�$�e?���Z���u�B�����?	��ǁ��R���x��bq��V�p�:�.b��9��   �   &Rώ칽BT��P�g��-���� ���8�i��6��	:��<u��E��� �	�1���i��)���b����ѽ��ｴ��A��� ��,��X5�: <��Z?���>�U�9�ȷ0���#��u�	�F��-�νHM��񗴽F��t)ʽY'罥 ������5��4M��ba�Bzp�py���z��:u���i�'�Y�lCF��1�R'�����   �   ׻��A�ֽ����Zs���@����������*6缳?�R�'��V��'���~���ǽ����1��B�Q��<#��*��.��1��01��.�?N)�f� �����8��d��ӽ&j������ ���࢈����tO��,���@�ӽ�A��D��@<&�o8���F�u�P�xU��UT��N���E�I�9���+�V��K��   �   &�¹���J߽���8����c��[�g���J�9n=�L?B�XzY��������f��3� ��~]�O�!�T�,�$�4��8��_9��*7�s2���+���"��:�������G߽���T����`��	�g�_�J�/i=�,:B��tY����t����b���/�
��S[�!�!�>�,�>�4�X�8�m^9��)7��r2�ݓ+�6�"�q;��   �   �� ����`:�Th���ӽ8m���㟽ũ���������XR��N�����ӽ�E��j���>&��q8��F��P��U��WT���N��E���9���+��U�@K�2���0�ֽ��������Us���@�������}��,��:��'�V��$��V{���ǽ"��0�.A��O��;#��*��.��1�11�ˬ.�tO)��   �   ��9���0���#�_w���~��6�ν"P��������h,ʽ�*�r����2�5�/7M��ea��|p�y�B�z�9=u�c�i���Y�mDF�'1�t'����Q�E빽�R��v�g��-����F|����i�86��9� ,u��<��=� �̍1�b�i��&���_��̉ѽ�ｚ��D@�%� ��,��X5� <��[?��>��   �   �>U�K�M��A���0��2��8������v��L	��X��:�$�`?���Z��u��������
���������}���cq�;�V�=�:��b��9��ӽ<�@�y�,(2����4���`�� ��./;0:; ��(f��@�f���ʼ�/�iQS�P-��%����ͽΙ����:�"�.�(>���J��yS�F,W��   �   ��p��kj���]���L�l9��%��A��	���� �4��z�&���@� _��~��d��������L��0���N잾����dH��?�i�A�F���$��N���ͽ�Y����W�+x
��}���Ҷ�p9~;0�(<@s`<��h<*D< ��; g��D^&�|M��B���T��_���ɵ��I�g��˯�p4�o�I���[�� i��`p��   �   �$��pK��O�w�nge��CP��";��(�*����@���K'��<�іY�q8{�A���៾����H趾:����������N��p5����{���S��,��S�Ha̽�a����A�N�ݼTG.�� ;�6C<��<XJ�<*�<�/�<n�<P�"<@-;:��2���˼/)��v��|����ֽ�P�T� ���;�z�U�Al��}� �   �   �i��Ό��.���y���b���K��G8���*���$�e�(��6���M�m�4����ɛ�����1����Rƾ��ɾ��ƾ<;���(����������y^�3���
��ͽ���t�4�����%�����;bt�<���<�$�<��<Zi�<�q�<Fh�<x�<`|U��Z��u�@�]�~j��@�ѽ*��$$�^�B��f`��Iz��:�������   �   .��0���ތ�߂�;n���V�B���3���-���1��{@���X�-�y�ԏ��ԣ� ����ƾ�GоL�ӾNeоpƾ�赾�~��������e�7�7��k��"Ͻ�ƍ��-�TB���7<��t.<Zi�<"0�<�6�<v�=,G�<<h�<�u�<p$M< {�:x&V�����*P����Ͻ�s���&���G���g��Ё�hь��͓��   �   �mB���?���8�CM/���%��Z�*~��"�G�2�i�N���v��/��������Ծ�x����
�2������!�>�����4
�����-Ѿ�¬������S�z��X�ؽ8؊�?���\e�p�i;�Y�<���<��<P��<���<x?�<ڨ�<�?<��;�t��Ƶ�p���Z�-`��A��E��4�k��3y*�̎7���?��   �   ��?��=�(�5��z,���"�[�� �����i�/�y'K��r�L�������<qѾ�_�>�R`�FE����N�`�\�>���ξ�K���凾h�P����@�ֽ
��}����j��8F;�	{<�߾<�<�X�<���<f��<>:�<T�< P�U;�4�ȼ�| ��c��ɕ�䆼�/���L�o
��M)�?�5�D�=��   �   `�8��#5���-��U$������]������&��@�Ozf��k��h���M&Ǿ�}澎���&�A���]�A��a�z��� �kž6������I���JJѽ�����i��|����:D�V<��<��<"u�<*ֺ<t)�<x�@<p[;�޻�~���f�p`<��c|��~��w�Ľw~�6����&���0��N7��   �   c�-�x()��T!�����l�՜����S�
�����0���S����e�����
�Ӿ�n����Pw�BE	�ƌ�����<վ�B���a��'u��[>����ɽ����7i�v@����|s<�Ё<�;�<���<��{<� <p9	;�V��Ŗ����P�3��5m�����ѳ�1�ӽ�>�����$�!���)�`.��   �   5� �֔�y��T	�F|��:
�,��؁������J�)Z;��Bc�T&��*ʢ�k����9Ծh����j����s������׾ob���0�����֨a��'1��J½����Z�$�U��(Tۻ�DN;��<��/<L�<࿗;�%�B����y��zF�,~��������n�ѽt�뽋)��L����3��p"��g#��   �   �V�4�;'�*`�,fڽ3�̽��ǽ��ν�����e��BzB��Pk��勾�D��+Ӷ�ؚǾ��Ҿ<�׾�վ��˾�Ӽ�k���ࡓ�0�y�	<M���#�L]��4ټ��S���%3�\�ؼ�W_��襻@� r�5O��}�(뙼:���(�2�Z]m�ح�����ͽ���T������"����G��f�1���   �   �P�C���P�fʽ�i���������Ȧ��J����׽���� ��B�77h����l��Y䦾�Ӱ��Z������P���ơ����^U��.5^��+:�b*�El�"������J�������N�� �M�\�^��T��Zl߼�y ���[��)������sԽ
a��+�j����_!�B,$��z$�b�"�������J���   �   t��	~߽��ý����"��,Y��iuy�&�}�r���R����˽�&������9��)Y�_v�Xh���)������sƔ����'y��, {�ȅa��F��k*�����������)�l���5����$�꼐)ݼ���҅��fF��U��̊��ڙнT�����]�#�u-2��q<��B��9C�@E@��9���0���%� p�F��   �   ^��_s̽�쪽]e���Kj�G���3���2���E��m��䔽���}�H���f(���@�wU�I*e��n�R�q�M�m�m�d�@�V��E�3��P�ʗ����nt̽`g���Oj�!G�S�3�`�2��E�!�m�蔽����������i(�ޮ@��zU��-e�c�n���q�G�m���d�C�V���E�3�IQ�֗��   �   ����������v�l�^�5�|��n��,!ݼ��d��y`F�RR������,�н���2��i�#�s*2��n<��B�?7C�>C@���9���0�T�%��o���~���߽��ý�é�D
��k[��1zy�O~�Q������t�˽+������9�W-Y��bv�Rj���+������[Ȕ������z���"{���a�-F��l*�P���   �   �l�꯻����ߔJ�8 ��y��4H����M��^�dK���a߼�s ���[��%��x��JoԽ6\�����g�����]!��*$�sy$���"�E��ˢ����|Q����R�Ghʽ�k�����b��w˦��M��T�׽��� ���B�`:h��
��h���u榾�հ��\������R��Oȡ�u���sV���6^��,:��*��   �   �]��Lټ�PS��L$3���ؼ�N_��ӥ��`� �d�P�N��k�>ᙼ ���д2�}Vm�0��� ���ͽ(�� ���.������F��f�����eW�.�N(�nb�hڽ��̽j�ǽM�ν�佒��Y���|B�xSk�=狾xF��+ն���Ǿ��Ҿp�׾վ��˾Yռ�ׄ������y�8=M�B�#��   �   t�eJ½����v�$�hR���FۻdN;��<��/<\�<Pۗ;��$���A�^����s�fuF�p&~������-�ѽ����(��L����r�Tq"�Mh#�� �ϕ����h
�q~��p�p��>������6L��[;��Dc��'���ˢ�����;Ծ�j����~����u��|�龃�׾�c���1������a�w(1��   �   ��&�ɽ��h��>�����`y<ԁ<X?�<H��<ȗ{<* <�l	;�:�\������]�3�2m�X���:г��ӽ�=���+��w�!�|�)�.�0�-�V))�nU!����{m����t��R�
�%��E�0�.�S����3f�����Ӿ�p�n�����2x�F	������$>վ�C��Hb��-u�;\>��   �   ���Jѽ����(i�4|�`̫:0�V<D��<���<x�<�ٺ<0-�<�A<<[;��޻�y��$d�^<��a|��}��ڒĽ$~�5��:��c&�#�0�DO7���8�.$5�G�-��V$����R����@����&��@�z{f��l��=���C'Ǿ�)��3'���y^�����a������ž�6��z����I��   �   ��J�ֽ�	��/�� �j� @F;{<��<f�<ZZ�<\��<b��<n<�<�< ��,P;�ַȼ�{ ��c�Jɕ��������L��
��M)���5���=� �?�%	=���5�E{,�
�"����_�����/�(K�ԕr���������qѾr`��>��`��E�0�5O�h`������7ξ-L���凾��P��   �   Z��$�ؽ
؊�����[e� �i; Z�<4��<R��<x��<2��<�?�<�<L�?<@�;�t��Ƶ�p���Z�C`��^��,E��4�y��By*�؎7���?��mB���?���8�DM/���%��Z�3~���"�b�2���N��v��/��������Ծ�x����
�?����ī!�>�����4
�	����-Ѿx¬�����̎S��   �   d��A�ֽ9	������j��IF;�{<l�<	�<�Z�<���<̌�<�<�<�< ��dN;���ȼ�z ��c��ȕ�腼�1��eL��	�M)���5���=�G�?�M=���5�yz,�I�"�������Y���/�&'K�Ôr����W����pѾg_�N>�`��D����N��_�	����XξuK��`凾��P��   �   v��Hѽ9���g��|���:P�V<���<���<�x�<4ں<�-�<�	A<pD[;h�޻�w��c��\<��_|�~|��a�ĽZ|�&����&���0��M7�b�8��"5���-��T$�J��������ә�k�&�J�@�oyf�Pk�������%Ǿ}����%����1]����``������pž/5��b���ǂI��   �   ��b�ɽݣ���e�4:��`N��}<�Ձ<�@�<x��<��{<0, <pv	;05򻐼��`��ο3�	0m�����γ��ӽh;���{����!�l�)��.��-�')�<S!����tk�͛����Z�
� ����0�V�S����-d�������Ӿ�m����(��lv�]D	�����{;վ�A��e`��%u��Y>��   �   @�G½@�����$�M��(7ۻ�yN;��<<�/<�<X��;��$���A������r��sF��$~��������8�ѽ4��j'��J����+��n"��e#�e� �!��������y������n��\��HI��X;��@c�0%���Ȣ�ܒ��8Ծ�f����H����q������׾�`���.��\��f�a��%1��   �   *Y���ռ��P��N 3���ؼ\F_�xǥ��� �`���N�i��ߙ�p���߳2�KUm�p��������ͽx����������*��D�#d�����zT�@�o%��\�$cڽ]�̽B�ǽ��ν�V�����$xB�<Nk�-䋾�B��@Ѷ���ǾU�Ҿ�׾�վ��˾�Ѽ�p�������y�K9M�)�#��   �   �g�,���C�����J�6��lu�� E����M�T�^��I��4`߼�r �	�[�~%������nԽ4[����f�����\!�$)$��w$���"�ɋ�������N����@L὘bʽhf���	�����Ŧ��G����׽��l �n�B�14h���w}��2⦾aѰ�OX��g���N��uġ�����S���1^��(:��'��   �   ��O���0���w�l�m�5�V��f���ݼ6����_F��Q��I�����н����ծ��#��)2�n<��B��5C��A@���9���0���%�bm��
��
���y߽߃ýZ������*V���oy�i�}�x���
���˽["������9��&Y�V[v�If��l'��p���*Ĕ��}��w��){��a��F��h*�K���   �   ��p̽tꪽ�c��<Ij�G���3���2���E�[�m�4䔽o���|���Jf(�>�@��vU��)e�,�n�p�q�-�m��d���V�3�E��3�qN�C�����#o̽%骽�a���Ej�JG�r�3��2� �E�ӝm�ᔽ���Jx꽒��sc(��@�8sU�D&e���n��q�$�m�f�d�m�V���E�� 3��M����   �   ���#{߽��ýE������MX��+ty�=�}�������W�˽]&��\��Խ9��)Y��^v�,h��c)��i���Ɣ�w���x���{�!�a��F��i*�ž������K����l���5���@��ݼx��z�ZF��N��r���T�н����$���#��&2�*k<�B��3C��?@� �9���0�>�%�m��
��   �   ,O�ѵ��:N὾dʽ�h�����b��hȦ�`J����׽ո�~ ��B�7h����R��6䦾|Ӱ�oZ��y��pP��-ơ������T���3^��):��(�mh�0���͏���J���>p��
?��\�M�h�^�fA��tV߼3m ���[��!�����jԽ�V�����d�����Z!��'$�Wv$���"�r��"��D���   �   BU�8�~&�_�jeڽ��̽��ǽa�ν�����G��(zB��Pk��勾�D��Ӷ���Ǿu�Ҿ�׾�վ��˾FӼ�����X�����y��:M��#�1Z���ռ�uP��P3���ؼd>_����@l� U��N�Y��֙�ޑ���2��Nm�楔�^����ͽ�潾���r��c��b �(D�d�,�b��   �   ;� ���������{���	���뽚�������J�Z;��Bc�H&��ʢ�^����9Ծmh����M����s��r�龟�׾b��0��P��ӧa��&1����G½b���^�$�,K��,ۻ�N;�<��/<��<H��;А$�@�A�`����m��nF�~� ��񸶽ڽѽ7�뽫&�TJ����P�Fo"�Zf#��   �   ��-��')�$T!����[l����i��<�
�����0���S����e������Ӿ�n�����Hw�4E	��������<վ�B��@a��ou��Z>�F��ɽ$����e�,9��`3�<�؁<D�<l��<��{<�6 <��	;h�B����	��޻3�!,m�:����̳���ӽv:����w����!���)�z.��   �   �8�4#5�_�-��U$�������J��q���&� �@�Czf��k��d���G&Ǿ�}澌���&�=���]�:���`�l��� �@ž�5��☂���I���&Iѽ����2g�(|����:�V<:��<���<:{�<ݺ<@1�<,A< f[;��޻�r���`�#Z<��]|�v{����Ľ�{�����4&���0�'N7��   �   ��?��=��5��z,���"�R��������b�/�t'K��r�I�������9qѾ�_�>�P`�DE����N�`�V�,���ξ�K���凾+�P������ֽ�	��P���j��KF;�{<�<�	�<�[�<��<b��<�>�<(< �۷�I;��ȼ�y ��c�$ȕ�v���ޮ�OL��	�.M)���5���=��   �   q%���.�'Y����*���Aq�Q'���M�pɁ��}���ξNv�������1��qH�kwZ��f�Tj��f��hZ�T2H��.1��i�4���uǾX��$db�����Խ�π�����)�PO�;��<�̺<|��<��<8A�<�S<(��;�]S��"R��H��y�
��[8�}g�A��5���(��XMͽ�:޽��	��   �   e+�^��$#�,O�d4�ڲ��e��?$�ScJ� :����O"˾�:���)��.�D#E���V�Sb��Kf��[b���V���D��Y.������<ľ�ϖ��6_�f��R4ҽ��~�P���H�; y�<���< ��<�1�<J��<�c*<P�*;нлt����ټ_%��HF��	t���h��Ӟ����Ͻ�M߽L��X���   �   �����罰
�a޽�߽�C����	��XG@�Ǘr�ș��'�������[T&���;��uL��eW��8[��W���L�"�;��'&� �c��b���Y���V���@�ʽ'zw�Rf��������;\�e<�V�<�s�<�~<0�%<6;`@ƻ䆂���ؼ)��N.E��q�獽Ћ���	����ǽ$׽���꽀��   �   a>彊ݽ�|Խiν�zν��ؽz�����l0�;�^�4Y�������ھ�Y�E�Z�,�35<�lWF�]�I��F��<�-��m��b�xyپk����o���(H�P��\����.m�����4� �	;�z<4�I<��3<���; y���&�tx���N���4��Bd��Ĉ�H�������2���4&н�$ܽw:�B��"�콍���   �   ��ݽ�н�{Ľ�]��I���[=��СսǑ���&�۝E�V{����7�¾:��*������'�)�0�4�01�z(����ki	�"����þ�L���]t��7�����]��s�b�hu��d�^�`5$�вF;�r; �90��V ���v�,�ܪe�&��|������/�Խ|��i�m�������V��S����D���   �   2hٽR�Ž�M��7���ܠ�����.���l�ֽ�-�(�{DW�٘��LS��dɾo��Q��r��i�{j�&����`H�D!�Uξ�����ӿY���$�M����j�Z��6�ꯐ���pX»� ��ti���ȼ37��s[�롐��;��f\ֽ	���#��~��p�Q���c���D��
v�7����8��   �   *�ٽI1���+��^���z���@S��h���y��LJٽ�
�y�1�3�`������C���:þ��ܾ�<������e �m:��P�⾵�ʾ�Ư�Nܓ�h�q�O�?��Z�M۽�3��G�X�A�^��p��ʢ���{���=�{�>��у�?ԭ��ڽE��L��O+�K[9��hB��#F��D�ܯ>���4��u(��?�>'�h����   �   m`�nӻ��𛽼,���%f��Z��f�Sچ��٨���ٽ��x-3��^�(h��;�����E�¾RGξ�8Ӿ�DѾ�Ⱦs����*��j9��w�z���O�P�'��(�"�ʽ{h���V^��Q$�=� B�O� �v#���\�"l��HAŽ����m����7�AR�<Ch�:rx��^]��j�|��*p���^���I�`3�H��a���   �   ���>´�ܖ�:�m�BA��*��H*��OC�,v��k����ӽ(���^+��5P�%�t�H��귘��H��I覾�F�����������U���s�lVS�Y�2��Q�����࿽�ܖ���m��A��*��L*�|TC��1v��o��@Խݨ��a+��9P�w�t����z���MK���ꦾ�I��������W���s��XS���2��R��   �   R)���ʽ�h���U^�P$���d;�� ��p#�B�\�6h���<Ž���(���7�-R��>h��mx�����8[��w�|�T'p���^�J�I��3�������_�wӻ�6񛽾-��l(f�h�Z�7�f��܆�(ݨ���ٽ���r03���^�Cj��~=������)�¾RJξ�;Ӿ�GѾ��Ⱦۏ���,��;���z�s�O���'��   �   �[�N۽4���X��?�Z����������r��8�Ԃ>��̓��ϭ���ڽ8����XL+��W9�-eB�. F���D��>�B�4�"t(�E>�i&������ٽ�1���,������
��$U������|���Mٽ,�
��1�V�`������E��p=þ��ܾ7�s���/
�{g �T=�����ʾ�ȯ��ݓ���q�̍?��   �   �$�TN�Z��u�Z��5�ܬ���� A»�{ ��bi���ȼ�0�?l[������6��Wֽv���H�,|�n�����a������(u�6���N8�mhٽ��Ž�N�����fޠ�����n����ֽ�	�:�(�	GW�l���6U���ɾ�q�ZS�t��k�l��'����I��#�3ξ�����f�Y��   �   �7�L���^����b�ht���^��$���F;@;r; Z9H��L���L����,�l�e���D���W���Խ��住e�t�������T���Q��W�I����ݽ��н�|Ľ	_��׿��+?���սL���>(�ȟE��{��᝾�¾X��M+�S����'���0��	4��11�c{(����yj	����(�þN��_t��   �   �)H�֡�����/m�B����4�p�	;d�<��I<��3<���;@*x���&��n���I�2�4��<d�����[���γ��Г��6$нQ#ܽa9彫���������>�Wݽ ~ԽGjν�{ν2�ؽ=�����cm0���^�=Z��^���`�ھ�Z�Q���,�q6<��XF���I�V�F�=�<�-��n��c��zپL���"p���   �   hV�o����ʽ`zw��e�������;��e<�Y�<jw�<p�~<�&<0G6;�&ƻ���p�ؼY���*E�J q�Y卽Z��������ǽ�׽��
����x�콢��w�F޽
�߽�D콊�����XH@��r��ș��(�������$U&���;��vL�}fW��9[���W�{�L�ޣ;�N(&���3�꾲b��Z���   �   �6_����e4ҽ��~��@�H	�;Hz�<*��<��<4�<ԑ�<di*< �*;P�лک��H�ټ�#��FF�t�>�~g��x���O�Ͻ{M߽`�꽌��+򽿂ｔ#뽰O��4뽊�����@$��cJ��:������"˾�;��*���.��#E��V��Sb�{Lf�8\b�(�V���D�Z.�+�-���ľЖ��   �   �cb������Խ�π�����(��P�;�<ͺ<̴�<
�<rA�<��S< ��;�\S��"R�zH����
��[8��g�,A��J���?��lMͽ�:޽.�꽊	�%���.�2Y���K���Vq�o'���M��Ɂ��}��@�ξxv�������1��qH�zwZ��f�Xj��f��hZ�I2H��.1�}i����XǾ<���   �   �5_����[3ҽC�~���4���;"{�<�<t��<�4�<4��<j*<p�*; �л.���p�ټ#�*FF�Gt����f������}�Ͻ�L߽[��v��*򽘁�o"뽋N��3�R��� �M?$�	cJ��9�⾡�"˾�:��m)���.��"E�)�V��Rb��Kf�E[b�C�V��D�ZY.���&���ľaϖ��   �   �V�����ʽuww��a��������;��e<�Z�<@x�<��~<\	&<�L6;$ƻ��L�ؼ����)E��p��䍽c���g��O�ǽ�׽���꽰�X��t��K	�޽��߽�B�F��c���F@��r��Ǚ�5'��������S&���;��tL��dW��7[�0�W�ƠL�M�;��&&�T�<�� a���X���   �   %'H����+m�f�����4���	;̅<��I<`�3<���; x�l�&��m���H�m�4��;d�������������v����"нf!ܽ*7�.��G������;�Rݽ�zԽ5gν�xν��ؽ�������j0���^�bX�������ھY�[�P�,�4<�4VF��I�טF�ߨ<��-��l��a��wپ"���pn���   �   �7����4[��̗b�\m����^� �#�`�F;�Jr; 9H��"�����$�,���e����������� �ԽL���c���9���9R���N������g�ݽ<�нLyĽ\[�����8;����սi���V%�6�E�M{��ޝ���¾W���(����$�'���0��4��.1��x(�h��0h	������þlK���Zt��   �   ��$�GI����Z��1�B������5»�w �\_i�T�ȼ0��k[�5����6���Vֽ�������{�Sm����`�������s������4�dٽ�Ž�J�����Dڠ�=���������ֽ��S�(�6BW�q����Q��Uɾ�l꾊P�q�Vh��h�l$����F����	ξ���Y��   �   AX��H۽@0��^�X��;������������p��07��>�n̓�=ϭ�M�ڽ����L+�:W9��dB�}F��D��>� �4��r(��<��$�´���ٽ�-��i(��r��������P������v��Gٽ,�
��1�P�`������A��k8þ��ܾ������Fd �@7��Y���ʾmį�@ړ��q�_�?��   �   &��ʽ�d���P^�4L$���t7꼯� ��o#���\��g��<<Ž���������7��R��>h�Zmx�r����Z����|�U&p���^��I�3�a��ח� \Ὂϻ�6훽�)�� f���Z���f�p׆��֨���ٽξ��*3���^�'f���8��g���d�¾EDξ�5Ӿ�AѾ�Ⱦ����F(��7��p�z��O�_�'��   �   ���ܿ�8ٖ�?�m��A�G*�2G*�dNC�+v��k��w�ӽ���^+��5P���t�.��ȷ��yH��覾�F��6���"���JU����s�US���2��O�Q��Dݿ�.ٖ�'�m��	A��*��C*�)JC��%v�Gh��t�ӽ����[+�%2P��t�� ��O����E��u妾)D��К������lS����s��RS��2��N��   �   '[�hϻ��훽�*��z"f���Z�X�f��ن��٨�Z�ٽ���U-3��^�h��;������+�¾1Gξ�8Ӿ�DѾ¹Ⱦ���l*���8��C�z�5�O���'�'��ʽ4e��P^��J$����1�� �k#���\�Td���7Žj������3�7�R�b:h��hx�<����X����|��"p���^�r�I�-
3�������   �   ��ٽ�-��)������*���PR�����Yy���Iٽ��
�Z�1��`������C���:þ��ܾ�$������e �4:��	��Z�ʾ`Ư��ۓ�O�q��?�kY�]J۽�0����X�	;�h�� 
��f����h��M2�|>��Ƀ��ʭ�8�ڽ����H+��S9�aB�F���D�:�>���4��p(�:;��#������   �   �dٽ��Ž�K������۠�������ֽ���(�cDW�͘��BS��Yɾo��Q��r��i�qj��%����DH�� �ξ �P��޾Y���$��J�����Z��1������"»�j �POi�|�ȼ"*��d[�!����1���Qֽa�����x��j�����^���&���r�~���4��   �   ��ݽ��нJzĽ�\��~����<��n�ս�����&�ŝE�B{����.�¾1��*������'�$�0�4�01��y(����Si	�����þ�L���\t��7�؛�6\����b��m��|�^� �#��G;�qr; .9ȶ��뉼F��Ն,���e��������V����ԽU��W`�`������HP���M��t����   �   b<�ݽ�{ԽFhν�yνA�ؽ.������k0�.�^�-Y�������ھ�Y�B�X�,�25<�jWF�Z�I��F��<�-��m��b�Hyپ2���@o��O(H�������,m������4��	;Ċ<��I<T�3<��;@6w���&��d���C��4��5d�ܽ������򯰽���j н�ܽ�5�b���������   �   ������	��޽��߽gC�������JG@���r�ș��'�������YT&���;��uL��eW��8[��W���L��;��'&���F���a���Y��yV����k�ʽgxw��b�����p��;��e<�\�<�z�<��~< &<0u6;�ƻ�x��,�ؼײ��%E�Y�p��⍽ʇ��	��:�ǽ2׽S�������   �   �*����"��N�84뽿���Z��?$�OcJ�:����M"˾�:���)��.�E#E���V�Sb��Kf��[b���V���D��Y.������,ľ�ϖ�Y6_�8���3ҽ��~�g���0�;�{�<���<���<6�<:��<�n*<P�*;��л������ټ,!�TDF��t���1f��0����ϽRL߽G�꽈���   �   �?���՚�����_���<��9�轚���`A�_b������^޾�&�<�0���T�y0x��ʋ��1��(��Y袿|(��R(�������w�^�S��/�ޅ��־8���
c��U��sĽ�`���μx���xl<�q<���< �r<&<�)f;����[V��2������v���>�QsZ��s�&���Č�Vf��kᗽ�0��ݢ���   �   姚�hE��V����%���?��"��*�0'>�L�|�<M����ھ�����-�rsQ��!t�Y���t���/����L��D���컕��n��%�s��P�t=,�	R	��PӾoʜ��_�5�*����+^���ͼ�1��n�;<�\<�1t< �M<8��; z9�"��ȍ��ټ����4�D�R���m�����������٘�P�����%���   �   ~@��r[���2䡽X�����ٽb�	�j�4�&p�x��D�Ͼ����V%�:GG�Xh�삿�������Ƿ��]+��������.h��F��+$�J����ɾ�ŕ�H�U�����#���V�̼H1һ��;,:<��<���;���������p���U&�m�N�$�r�䀈�є�X2�������x��ɶ��ީ��9���l���   �   _��z◽�_��G�������?�Ƚ�����&�_�\�Q���G���������g7���U�06q��j���c���،�҆��������q��AV�&i7�	��N򾊫���ꊾ�F����h���DL�zp̼�U� p�8�!7; ��9xp���Qy� %ڼ�� �'�U����Ǜ�	P��'d��e�Ƚcν��ϽI2ͽ��ǽ�`��zw��ڜ���   �   ����gɘ�kD���7��^𘽩1��d὾\��D����^!��٘پ�\�>F#�J�>���V��cj���v�zp{�aw��%k�=�W��~?��	$�����%پ#ߧ���z��64�_����נ�Q�A��vҼ8�M�H�ڻXa滠)O�ԝ��<1�O;Q�z���:ʬ���̽ �轾����
�.�2���%�^����0⽊eν\{���   �   tɵ����$�����10��xa�������9���(��l_�3G���3��<�T���.$��Z9�H8J�0U�.Y���U��SK���:��%�rK�\
��_������\�E��b�ݽ�Ē���8�⼺Ҕ����⡥��a��}�6�:ـ�|z��N�ؽR��;��)�d6��=���?�Ɍ<��m4��~(����.�	�+����ҽ�   �   �k˽�������\x���p�Zf��6ǟ���Ͻl�
��9��r�ਛ�����*�j������(�v2���5���2��K*�g��re�B��g�Ǿ�	����{��e>��D���ĽG��B�4������9Լp�強\��4U������fǽ�G �b�<��W��~m�(`}�%Ƃ�Aɂ���}��7o�'f[��'D��M+�bt�O����   �   �5꽈Ը�<��I�o��U��AZ�����A��ؽ۽�Z��VB���y������~�ܾ�p���O����U����RT
�W>��`���ľ� ������S�"�>�٢����y���7�����p�/���j����T�ٽ����d4��\�����t3��C����~�����Pծ��9��>�Q!���;z�<vV��@3��`��   �   JT	��^ѽ������o��B���3��JE�F�w�|����'�� ���@�N�q�/�����m�¾l6վ��~��<�UqھHiʾٸ��=��υ��\�o0��R	�]ѽɌ����o�3�B�n�3�UNE���w� ���,��#� A���q�ʲ������¾:վ��J���?��tھdlʾ����Z?���Ѕ��\�h0��   �   �"�C�죮�H�y�>�7������/��j����N�ٽ|��"a4�l\�����0��3���p{��w���3Ү��6������7z�AsV��>3�A_��3�ZӸ��;��ӥo���U��DZ�F���D����۽R]��YB���y�k�t���ܔܾ�t���Q����x����EV
��A��m�㾜�ľ���t��`�S��   �   {g>�F���Ľ�G����4����Z4ԼƟ开W�.U������aǽ�D �m^��<��W��ym��Z}��Â��Ƃ��}�a3o��b[��$D�[K+��r�����Fj˽S���򮌽^x�Ȫp�h���ɟ���Ͻt�
�i9���r� ���6���#-�6�����(��2��5���2��M*�G��g���ﾗ�Ǿ=��,�{��   �   �\�x����ݽJŒ���8�⼦Δ��ق�z����V����6�Հ�zu��v�ؽ�����)�Z6��=���?�.�<�Qj4�|(�Y��d�	�����ҽrȵ�B��D$��W ��d1��0c������<���(��o_��H���5������]0$��\9�r:J�P2U�`0Y���U��UK���:���%��L��쾭a��A���   �   K�z��74������ؠ���A��uҼ@�M��|ڻ8G滈O�����*��3Q� ���0Ŭ��̽�轲��� �
�~	�����#����*.⽫cν/z��X���Oɘ��D��W8����W3����2^��D�����"��ߚپ6^��G#���>���V��ej���v��r{�cw��'k���W�a�?�:$����3'پN৾�   �   �늾��F���������L��o̼�Q� ��8`H7;�J�9�P���>y��ڼ�� ���U��������K���_��R�Ƚ�_νH�Ͻs/ͽ��ǽ_��Dv��&������◽`�����������Ƚ����&��\�!R��(I���������h7�>�U��7q�wk���d���ٌ�����Ȥ�� �q��BV�2j7�����򾃬���   �   �ŕ���U����#��@�V�~̼0+һ��;x@<�<���;�@�����2렼���P&��N��~r�4~��tΔ�0������6w��`���Ш��������h@��������䡽5�����ٽ 
�_�4�hp�J��V�Ͼc��ZW%�0HG�Yh��삿-���b��k����+�����������.h�ֵF�4,$����Q�ɾ�   �   �ʜ�K�_�N�:����+^�Z�ͼx-���s�;�\<T6t<\�M<@��; �{9��Xč���ټ9���4���R��m�����Q����ؘ�������%��꧚��E������@&��8@����E+��'>��|��M��J�ھ4��Z�-�tQ�1"t�����ͼ������ M������5����n����s�:�P��=,�<R	�6QӾ�   �   �7��[
c��U��sĽ��`��μ����Hm<��q<$��<��r<�&<�+f; ����ZV�h2������m���>�ZsZ��s�8��
Ō�cf��}ᗽ�0��𢚽�?���՚�����_�� =��p�轾��aA�b��	 ���^޾�&�X�0���T��0x��ʋ��1��%(��[袿|(��N(��񧋿�w�H�S��/�ʅ��־�   �   �ɜ�Q�_���9���_*^�^�ͼ�'���w�;,�\<d7t<<�M<(��; |9���Í���ټ����4�:�R�}�m�����0��֌��Vؘ�=�����$��&����D��Ι��\%��@?���彗*��&>��|�M��Z�ھ�����-�sQ�+!t����/���㔝�xL��򙝿����en����s�]�P� =,��Q	�SPӾ�   �   �ĕ��U�ķ��!����V��̼� һ�'�;8C<��<ț�;`5������꠼l��AP&���N�~r��}���͔�^/��ٯ��Pv��U�������>�������>��혽&���㡽R�����ٽ��	���4�Np������Ͼ?���U%��FG�(Wh��낿����%��)����*��w�������-h�0�F��*$������ɾ�   �   �銾V�F����N����{L�Dj̼HJ� l�8�V7;���9 M���<y��ڼ� �w�U�H�����TK��[_����Ƚ�^ν<�Ͻ6.ͽ6�ǽj]��~t��<�����|����]������������Ƚލ���&��\�:P���F���������f7���U��4q��i��c���׌�����(����q�,@V��g7������*����   �   �z��44�2���^ՠ� �A�"oҼ }M�pڻ8>�\O�䑸�<*�3Q�ƒ���Ĭ���̽���4������
���,���"�M���7,⽒aν�w�������Ƙ�B��v5��f�/��,�t[�[
D���� ��#�پ�[��D#�Ì>�6�V��aj���v�in{�_w��#k�d�W�6}?��$�|���#پ�ݧ��   �   R�\�����ݽ�����8��⼪ɔ�xւ����U����6��Ԁ�6u��2�ؽ���k���)�6���=���?���<��i4�>{(�l��X�	�<���ҽ�ŵ�t|��T!��,���-��%_��4����6���(��j_��E���1��������,$��X9�66J��-U��+Y�j�U�iQK���:�=�%��I����]��: ���   �   �b>��B��Ľ�C��ʽ4�����N/ԼJ��UV�E-U�b���Eaǽ�D �M^��<��W��ym��Z}�bÂ��Ƃ���}��2o��a[��#D�MJ+�rq�S����g˽x���꫌��Wx���p��c��zğ���Ͻ��
�_9�s�r�����8���&'꾼�������(�>2�X�5�o�2��I*�d���c��ﾷ�ǾS���{��   �   9"������,�y�,�7�g��C�2�/�b~j�������ٽV��a4�N\�����0�����S{��P���Ү��6��R����6z�@rV�{=3�
^�51꽖и��8����o���U�y<Z�t��>���۽xX��SB�0�y��훾Ί��K�ܾ]m���M�|��-�����DR
��:�����	�ľ-��������S��   �   :P	��Xѽ����2�o�E�B���3�HHE���w�����&'�� �c�@�1�q�"�����`�¾Z6վ��`���;� qھiʾ�����<���΅��\�T0��Q	�|Zѽ�����o���B���3�EE�5�w�榥�#�,�!�@�*�q�����.�¾�2վT�ᾞ��=8侢mھ�eʾ����\:���̅��\�"0��   �   �.�"ϸ�8����o���U��>Z����@A��c�۽�Z��VB���y��~���r�ܾ�p���O����J����=T
� >���㾺�ľ^ ��t��!�S�"�
�q���j�y��7�����C�/�yj�"�o�ٽ���]4�&\������-��&���6x��&����ή��3���윾V��3z�oV�;3�B\��   �   �e˽~�������Xx�#�p�$e��`Ɵ�I�Ͻ;�
��9�c�r�Ԩ�������)�f��ݔ���(�p2���5���2��K*�T��Xe����Ǿ2	���{��d>��C���Ľ�D��'�4����8+ԼΕ��Q�N'U������\ǽ�A ��Z��<�ZW��tm��U}�����Ă�ڿ}�n.o��][�� D��G+��o������   �   �ĵ��{��L!������.���`�����9��g(��l_�'G���3��4�P���.$��Z9�F8J�0U�.Y���U��SK���:���%�ZK�"
쾲_�����o�\������ݽ����8�*��Ɣ��т�����HK����6��Ѐ��p����ؽ�����
)�!6���=���?���<�Vf4�[x(���p�	�a���ҽ�   �   %����Ƙ�NB��6��J�0���ὖ\��D����V!��Әپ�\�<F#�G�>���V��cj���v�xp{�aw��%k�4�W��~?��	$����l%پ�ާ� �z�64�����֠��A�oҼ�yM�xaڻ�(�|O�H���A$��+Q�����"���x�̽��@���
���
�B����� �ď��v)⽌_ν�v���   �   ���l���^��,���¹����ȽD����&�H�\�Q���G��������g7���U�/6q��j���c���،�҆��������q��AV�i7����+�b����ꊾ��F����\����|L��j̼@H� ��8pu7;���9@1���+y��ڼ� ���U���������"G��$[����Ƚ[νǫϽ<+ͽ�ǽ�[��!s��Z����   �   �>��혽^����㡽޲��r�ٽH�	�T�4�p�s��B�Ͼ����V%�9GG�Xh� 삿�������ȷ��]+��������.h��F��+$�@����ɾkŕ��U�t���"����V�f̼ һ -�;�G<��<8��;�ހ�t���⠼���pK&�s�N��xr�"{��[˔��,������jt��ʲ��v���b���"���   �   ����D��䙝��%��w?�� ��*�%'>�G�|�:M����ھ�����-�psQ��!t�Y���t���0����L��E���컕��n��#�s�ނP�p=,�R	��PӾaʜ��_������$+^�"�ͼ�(��0y�;�\< :t<��M<���; �}9��п����ټz��4���R���m�f�����苓��ט���x�$���   �   O�N��/T� Pj�����?ε�����)+���n�V���^�O��lA?�Fn�Dk���Ȧ�s���˿S*ֿ?�ٿ/*ֿ#�˿6A���e���Ў�Εl��<�;��r`ؾK����BU�\���m��@}9�� �� Ee�  �;���;p�;@,��	�����pJڼ�4�ê3�w�O�The��Ft�||�L}~�H!{���s�A-i��]�X�S��   �   �S��WV�;j��h��J��^��3c(�'�j�iA��_hܾ���<�[`j��������v��%ȿ��ҿxZֿS�ҿ}ȿLV��$̣������h��9�0K��Ծ旘��R��	��8���8�>s�� ����X;���; M	;6��GM��a��%��H�*���M�2 k�1e���w���͊�.�������I��0�v�~Eh�-[��   �   �`b��i]�D�i��އ��,�����3U ��e_��^��ʧѾ&�
���2��_��X���T���ɯ�����ȿ�h̿}ɿQ>���֯�d9��	����]��G1�J���$˾4���Q�H����C񡽱Q4�����0�컀;��@�ź�	ѻ 7p��=μ+
���G�cv�^-���9���]���Z���X��lέ�����h�����p��J�r��   �   ?}�<,k�q�k����񛡽}ֽ����M�������������$��`M�2�w��'��]4���p�������ռ�]ʹ�����}���S��w�\�L���#�	U��$ѻ��↾�O:�ǜ������s�/������G�����uN�敪������?�Ť~�vɞ�������Խ��MI�v���j��"��Aܽ��ɽ����X��b��   �   0���6���Ir��}��,���V������07�~�|�ذ�������+�6���\�Q���������������z�B���)���e������a]��67��a�z��Mx���r�`/(�r߽ë�� �,�2׼P࠼�������߲*��Jp�.F����ʽ������^��	r)���/���0�L,���"�Y�:��߯���˽�A���   �   ����Q7��B[��l�w�)���dU��֡�-����Y��Γ���þ�n��_��<O>�:^��ez��i�����L������ ����{�۝_��?����*���EVľ֒�NT�C%�ԏǽ
낽��-�TX�֒��ō�\M��T���o������K���75�I5O�\zd�UHs��qz��y���p�2�a�6M�z|5��]�����5ٽ�   �   ��ڽD����H�x�a�{�V���nu��Z��x+5��v����9Ҿ�L�/��C_9�f>Q�l9d��p��u��Tq��e�e S���;��� ��_�O�վ�쥾%Oy��`5������i��t��>5�Lr �k92��`g��=����ֽ�/�e�2��Z������@���y������V��	Ԭ�Mإ��%��劾O�r��oN�Q�*�b�	��   �   J����Ͻ��������
�l���~�����s	ԽPn�n�E��6���A���Ӿ����Ț�d)��8�պB�&�F���C��=:��\+��_����Z�پ�P��������N����Uڽ����h�:�D� J�wlw�������ۈ��
E�,�w�hV��4S���Ǿs�ھ�=羁Z쾋��l;߾oξ�ϸ�tO��dᆾFo\��9/��   �   ��(�{���T鹽�H��v1f�m+]�Q,~����>����3�K����������ǾP�����_��w�R���w��Q�����v�lϾI���Y����\��(������繽>H���1f��-]�e0~� ����������K�♃�t¤��Ǿ\��2�5b�6z���Zz�[T�����z��oϾ�K���[����\��   �   '�N�q��Wڽ�����h���D���I�5gw�Թ���⽟���E�,�w�pS���O��'�ǾH�ھx9�V�A��h7߾pkξO̸��L��8߆��k\�J7/����P�Ͻ����6����l�Z�~������Խ�p���E��8��vD��T�Ӿ�������)�̖8���B�
�F�ʜC�L@:�0_+��a����>�پ4S��a����   �   �Qy�Sb5�����j���t�=5��o �52��Zg��9��I�ֽh,�J�2��Z�.���s=���v��b��QS���Ь�ե��"��|⊾��r�llN���*�W�	���ڽ��� �:�x���{������w��.��.5�-	v�( ��T<Ҿ�N�G���a9�AQ�S<d�	�p��u��Wq��e��"S���;��� �a���վ��   �   Uג��OT�g&��ǽt낽��-�FV�؋������M�4P��Tj��s���w��]35�i0O�ud��Bs�`lz���y���p���a�2M�y5�>[�����2ٽ⭱�6���Z���w����W��n����b�Y��Г�*�þ�q��#��XQ>��^�7hz�ek�������M��
�����2�{��_��?�������Xľ�   �   ~y����r�o0(�Bs߽>�����,�/׼۠�����h��(�*�ZBp�5A����ʽ:����n���m)���/���0��,�0�"�`����ӫ콬�˽{?������.5��2Ir��}��-���X��:���27���|�u���ޕ�?����6���\�q���␿���%�����qC��+���f������c]��77��b� ���   �   һ�.ㆾ^P:�Ý��d���O�/�j���G� ���fN�*�������?�_�~��Ğ���"�ԽZ�罊C�hp��je��^���<ܽL�ɽᛵ�.����=}�K+k�v�k�"��朡��~ֽ����M����W���������$�bM��w��(��k5���q������ּ�{˹�����~���T��*�w���L���#�dV���   �   J%˾������H����񡽎Q4�t������@����Cź��лH'p�`4μ��x�G���u��)���5��&Z��W���U��l˭�j}���f��I����n��d�r��_b�Ti]�|�i�2߇��-��*��V �%g_��_���Ѿ��
���2��_�kY��PU���ʯ������ȿ�i̿Jɿ?��nׯ��9���	����]�KH1�����   �   I�Ծ����R�$�	��8���8�2r��(��� �X;���;`h	;�%��l=M�R\�� ����*�`�M���j�dc��v��(̊�����ɞ���H����v�CDh�G,[���S�kWV�vj��h���J��*��c(���j��A��iܾ�p<� aj���9��jw���ȿE�ҿ�Zֿ��ҿd}ȿ�V��j̣�X���)�h�b�9�aK��   �   G`ؾ(����BU�/���m���|9����� @e�0"�;���;X�;�,��	�&��� Jڼ[4���3�f�O�@he��Ft�||�`}~�b!{���s�a-i�7�]���S�{�N��/T�VPj�Ĵ��|ε�`����)+�;�n�������p���A?�@Fn�Xk���Ȧ�%s����˿Y*ֿD�ٿ.*ֿ�˿+A���e���Ў���l���<� ���   �   c�Ծj����R��	��7��S
8�|p�����@�X;���;�k	;�$���<M�.\�������*�7�M�n�j�Dc���u���ˊ�|���x���dH����v�hCh�T+[���S�AVV�2j�:h���I������b(��j�9A��hܾp��<�`j�{������v���~ȿk�ҿZֿ��ҿ�|ȿ�U���ˣ�Ǒ��5�h���9��J��   �   �#˾g����H�����#O4������컀欺�4ź��л,&p��3μ��B�G���u��)���5���Y���V�� U���ʭ��|���e�������m����r��]b�g]���i��݇��+���罕T �+e_�-^���Ѿ��
���2��_�MX��T��/ɯ�	��M�ȿ�g̿�ɿ�=��֯��8��}����]��F1�����   �   �ϻ�tᆾ�M:�H���������/������G�����cN�&������4�?��~��Ğ�����Խ��3C��o���d�����<ܽ`�ɽϚ������E:}�)(k��k���j���g{ֽ��ƫM��������������$�v_M�Ȓw��&��l3���o��ߙ���Լ�>ɹ�����|���R��!�w���L�}�#�:S���   �   �v��f�r�y-(�o߽P�����,��)׼Lנ�R�ʕ꼃�*��Ap�A����ʽ�����S���m)���/���0�=,���"���+�����D�˽�=������P3���Dr��}��*���T�����P/7�~�|�������������6�ӳ\�N����ߐ�m���r�����@��x(���d������_]��47�+`�\���   �   FԒ�TKT�*#�}�ǽ:肽|�-�<S�ć��\���M��O��j��<���]��D35�R0O��td��Bs�,lz�`�y���p�4�a��1M��x5��Z�А�.1ٽ
����3��rX��z�w�̫���R����q����Y�R͓���þkl��͕�WM>�^�cz��h�������J�� �����	�{�w�_���?�˷�O����Sľ�   �   �Ky��]5�r���4f���t��85�}l ��22�QYg�,9���ֽG,�.�2��Z�$���i=���v��Q��9S��sЬ��ԥ��"��:⊾]�r��kN���*�~�	��ڽ`�����x�2�{�����er�����#)5��v�����6Ҿ_K�B��]9��;Q��6d��p�}u��Qq�7�e��S�V;��� ��]�o�վo꥾�   �   C�N��QQڽk��S�h�$�D���I�.ew�+���)�v��cE��w�eS���O���Ǿ>�ھh9�V�'��A7߾?kξ̸�|L���ކ�(k\�z6/����G�Ͻ2���~���w�l���~�x����Խl�y�E��4��_?���Ӿ�������
)�f�8��B�F�F��C��::�:Z+��]���� �پ5N��~����   �   G�(�t���x㹽�D���+f�X']��)~�����������K�t���~����ǾI�����_��w�L���w��Q�����v�qlϾ�H���Y����\���(�ĸ���幽�E���+f��%]�I&~�������S����K�L���ʼ��M|Ǿv����^]�u����Au��O�����r�iϾF��~W����\��   �   �����Ͻ����ҹ��Իl��~�V����Խn�B�E��6���A���Ӿ����Ś�d)�
�8�ҺB�"�F��C��=:��\+��_�����پ�P��^����N� ��Sڽ���2�h�7�D��I��`w�ﵥ��	⽍���E�w�w��P��zL��n�Ǿ6�ھ%5羮Q�އ�.3߾�gξ�ȸ��I���܆��g\��3/��   �   �ڽN��r��x� �{�թ��lt����A+5��v����u9Ҿ�L�-��A_9�e>Q�l9d��p�~u��Tq��e�[ S���;��� �w_��վw쥾�Ny��_5�=����g��Zt��85��j �\/2��Sg�z5���ֽ/)�a�2�]�Z�z���h:��Js������O���̬��ѥ�����ߊ���r�hN���*�H�	��   �   ����x2���W��K�w�\���*T��
�������Y��Γ���þ�n��\��<O>�7^��ez��i�����L������ ����{�Н_� �?�{�����Vľ�Ւ�MT��$�D�ǽ邽��-��Q�B���!���	M��K�� e��.������/5��+O��od�V=s��fz��y���p���a�~-M�u5��W�����-ٽ�   �   B���A2��	Dr��}�<+���U������07�]�|�Ͱ�������)�6���\�Q���������������{�B���)���e������a]�x67�qa�T��!x��y�r��.(��p߽G���8�,�(׼^Ӡ��쪼��꼌�*�E:p�b<��C�ʽ�	��t������i)�w�/�ŋ0�t,�W�"������J����˽p;���   �   �7}��&k�l�k�>��򚡽]|ֽ���٬M�|�����������$��`M�3�w��'��]4���p�������ռ�_ʹ�����}���S����w�T�L���#��T��ѻ�^↾%O:����ߖ����/�<����G����VN���������?�H�~�������Խx�罂=�dj���_������7ܽ��ɽʗ��������   �   \b�6f]���i��݇�A,�����U ��e_��^��ŧѾ%�
���2��_��X���T���ɯ�����ȿ�h̿~ɿR>���֯�d9��	����]��G1�B���$˾����H�������O4� ���P�컠��� �ĺP�лXp�p+μ�����G�,�u�D&��.2��KV��2S���Q���ǭ�z���c������ml��_�r��   �   ʃS��UV��j�<h���I��0��!c(��j�fA��^hܾ���<�Z`j��������v��%ȿ��ҿyZֿU�ҿ}ȿMV��#̣������h��9�,K���Ծۗ���R��	�h8���
8��p��������X;�ȣ;0	;����4M��W��F����*���M��j��a��.t��Nʊ��������>G����v��Ah�3*[��   �   D��a	)���K�&����ý����rP������gӾ�:���A�1cy����U��!�׿]��a��
��l�<
��T����)׿K;������R�v���>���� ̾�A��$�;����D��0L��)���ػ`�x���ԻgV�J���?��-0�iX�΢z��H���f��(n��Q����:���l��Y�n�9kT�4�;��I(��   �   (���-��LM��	���)��
���$M������Ͼ���p_>�'Qu�M������SԿV,�{O�H���6
�����L�����ӿ)b��"���|
s���;�b����Ⱦ���� 9�w�L슽�T������f	�(�лD@"�;����߼z��/UL���w�r
��춛�]�������fT��
ᐽ�₽°g�1�J���3��   �   CA��=��S��S��k���:���C��z��!�žb���5��~i�9J������pʿ�������T��v������g0��Gʿ��&���ټg���2�.B�7���g҄��"1��὚������"����c��)i�X��l���A[0��`i��:���v���S��a8ѽ�#ڽ��۽�Tֽ�ʽ�(���l��&^���	z���W��   �   k�l�N7X�۶^�����<�~���J�4�>����1�����C�&��W�j������j�ѿ������D���Z俏Cҿ�0��� ������ V��3%��������v�~�$��Խ�g����!�d�ټBվ����Ԥ�W�W�Ǒ���ߵ���۽�=���F��<�pI��.�� �(���� ��*���Ľ)䥽�؊��   �   �N��z��)�r�d@��������<"��Eg��_��5�޾�k�H�?���n��ӏ��5���ݻ�C'̿��ֿ�pڿ�׿	�̿����&ϧ�c7��04o��[?����*Bܾ�Ş��h]��`���ý&�~��P/����1��VA�L����S������
�T�$�*�<�ߪO�A�\���b��_a�_�X���I��i6����6�$S�׸��   �   �Ľ�ݞ�V8�����Û���˽���_2H�����쿾\����%�s&N��x�Ƹ��Ң����7Y��Ʊ���˺�lⱿ����柑��z��7O�F�%�0����*��;����A��~�X+��Fvz�r�E�"�@���d��g��eTɽ���N.'��,L��jp�������r���a������ݲ�� ��H�^��=<�ю������   �   �^ �� ǽ�<���c���������~�.(��/j����,վ#�	�� ,�H�O�)@r�)}�����󊜿�m��b������叉��t���Q�>�-��H%׾�$���1j�v�%�de������|���f�	���4ң�P۽Q���=�`<n�����\���"���>Ҿ�E޾�@�f"־�ž�����ᘾ�/����P��C%��   �   7%&������j��j����]��QC����ɽgM	�-�=��:��H�� ޾9�
���'���C��&]�y.q��9~�n����,���r��y_�N�F��c*�9A��p�ѳ��6��&�A�(-�w�ȽW�����������4���������I������m����ž��羹�:?�^E��[�z8���s��";���
H���Y��   �   �S�/��s�����ȑ�V������6ڽ�{���I����&��T�ؾ��]4��-�U=��oG��XK��`H�X�>��/���r��޾�:������S�$���置���ȑ�v�����:ڽz~�P�I���&)��$�ؾ�� 7��"-��
=�sG��[K��cH�w�>���/�<�� ���޾@=��,����   �   �7��t�A��.� �Ƚ����$�������1��N�ར����I���Vj���ž2��6��<��B��X��5�.������;����E��UY��"&�k����h�������]���D��nʽ|O	�'�=��<���﫾�޾\�
�M�'���C�F*]�2q�>=~�L����0�=�r��|_��F��e*�'C��s�����   �   r&��d4j��%�,g罊����|���f�w���iΣ� ۽�����=�7n�r����������$:ҾA޾R㾅;�־)�ž9����ޘ��-��4�P��@%��\ �Eǽ;��"c������������0(��2j�.���/վ��	�C,���O�ECr��~����ጜ��o��H������������t��Q�F�-����'׾�   �   i,��R<��g�A���,���uz�C�E�~@���d��c���Nɽ���(*'��'L�:ep�ڊ������ܛ��w]��~����홾ү��S����^�,:<���l�����Ľ�۞�J7��q���Û���˽8���4H�l��￾G����%��(N���x�R����Ӣ�\��[�������ͺ�.䱿#���Q���Pz��9O�ݷ%������   �   �Cܾ�ƞ�#j]��a�p�ý�~�.O/�t�����PA�(���zN�����@�
��$�q}<�ʥO���\���b�jZa�m�X��I��e6�}��<3��N⽲Ӹ�dL������r��@���	����b>"��Gg�a��L�޾m��?���n�#Տ��6��߻��(̿��ֿorڿ�׿��̿&���mЧ�}8��6o�[]?�·��   �   � ������v�1�$��Խ�g����!���ټ�ξ�>��Ğ��W�>����ڵ�ļ۽�6��GC�9��E��*�r����� �&�ӕĽ᥽r֊�;�l�f5X�3�^�>���,���/�����4�1���'3�����v�&�4	W�U2��������ѿ���k��{����K\��Dҿ�1�����Q���1V��4%��   �   �B�΋���҄�:#1�w�὞�����8����c�$i�f ������yU0�Zi��6��Nr��LO���3ѽ;ڽH�۽�Pֽ�ʽ%���i���[���z���W�PA��=��S�"T��>������C�F{��*�ž���5��i��J�������qʿ� ����x������������@1㿝Hʿ���������g�`�2��   �   ���	�Ⱦ���!9�w�4슽TT�䔑��a	���л�7"�6����߼��^QL���w�:��������`����죽~R��\ߐ�xႽm�g�]�J���3�D(�"�-��LM�
��Y*��~���%M������Ͼ2��`>��Qu�����{��wTԿ�,��O����87
�4���L�C��i�ӿrb��]����
s�ʼ;��   �   ��� ̾�A����;�A�����K��(��ػ0�x�h�ԻfV�������-0��hX���z��H��yf��"n��V����:���l��r�n�ZkT�a�;�J(�t���	)��K�\���W�ý���rP�%���,hӾ�:�܏A�^cy����o��8�׿p��a�
��l�:
��T����p)׿7;������,�v���>��   �   ���0�ȾX��7 9��u�n늽JS�p���`	��л 7"��5��f�߼���HQL�o�w�,���������F����죽VR��&ߐ�=Ⴝ߭g���J���3�s(�.�-��KM�J	��`)������$M�{�����Ͼ���2_>��Pu��������SԿ�+�@O����6
����zL�S���ӿ�a�������	s��;��   �   �A�1����ф��!1�I����������Dc��i��������9U0��Yi��6��8r��8O���3ѽڽ�۽gPֽ��ʽ�$��i��$[���z�Z�W��A��	=��S��R��h������P�C�z��z�ž����5��}i��I��2���oʿ������n�����������v/�GʿM��}�����g���2��   �   �������v���$�~Խ�e��!�@�ټ̾����;����W�����ڵ���۽�6��9C�9��E��*�H�̺��� �o%� �ĽCॽ�Պ�$�l��2X��^�H����񰽳���/�4�����0�����V�&�~W��텿8������9�ѿ��㿎�ￓ����ￕY�EBҿ�/������������U��2%��   �   @ܾĞ�Zf]��^���ý�~��K/�>����OA�Մ��GN�����0�
��$�g}<���O���\���b�HZa�=�X���I�ve6�#���2��M⽘Ҹ�K��~��&�r�->������};"��Cg�E^����޾�j�Β?���n��ҏ�E4��xܻ��%̿Q�ֿ�nڿ#׿c�̿'����ͧ�(6��2o�2Z?�M���   �   m(��l9��D�A��|�(��jpz���E��{@��d�8c���Nɽf��*'��'L�,ep�Ԋ������ӛ��j]��m����홾����)��U�^��9<�Y��6���}�Ľ�ٞ�B5��� �������˽��G0H�j���꿾ڷ��R%�k$N�~�x�[����Т����_W��寽�ʺ��౿ؽ��_���7z�J5O�p�%�J����   �   r"���.j���%�Fa�r���|��f�:����ͣ��۽�����=�7n�k����������:ҾA޾H�t;��־	�ž���jޘ�\-����P�R@%��[ ��ǽ9���`�����񳽑z�l,(��,j���*վ|�	���+�˯O�@=r��{��K�������k��y��
��/����t���Q���-�G�`"׾�   �   �3��ޝA��*�L�Ƚ����n������`0�����g����I���Lj���ž.��4�<��B��X��5�$�������;���|E���Y�"&�̽���f�����|Z��3@��.�ɽ8K	�\�=�9���꫾f�ݾB�
�^�'�%�C��#]�+q��5~�����@)�D�r�wv_�[�F��`*�?�[m�����   �   1�S����潢��2ő��	�����5ڽx{�x�I����&��N�ؾ��\4��-�V=��oG��XK��`H�Q�>�ڔ/���^�P�޾P:��ݺ����S�j���V���ő�8	��U	���2ڽ0y�C�I�t��<#��̍ؾn���1�#-�>=�flG�=UK�X]H�(�>��/��$���޾c7�������   �   6&����ud��Ɉ��RZ��A��K�ɽ�L	��=��:��9�� ޾6�
���'���C��&]�x.q��9~�n����,���r��y_�B�F�vc*�$A��p⾙����5����A�Y,�b�Ƚ���� ��s����-����ར���I��|��Ng��m�ž���
��9��?��U��2�r�}��C�
;y��C���Y��   �   �Y �qǽ7���_��)����|�@.(�h/j�����,վ�	�� ,�G�O�(@r�*}�����󊜿�m��b������㏉���t�|�Q�/�-��%׾x$��j1j���%��c罓��%�|��f�!��^ʣ�	۽�����=�2n�v���=������5Ҿ�<޾�
��6ྡྷ־�ž����_ۘ��*����P�==%��   �   ��Ľ�מ��3��Y ������)�˽8��2H�����쿾S����%�p&N��x�Ƹ��Ң����9Y��Ǳ���˺�kⱿ����㟑��z��7O�8�%����}*���:��D�A��}�k)���pz�?�E�xx@���d��_���IɽE��7&'�$#L��_p�ȇ��=���N����Y��㵠�D꙾����h����^��5<�;��j����   �   ~H������/�r��=������低<"��Eg�t_��+�޾�k�F�?��n��ӏ��5���ݻ�D'̿ �ֿ�pڿ�׿�̿����$ϧ�`7��*4o��[?����
Bܾ�Ş�Fh]�*`�+�ý �~�K/���>�JA�"����I����ཱ�
���$��x<�ɠO���\�6�b�Ua�A�X�;�I�^a6�����/�I� ϸ��   �   c�l�u0X�ױ^�(����񰽭����4�*����1�����B�&��W�i������l�ѿ�������E���Z俏Cҿ�0��� ��������U��3%�������Sv��$��Խf����!�d�ټ�ƾ���������W������յ���۽�0���?�f5��A�'�������� �� ���Ľ�ܥ��Ҋ��   �   ^A�A=��S��R���������ݖC�{z���ž`���5��~i�9J������pʿ�������T��v������h0��Gʿ��%���ּg���2�&B�#���N҄��"1�Z�Ὓ�����蛫��c�i����������O0��Si�,3��6n���J��/ѽxڽ��۽Lֽ��ʽ!���e���X��} z��W��   �   .(�D�-�#KM�*	��b)������$M������Ͼ���p_>�'Qu�M������SԿU,�{O�H���6
�����L�����ӿ(b��!���z
s���;�^����Ⱦ���� 9��v��늽�S�����]	��л 1"��1��r�߼���ML���w���`���� ������ꣽ_P��`ݐ��߂�;�g���J�"�3��   �   �Y�H�"���P�9A����⽍u+���������)7�:t�=����¿#��J��.��t$��.-��>0��,-�D_$����I���Z���r��Vq�v4���&��
�q�L���㿽~�`����p���L>�ƶ��2Iټ%�C)I�,�z�Oۓ�w�������c���u��������<��������va��=��!��   �   φ!���)�j"T�����/$�)���{�X���Q��&4��<p�
s���m���l�����6�!��T*� W-�|[*���!�ؚ��?��俙'��Q���Tm��41����O����m�ƿ��;��{a�(��,������$'��f����1��Qg�P~��r���k��K/ɽ�Cн��ϽA�ȽS���I���>���,z�{Q�:A1��   �   ��C�z@���^�Bz���kٽ�"��Bp��쮾����g+�c�d�%��7u��1mڿ����f����~'"�:%��C"��:����̢��$�ٿN������Nb�%�(�0>�!:����c����יּ���d�������&B弨��.B����#ԡ��Yýj��@���N��y�	�:	����':��ʰܽ�e��񢽢$����`��   �   �J�z�f�SPr��ɕ���Ͻ�m��z^�\����侕��X�R�����ai��c�ɿ1�鿾�G�n��D�b��З��L�	�u�ɿ������? Q����T��o���Q�S���
��b��9l�~M-����Jc4�W�g��s��f�ý���;���)$�R�4�2�?�@�D��.C�� ;��-����	z����@��B-���   �   򥫽����lވ�p���|	Ž�
��GH��H���̾����;�b�q��|������
_ѿn��\������Z^��G����7���1ҿK��������q���:�Xv�0;ɾeÌ��?��D �����tz�C|U��a�n3���೽F�����*4��T���p���5���R܎�xC�����$�y��_��A���"�@"�iyս�   �   0�罟����(��\r��ٌ������p�/��sz�@F��e_���!���P�����v��������˿�ݿ���������޿`8Ϳ ߶�2d��ɷ��CjQ���!�����Ԯ��
v�Z�)���d���F��r��K7��˽���+���W��Ђ�[Q������ݽ���Ⱦ��̾DCʾJ��O��H���L����e�"�:����   �   G�R|ｗ���nC��ab���A߽��P`S�����#dʾ:��O.�
�Y����%�������f����@ĿQ�ǿ��Ŀq���Y鬿��M���s[��/�R��$˾����b�Q�����Hս<��ا�����,�ٽfQ���<�pgs��8��Q=��p�׾���8�_��υ�4�����n��@,ݾ;l������H2�� vI��   �   A~L������G5��LA����Ƚ���}�-��p�_���a�پ�����/�}PT�N�w�!w��Qᗿ��S�U���
����Ԍ��yz��	W��62�ѧ�J�ܾܥ�j�r��	/����"uĽ-���#h��ZCݽ`���C����W����Ͼw��G��&��c5��c?�()C��T@��+7���(����	� ���վ�����@���   �   �Ӄ�C����I�۽�5������ֽ����=��d���n���۾Fs	�$&��B�R[���n���{�<R����|�/�p�{�]�9�D��)�J$�i��錮�
҃�ZC������۽�5��7�����ֽ��)�=�g���q����۾�u	��&&�2B�[���n��{�VT����|��p��]�d�D��)��&��ྒྷ����   �   9ޥ�e�r��/������uĽh����e���?ݽ���	C�4���S����Ͼ;r��s��&�`5�O`?��%C�0Q@�@(7��(������ ���վ�����>���zL����	�	4��wA��W�Ƚ>����-�Ep�������پ�����/��ST���w�+y���㗿A����󢿗���/����֌�s}z��W�"92�ũ�B�ܾ�   �   H&˾+���r�Q���{Iս���&�������|ٽ;N�t�<�bs�@5��\9��ؓ׾]��I5�q��ׂ�L��"��i���'ݾzh��p����/��PrI�ZD��x�q����B���b���C߽��cS������fʾ��hQ.��Y�w�����Ŋ������CĿ��ǿ�Ŀ����c묿�� O���v[��/�����   �   Ŵ�k֮��v���)���H����D�����3��˽��S�+���W��͂��M�����@ٽ�+�Ⱦ��̾�>ʾ	��m����0I���e�U�:�2�����΅��['���q���������C�/��vz�BH��*b���!���P�:���x��������˿#�ݿ=��7�a��&�޿[:Ϳ�඿�e��	���FlQ�+�!��   �   ]w��<ɾWČ�%�?�YE �	��sz��xU��`��/���۳���8��	&4��T���p�U���ۨ���؎�&@��v��f�y��_���A�A�"�f�uսբ��뾐�f݈�d���t
Ž�
�uIH��I���̾Q��H�;���q�=~�������`ѿa��s���� �r_��H������c3ҿ�������Z�q�4�:��   �   �����5���<�S�,�
�c���7l��J-�����]4��g�"o���ýy�񽃢��%$�޸4���?���D��)C�l;��-�Q���v����7��2*��=F���f�Or�ʕ���Ͻ�n�p|^�5]��^�侺��ْR������j����ɿ��鿒��G�^��E�F������M�]
꿏�ɿ���� ��`Q��   �   ��(��>�:����c�6�������d����F���:��{�CB�[���ϡ�Uý4�ὢ��`����	�X	����"5��V�ܽ b����"��`���C��@��^��z���lٽ�"�Dp���f����h+���d����v��/nڿ�����D�0("��%�rD"�f;���������ٿ�3	���Nb��   �   �41�5��HO����m�տ��;��Zza�$��)������*"��X��M�1��Mg��{���������r,ɽ�@н��Ͻ��Ƚ����*���3<���)z�Q�o?1���!��)�`"T�D����$བྷ)�i�{������&4��=p�ws��Ln���忾�������!�@U*�`W-��[*���!����?����'�����%Um��   �   Q4�Ҙ����œq����㿽��`���������<�����Hټ�$��(I��z�0ۓ�w��s����c���u��������D��������va�=�A�!��Y���"��P�|A�����u+�/��"���ɾ��)7�::t�Y����¿A��X��*.��t$��.-��>0��,-�>_$����I����@���r��,q��   �   41�$���N����m�$���:��+ya�D
��(��ض���!��>��>�1�~Mg��{���������k,ɽ�@н��Ͻ��Ƚ����	���
<��|)z��Q��>1���!�1�)�@!T������#��)�P�{�$���*���%4��<p��r���m����4��T����!��T*��V-� [*�.�!����X?��!'���
��-Tm��   �   L�(��<�49����c����6�����d�^��(�ༀ9�y{�B�A���ϡ�Uý,�Ὑ��Z��|�	�J	�����4���ܽ�a�����!����`���C�8@��^�y���jٽG"�Bp�*쮾J���8g+���d�����t��mlڿ������ ��&"��%�C"�*:��������5�ٿ������Mb��   �   ������9�����S�V�
��`���4l��H-�&���\4���g��n��èýe��}���%$�ڸ4���?���D��)C�S;���-�'���v��佤���)��}D���f�+Lr�ȕ��Ͻ�l��y^�$[��s�侹��1�R�����sh��D�ɿ�� �2F����.C�z����L���1�ɿ���������P��   �   u�C9ɾ�����?�#C ���'oz�&vU�l�`�/��x۳����(���%4��T���p�S���ب���؎�@��h��A�y�ԭ_���A���"��4tսʡ�������ۈ����Ž��
�FH�yG��-̾��� �;���q��{������s]ѿ���d������H]��F�����Q��0ҿ���>���i�q��:��   �   ����Ү��v��)��������B������2���˽��9�+�}�W��͂��M�����?ٽ�(�Ⱦ��̾�>ʾ� ��X����I��Ƚe���:�������W���l%��Zo������ށ����/�uqz��D��	]�g�!�{�P����Yu�������˿��ݿ��迉�Ő�Ü޿O6Ϳ!ݶ��b��c����gQ���!��   �   =!˾����@�Q�H���Dս| ����,���{ٽ�M�E�<�bs�85��Y9��֓׾\��H5�p��Ղ�H����i���'ݾZh��H����/���qI��C�.w�w����?��#_��4>߽���]S�ҥ���aʾ���M.�v�Y�;��Z�������5���l>Ŀ��ǿk�Ŀ-���<笿�왿�K��q[���/�����   �   r٥�p�r��/������pĽ,����c��=>ݽ-���C� ���S����Ͼ7r��s��&�`5�O`?��%C�-Q@�<(7�و(������ ���վ����T>��mzL����2�m1���=��(�Ƚ�����-�*p����T�پ���^�/��MT�ڑw�0u��5ߗ���	������Ҍ�Ivz��W��32������ܾ�   �   �σ��C�����۽�1������ֽ5����=��d���n��
�۾Ds	�$&��B�T[���n���{�<R����|�,�p�u�]�.�D��)�:$�C�ྻ����у��C���2�۽O2��r����ֽ^����=��b���k����۾q	�`!&��B���Z���n���{�$P��o�|�5�p�ȕ]���D�)��!�}��Չ���   �   �vL�J���뽥/��i=���Ƚ`�����-�Ip�G���T�پ�����/�~PT�N�w�"w��Rᗿ��R�U���	����Ԍ��yz��	W��62����"�ܾ�ۥ���r�<	/�i���(rĽ����5b��#;ݽƖ�^
C�� ���P���Ͼ�m������&��\5��\?��!C��M@��$7���(���A� ���վy����;���   �   �@�s�ׄ���>��_��o?߽8��_S�x���dʾ5��O.�
�Y����&�������h����@ĿS�ǿ��Ŀq���W鬿��M���s[���/�B���#˾\�����Q�Ը�Fս� ��̢�������wٽ'K���<�]s�%2���5��v�׾e��2������`�V���c��-#ݾsd�����-���mI��   �   9��"���n#��~n��.���:�����/��sz�(F��W_���!���P�����v��¯����˿�ݿ���������޿_8Ϳ�޶�0d��ŷ��;jQ���!�b��Ԯ�
v���)�z�t����A������/��
˽��\�+���W��ʂ�cJ��@���ս���Ⱦf�̾::ʾ����d��<
F��ȸe��:�����   �   M���.���0ڈ�r��mŽI�
�DGH�zH���̾�����;�a�q��|������
_ѿp��^������\^��G����8���1ҿJ��������q���:�Kv�;ɾ4Ì�v�?�D ����rnz��sU���`��+���ֳ��齋���!4��T��p�8탾�����Վ��<��@��l�y���_��A�:�"���oս�   �   �?��f�-Jr��Ǖ�6�ϽXm��z^��[����侒��X�R�����ai��d�ɿ1����G�p��D�b��З��L�	�u�ɿ	������8 Q����<��L����S�(�
�Ea��x4l�"G-����"X4��g��j����ýS������!$���4���?���D�M%C��;���-�����s�Α�[��"&���   �   [�C��@���^��x���jٽ�"��Bp��쮾����g+�b�d�%��6u��2mڿ����h����~'"�<%��C"��:����̢��%�ٿM������Nb� �(� >�:����c����ૹ���d����r�༜3�sw��B���̡��Pý4��8z�������	�p	� ���/����ܽ�]��4ꢽ���d}`��   �   K�!���)�w T�K����#��)���{�Q���N��&4��<p�
s���m���l�����6�!��T*� W-�~[*���!�ؚ��?��俘'��Q���Tm��41����O����m���� ;���ya�
�8'��J���2��ظ�?�1��Ig��y���������)ɽ>н�Ͻ�ȽZ�̎��:��/&z��Q��<1��   �   �9$� �3�{�l�����}���UM����������!�d�_�M͔�f����뿾���W#��)8�yI��U�hCY��U�WI��7���"�������2���"����S\�����jݾ_*��ÍB�n�������B;��� �v��������$�� W�x���}ߣ�$q���(ҽRB�&������ڽ�1ʽE���B��������T�]{2��   �   ,2��<��q��}����mJ�!���N߾LR�*�[��e��Y���g���
��� �5���E��IQ�8UU��RQ���E�`�4�P1 ���	��,濹๿�����X��w�<�پL񒾖�?��z�l��_�@��
����!����=��Uu�ҝ���m���RԽ��l'��s �[���$��F���Ƚn��ܬ��.Um���E��   �   +�\�o"Y�Ό��Į�
��aB��<��^�ԾK��[Q��i���Ѳ��ݿb��b,,���;��iF�j2J��F��<�;,����0��R�ۿ����/��r�N�R+�%�Ͼ�����8�ȝ�*��A�Q��H)�U',��`O�X̄�\����н����b�P��
%��)��K'�$�����+�����츾�
��.���   �   �h��D���댽�}������a6�F���Eľ`����@�6~��a���F̿�2�� T���
�,��6�>�9�m6��5-�����%���˿�J��>9�*�>�w�	��h�����W�-��]�zÜ���o��-^�k.y��A��1wƽ����0�8	3��0K��^�nxk�f�p���m��c�.�Q��=;���!��c�`�ܽ�(���   �   ��ɽD��E���2l��@L�k!'���r�U���� ��S�+��5e��q���ն�%�ڿ�6�����A�._"�hZ%��"�h����zQ���rۿ����I��eld�-�*�����ɬ���l��. �W�ܽ�P��pގ��2�������Q���8�h�_�ゾ���hݡ�����U���<���J������Z���%i���B��I��T���   �   �A
�	ݽ f��Μ��4��M��U�؝��CN׾c8��E�M�~��m������=ܿ�������.��Xd��E�����_��c�ݿ����%��!��/�E�q��־jᖾ�]Q���dֽM���襯���˽�� �X '���U��_��>4���w����Ծ���������q ���]�h�ؾ�����!��Vz��-�_���0��   �   ��:���VX�M�н7
ݽ3L�q8�r��w��������2%��/U�
Ʉ�Ϝ���E���Ͽ;�Έ{�?��T��M�'�ѿ��������؅�v�V���%��T���u��rt���6����YԽ�Nƽ��۽���\�2���i�R$���T��K]�G��n��$#�� ,���/���,��$�����e�羺t������(�r��   �   	�w��K:������꽺ݽ^��|"��TU�����ȾÊ�zf,��&W�a���
ږ�Ϡ���w���¿Y�ſn�¿�͹�sH��;����'����Y��C.�e��9Yʾ����V����B��̎ؽ��l6
���4�k�p��О�8m̾�C���7�Q!4��PK���]��i��Wn���j�٭_���M��6� ��9��Ѿlʢ��   �   R���Lm���/�"���,�h�vS�w�,��ci�����'Ѿ���z(�:fK��9m����)����[���@��\�����������Wp��\N�+��	���Ծ�O��oIm�z�/���<,彻�U��,��gi�����B+Ѿ
���|(��iK��=m�C�������r^��KC������
���� ���[p�K`N��+��		��Ծ�   �   �[ʾ���6V�*���B����ؽx��94
�G�4���p��͞�<i̾�>�� 5��4��LK���]���i�!Sn���j���_�"�M���6�;��L7��Ѿ�Ǣ���w�I:����K���ݽ0��W$��WU������ȾҌ�i,��)W�O���?ܖ�?���<z��� ¿�ſ"�¿_й��J��T���e)����Y�MF.�8���   �   ^W���w���u��i6����{YԽ�Lƽ	�۽#����2���i�!���P��xX�BD��k�!#��,�Q�/�V�,���$�܏�Z��Ŋ��p��������r���:����U�<�н�
ݽLM�s8���ڊ��Գ���4%��2U��ʄ�Ԟ��H����Ͽ���a~���sW�fP㿕�ѿ���g��|څ���V���%��   �   ���־�▾}_Q�<�dֽ쐱�)���h�˽�� �d�&��U��\���0��-s���Ծʠ�V���	������MX뾢�ؾp���h��bw����_�:�0�?
��ݽd��=�����KN�-�U������P׾:�@�E��~�Qo�������ܿ��� ������e�XG���b��|�ݿi��q'������E��   �   o�*�ژ��"ˬ��l�Y/ ���ܽ�O��f܎�q/��D���潄��^�8�ވ_��߂�����١�����0���8��(G��&��?��l i�5�B� F�?O���ɽ������l��PM콫"'���r�򞯾#����+��7e��r��[׶� �ڿ�8����bB��`"��[%�Z�"����(��_S��qtۿ�	���J��nd��   �   .�>�.�	��i�������-��]����o�C)^��'y��=���qƽo���-��3��+K���^��rk���p���m��c�S�Q��9;���!�x`�q�ܽ(%��,f��^B���ꌽ�}��΢���6�7���rFľe����@������'H̿54���T���*�,�$!6�r�9�Fn6��6-������W&���˿�K���:��   �    �N��+���Ͼ���x�8��� ��I�Q��E)�#,�[O��Ȅ�����н<���~_�����%�j)�DH'�������v��/�������`����\�L Y����Į��
��bB�@=��{�Ծ��\Q��j���Ҳ��ݿ����*-,���;��jF�T3J�ȓF��<��;,�B������ۿG�������   �   X�X�x�u�پi񒾪�?��z�Bl��>�@�K�
�^ ��E����=��Qu�_����j���OԽ��� $��Yq ��������`�6�Ƚ5�����LRm��~E��*2�%�<��q��}��z���J��!��DO߾�R���[�_f��ۡ����F�
�� ��5�t�E�JQ��UU��RQ�8�E���4��1 ���	�-��๿�����   �   kS\�����jݾ6*����B����q��OB;�"� �������P�$�E W�P���Xߣ�q���(ҽ:B���۲���ڽ�1ʽ'E���B������+�T��{2�(:$�Z�3��l������UM�΅�����!���_�k͔�����6������W#�
*8�yI��U�jCY��U�WI��7���"��������������   �   u�X�pw���پ����?�ey�k��E�@���
��������ۛ=��Qu�X����j���OԽ��� $��Xq ������N�#�Ƚ��ઐ��Qm�~E��)2�W�<��q�
}����-J�� ��PN߾R���[��e������翶�
�f� ��5���E�"IQ��TU�RQ�\�E���4��0 �b�	�4,�?๿'����   �   l�N��*�	�Ͼ䅌��8�̛�R����Q��D)�X",��ZO��Ȅ�����н:���_�����%�g)�?H'�������`�����Ŵ����������\��Y�ȉ�Hî�`	�aB�<����Ծ̡�YZQ�si��5Ѳ��ݿ��v��+,���;��hF��1J��F��<�D:,������Z�ۿ�������   �   ��>�w�	�g��
�����-�[�������o��'^��&y�f=���qƽU��� -��3��+K���^��rk���p���m��c�>�Q��9;�ӹ!�I`� �ܽ�$��de��LA��H錽�{������26������Cľ�����@��}��|���E̿F1��4S� ����,��6��9��k6�v4-������#����˿�I���7��   �   ��*���DȬ�,�l��, ���ܽ\M���ڎ��.��������m��N�8�ֈ_��߂�����١�����/���8��!G����.��B i���B��E��N�� �ɽj��~��ni���I��'���r���������+�4e��p��gԶ���ڿ�4������?��]"�Y%���"�&����gO��qۿ���H��Zjd��   �   ����־�ߖ�<[Q�[�1`ֽe�������e�˽�� �5�&�f�U��\��0��.s���Ծ̠�W���������EX뾕�ؾ\���Q��Dw��3�_���0��>
�&ݽb��g�����GK�űU�V���-L׾�6��E���~�l��*�'ܿ0���Z������b��D�<��A]��%�ݿ���B$��_����E��   �   6Q��s���r��6�����UԽDJƽd�۽���H�2�{�i�!���P��wX�CD��k�!#��,�Q�/�T�,���$�׏�Q������p������4�r��:����S�^�н�ݽ:J��n8����S��������0%�D-U�|Ǆ������C����Ͽ����x�i���Q�
K㿞�ѿ�����
��9ׅ���V���%��   �   VʾN��@V���@=��2�ؽ ��n3
�ͫ4���p��͞�2i̾�>�� 5��4��LK���]���i�"Sn���j���_��M���6�1��>7��ѾsǢ��w�nH:�������{ݽG�� ��QU������Ⱦ��d,��#W������ז�{���u��>¿��ſ��¿1˹�F������%��D�Y�EA.�Q���   �   �L��Em�#�/�W��v'���VR���,��ci�䱝��'Ѿ���z(�<fK��9m�
���,����[���@��]�����������Wp��\N��+��	���Ծ}O���Hm���/�����(�P�$Q���,�2`i�y���?$Ѿ���`w(��bK��5m�禅�ؔ��~Y��A>������H�������Sp�}YN�+�7	��Ծ�   �   �w�FE:����E��/{ݽX���!�TTU�m��e�Ⱦ���vf,��&W�b���ږ�Ѡ���w���¿\�ſo�¿�͹�qH��8����'��{�Y��C.�T��Yʾm��V�����>��	�ؽ,�㽛1
��4�h�p��ʞ��e̾T:��42��4�IK�~�]�p�i��Nn�N�j���_�F�M�:�6�:���4�� ѾmĢ��   �   ^�:�B�\P轰�нbݽ�J�6p8�4��S���r����2%��/U�	Ʉ�Ϝ���E���Ͽ=�Ή{�@��T��M�%�ѿ��������؅�m�V���%�kT��\u��"t��6�����UԽ�Hƽ��۽M���2���i����L���S⾖A��h��#�{,��|/���,��$�����������l�����M�r��   �   �;
�*ݽ�_��B�����L�a�U�����*N׾\8��E�K�~��m������>ܿ�������.��Zd��E�����_��a�ݿ����%����%�E�c���
־,ᖾ;]Q�r��`ֽ����e�����˽�� ���&���U��Y���,��o��Q�Ծ������ry��d���S뾹�ؾ	������/t��A�_��0��   �   ��ɽj��J|���h���I콦 '�=�r�3���� ��Q�+��5e��q���ն�&�ڿ�6�����A�0_"�jZ%��"�j����xQ���rۿ����I��]ld�#�*������ɬ�!�l��- ���ܽM��jَ��+�����U������8���_��܂�~���ա�������3��CC���{������i�g�B�+B��H���   �   Ub��"?�� 茽/{�������6�����DľZ����@�5~��c���F̿�2�� T���
�,��6�@�9� m6��5-�����%���˿�J��:9�"�>�l�	�lh��蟂���-��[�������o��#^�]!y��9���lƽA���W)�~ 3��&K�M�^�Imk�	�p�U�m�.c�P�Q�5;��!�]���ܽv ���   �   ��\��Y����®�y	�vaB�g<��R�ԾG��
[Q��i���Ѳ��ݿd��b,,���;��iF�j2J��F��<�;,����0��R�ۿ����-��o�N�L+��Ͼ������8����v�����Q�B)��,��UO��ń�;��
�н����\����,%��	)��D'�z��������(�㽭���X��<���   �   �'2���<��q��|��׭�CJ�!���N߾KR�,�[��e��Y���g���
��� �5���E��IQ�8UU��RQ���E�`�4�P1 ���	��,濸๿�����X��w�4�پ<�g�?�	z��k��
�@���
��������=�Nu�6���<h���LԽ���� ���o ��������U�t�Ƚ���ܨ���Nm�r{E��   �   �>�[�P�~É��˽.��2�p��ε�t���B?�mჿ�	��O�߿�	
�4l%��*A�|�[�V�r�,��������\r�dC[�NU@�hX$�����cݿK���"��S<�Hb��s����h���@����+u��>2����01���Z�2ۉ�0ʩ��ɽ�E� M���R��}	�������R�BԽV6�������x�jO��   �   RO���[�S�����˽�D�b�m����*���$<����=>���!ܿ�����"���=���W���m�*}��:��P}���m��bW�R,=�b�!���� ڿ�Z������Y9�T�̮���e�B����}4{�6=�5�0�%|G��Vw��[�����fm�'o �V
��k����~�������]5�˽�#��2O����e��   �   ����b}�H`���̽�8�5d�0𪾣���N3�Bw�b����ѿ��>���[4��LL�`��vn���s���n�F�`��^L��4��s��� ��Yп힢�GXt�ʳ0����#��f]�\B�j���/���`���c��
���l���ѽ�L���q��|)���9�H'D��aH���E�4�<�q.��������޽h����   �   �5��A ��~N��b<Ͻ&l�ZV�Ņ������ %�"�c��f��+����p���t&�"D;��M��Y�V�]��zY���M�>�;�FI&��	������Bo��{�a��-#�K3�#S��(�O�2��m½���z$��x坽�c���S�1I�L�6�V�U���q�H���t��^O��b��ޅ���v���[��=�Kg��� ���Ͻ�   �   3�	�ǽ���0�ս�,���D�����GϾk3��K�3���w��ֿͅh) �Ja�v�&�L�5���?�n�C��j@���6���'���Ҏ ���ֿ�J���Ɔ�C�I�	���̾����
�?�P��:�ʽ���?ߺ���޽�x�}�1���\�<F��ꛛ���������/Oʾ�RξWe˾���k����䈾=ld��H9�Z���   �   9"���_��2�����G�2��8|��=��f����C/���i�>���8����޿B� �@�^�d%��(�0�%���j�����~$���+�����i���.�!]���Ĳ���x��.�ٻ�&$ٽ&Z׽o�����cH�2P�����
���D�߾"j��]�	�F���l��
�
�E����s�E�þ�����p��\_O��   �   T�[�ٟ)�b8	�ã���!��!��2Z�"����վJ���`C���{�vs��ڙ��kTٿV��*?�\�Z�����'������Yۿc>�������:}��*D����Iuվ{��bX��� ��a�:��T�$�ڻU�!V���y��Lf޾>������0�P�@��{K��eO��VL���B�S�2���ӓ�;��qe������   �   ,͑���[�<�(��a����*
��:�0�|��.��B��&�&�K� ~�F͘�r���2ǿ|bؿv��3���w俰�ٿ�ɿ�Z��0w���]����M�c[��o ��@]}�FI:����]����%�uwW�K-��d���؀�)N�P�6�U�@p�\傿�艿{����v���胿��r�z�W�K\9����G���տ��   �   ,+��N
���O�
K �����d��$�h�M�T�������h������iG�Yhp�u����x���P���P��
�������������͢��s{s��I��!�����V(��X����O��I �`���e�}&�w�M����� ����������ImG�nlp�����b{��gS���S������n
��K���0�����Rs�AJ��!������   �   2ﾢ��`}��J:�������,�%��sW��*����&|�=K�Ѥ6�U��;p��₿,承职�It��!惿��r���W��X9�������ѿ��ʑ�F�[�/�(��`����0�	�:���|��1�����A�K��#~��Ϙ��t���5ǿ�eؿ���e���z俩�ٿ�ɿm]��Ky��{_����M��]��   �   /���wվ ��CdX���� ��_�2��6�$�w�U�/S���u���a޾.;�6��,�0�L�@��wK��aO��RL���B���2���������a��h���f�[�,�)��6	�o����!�+�!�Z5Z�����վ?���cC���{�uu��1���WٿK���@�����()�a���\ۿ�@��s����=}��,D��   �   8�.�o_��nƲ���x���.�ܻ��"ٽW׽1j�����_H�HJ�켞��|��$�߾^d��=�	��B�@�'����
������n��þt���n��$[O��5"�
�����x��A����2�;|��?��F����E/���i��?���:��"�޿�� �������e%�؂(���%�&�Ґ� ���&��������#�i��   �   ��I��6�̾������?�p��,�ʽ����ۺ���޽{u��1�T�\��B��$���p������\JʾNξ�`˾����B{��-잾�ሾgd��D9�.���z��ǽR����ս�-�E�D�����IϾ�4��K�=4��y����ֿ|* ��b��&���5�Z�?�(�C��l@�8�6��'���ď ��ֿ�K���ǆ��   �   ��a�t.#�l4��S����O�22��l½k����!���᝽�^���M�_E���6��U���q����q�� L���^���څ���v���[�=��c��� �.�ϽO2��'���xM��n<Ͻ�l��V�݆��<���%�ªc�h��y���7r����&�hE;�NM�hY��]�v|Y��M�b�;�8J&��
���!	��p���   �   Yt�Z�0������#���]�rB�񌾽
��R
`���c�����h���ѽ�F��Jn�y)��9�$#D�f]H���E�S�<���-�`�"���޽����씽��_}��_��$�̽9�,6d������;3��w�.����ѿ������h\4��ML��`�xn��s�įn�J�`��_L�t4�:t�H� ��Zпt����   �   ���Y9�4T�=̮���e�6�����53{�E}=���0��xG�sRw�Y��8���)j�^m �j��i���������4��V2�z˽a!��xM���e��O���[�4�����˽E�!�m�J�����*%<�f����>��z"ܿ<��(�"�J�=�:�W�(�m��}��:���}�B�m�RcW��,=���!���mڿ�Z���   �   �"���R<�(b��s����h���맼�c+u�>2�z���1�*�Z�ۉ� ʩ���ɽ�E� M���R��}	�������X���BԽc6������x�CjO�l�>���P��É�n�˽k����p�ϵ����%C?��ჿ�	��u�߿�	
�Jl%��*A���[�f�r�1��������\r�TC[�:U@�VX$�����cݿ+���   �   ���Y9��S��ˮ���e�������"2{��|=�/�0��xG�NRw�Y��5���,j�\m �l��i���������.��D2�c˽A!��UM����e�O���[����� �˽tD��m������^$<�ܽ��>���!ܿ���z�"�t�=�6�W���m��}�/:���}��m�XbW��+=���!�����ڿGZ���   �   Wt��0�����$"���]�<A�\���	��	`�֊c�P���h���ѽ�F��Jn�y)��9�)#D�h]H���E�N�<���-�Q�����޽���b씽h���^}��^��s�̽�7�A4d��諭�����3�rw����D�ѿ|������Z4��KL���`��un�|s�r�n�0�`��]L��4�s�J� ��Xп)����   �   �a�n,#��1��Q��L�O��0��j½ ���� ��8᝽D^��uM�SE���6��U���q����q��L���^���څ���v���[���=��c��� ���Ͻ�1������K��:Ͻ k�V�����O����$��c�)f�� ���Yo�,�~&��B;��M�bY�ʀ]�vyY�$�M� �;�6H&���X�����?n���   �   l�I�� ���̾Q���Ͻ?�l����ʽ����ں�!�޽Pu���1�E�\��B��&���t������`JʾNξ�`˾����;{��"잾�ሾ�fd�WD9����y콬�ǽo���սj+��D����RFϾP2�rK�2��Iv��7�ֿs( �(`�$�&���5��?���C�Di@�&�6�*�'���ō �ÿֿI��Vņ��   �   ��.�7Z���²���x���.�����ٽ0U׽i��S���^H�0J�漞��|��&�߾cd��?�	��B�A�'����
������n��þ[����m���ZO�}5"�V����b����;�2��5|��;�����,B/���i��<���6����޿
� ��}���^b%�d(�~�%�����v��6"�
������\�i��   �   ���^rվT��>_X�z�D ��\�F����$�$�U�S���u���a޾-;�8��/�0�P�@��wK��aO��RL���B���2���������a��=����[�v�)��5	�Q���u��!�70Z�O�����վ����^C���{��q�������Qٿ���=������v��&������Vۿ<�������7}��'D��   �   Pﾬ���Y}�F:����z����K�%�sW�p*������|�;K�Ф6�U��;p��₿.承ꁌ�It��惿��r���W��X9���ˇ���ѿ��ʑ���[�-�(�_�q����$�:���|��,�������W�K��~�1˘��o��0ǿ�_ؿ_���翜t俩�ٿɿlX���t���[����M��X��   �   �$�������O��F �����b�j#���M��������W������iG�\hp�w����x���P���P���������������ˢ��l{s� �I�r�!�����#(������O�`H �T��|b�"��M� �������t�������fG��dp�@�Rv���M���M��!������Ɩ����t���Zws���I���!�V����   �   �Ǒ��[���(��]���s�Α:���|��.��(�� �$�K� ~�G͘�r���2ǿbؿy��4���w俯�ٿ�ɿ�Z��-w���]����M�T[���. ��v\}�H:�� �e�|��/�%��oW�(��`����w�H���6�8U�:7p������㉿\���q���ヿ��r�|�W�iU9����!����Ϳ��   �   ��[�r�)��3	�P���X�z�!�2Z�ߧ����վB���`C���{�ws��ܙ��mTٿY��,?�^�\�����'������Yۿ_>�������:}�w*D�t��uվ(���aX���r �5[����$�6�U�hP��br��]޾{8�����0�g�@��sK�_]O��NL���B���2�m
�4�����]��U����   �    2"��������}��� �2��7|�[=��L����C/���i�>���8����޿B� �B�`�d%��(�0�%���j�����{$����'�����i���.��\���Ĳ��x���.�
���ٽ�R׽�d��B���ZH��D�u���px��<�߾�^��3�	��?��������
�Թ��ji㾌�þ�����j��GVO��   �   �t�&�ǽC
��-�ս�+���D�i���GϾb3��K�3���w��΅ֿh) �Ja�x�&�N�5���?�p�C��j@���6���'���Ҏ ���ֿ�J���Ɔ�:�I�����̾y���!�?����/�ʽ6��q׺���޽.r���1�-�\��?������[��������Eʾ*Iξ�[˾����w��^螾�ވ�|ad��?9�{���   �   �-������TJ��{9Ͻ-k��V�����x��� %�!�c��f��,����p���t&�"D;��M��Y�X�]��zY���M�<�;�FI&��	������?o��u�a��-#�+3��R���O�1��j½�������ޝ��Y���G��A�w�6�!�U�O�q���bn���H���[���ׅ��v�b�[�'�=��_�p� ���Ͻ�   �   ����Z}��]���̽�7��4d�𪾕���L3�Aw�c����ѿ��>���[4��LL�ė`��vn���s���n�F�`��^L��4��s��� ��Yп랢�BXt�ĳ0�Լ���"���]��A���������`��c����e��SѽzA��4k��u)�<�9�'D�NYH�r�E�j�<�9�-���;���޽����J锽�   �   �O���[������˽fD�4�m����&���$<����=>���!ܿ�����"���=���W���m�,}��:��P}���m��bW�P,=�b�!���� ڿ�Z������Y9�T�	̮�\�e�������1{��{=�|�0�$vG�Ow��V������Ggὼk ����g���������s��"/콨˽���dK����e��   �   �]�`�q��^������2�`!���DϾ"��x;Z��7����ƿW���H��T=���^��;��v׎�:��Dy��Aޘ�����Z����]���;���}S����Ŀ#����zW����b�˾k��K1-�}�޽̾����^��%J�u$]�2����R����Ƚ ��2���g�$�����.��r��k������нh��掽��o��   �   :�o���}�����8齈�0�VJ��
̾$T�n�V�-Γ���ÿo����Q���9���Z�DT{�/ы�S�����������Ƌ�F�z��Z���8��)���������1���T�+8�J�ȾY����+�96߽N��rk��\�32v������������g�L���"��+��U/�P�,��$�������_���� ����z���   �   ,"������æ��e�Yv,����j�¾8��kL�eˌ�����3�L���0�x&O�z�l��R��Q6��r��!X���y����l���N�*
0��F� ������v���0J�.^��Ϳ�>�~�Q�'�0���s������Ɗ��w���ƽ�\�������,��HC��"U���`�ZOe��b�s�W���F�{�0��b�֤��hGн��   �   �YŽ�3���ֽ��P�_&�xt��ʹ��1��h<�>ԁ��L���'ܿ���
�"���=���W���m��}�GW���}���n��FX��>�h�"�0��HBۿ�Q���〿�:����5���To���!�Z�佐+���F���������&v/�l"S�B$v�Nʊ��W��M��������M������� �z�� X�9v4�]�l���   �   �s�佒ڽr �����`�kB��ı�((�,�g�C��K/ſ$v�B}�v�(���>�0�P�Z]��b���]�L�Q���?��)����S��ſ���~�f��'����F���\��^��d��ҽ�8ܽ{��K#���M�F~~�~��{���Eɾ&z۾�`���{O�U6ݾ�˾ *��R��	���R�A(��   �   9�֕��W����^�+L������;r��?H��M�����Ւӿ�����Q��[$��3�|=�F�@�(�=�f14�r�%�Z�WI���pԿn���X����G�o����̾�����ZI��c�YL��r�����H4��g�gʒ��<��X�۾* �J|�̑�&�C)�c�&�3��w��־���޾�r������j<l��   �   �cz��A�J����Nb���8��y�����)���'�):_�-������T(տ4���p=
�6,���� !����,��e�����`�ֿ�H��P��[�_��'�Q�����!x�_#7��=��u�z�r	>�Y�u����̾y������Hk3��UJ�y�\��bh���l�]5i��
^�)FL��5����tX��Ͼ�����   �   "S��g�z��A���	n���(�"�U������NǾ���L�4��i�����/���ɿ�6�<�����u�ԕ��A��':��˿�����?��!�j�6������Ǿ㐾��U��(��0�����>���w�8;���ؾ��
�Z@-���P�&�s�����?��;!���	������@A��a���4v��|S��m/�����ھ�   �   �׾o쟾�ym�s�7��C�O��]�6�P�k�b����"־f����6�s�c�;����@��w�¿Y�̿S�п8�Ϳ�Ŀiⴿ�5�������mf�E�8��@���׾0ꟾ�vm���7�uC� �e�6���k�����V&־�����6�T�c�g=��e����B����¿��̿��пw�Ϳ�"Ŀ?崿58��ʼ���qf�.�8�9C��   �   ]��d�Ǿ�䐾��U�t(�H0�����>�N�w�$8���ؾ�
�=-���P���s�5��"=��]����� ����>���^��z0v��xS��j/������ھ`P����z���@����n� �(���U������QǾ����4��i����������ɿ�9⿪���Y��v����YE��==�ʹ˿����A��V�j��6��   �   ��'����S��-x�9$7��=��t�4��>�a�u�� ��ʶ̾���n���g3�NQJ��\�^h��l��0i�>^�BL�^�5�k���U��Ͼz���2_z���A�r
�*���b��8�l�y����'-��N�'�=_��������*տ7���?
�.����!���x.�>g�������ֿ�J���Q����_��   �   ��G����D�̾�����[I��c��J������V��g{4�ug�
ǒ��8��O�۾; ��x�:��M&�F?)���&����<�������޾�n��b����7l��9�{��nV�.���^��,L�6����;�s��AH�O������ӿ2����S�z]$��3��=�\�@�,�=�@34��%�t[��K���rԿ�o��Z���   �   .�f�'���꾻G���\��^�zc�7ҽ�4ܽ�|�H#��M�x~�����v���@ɾ�t۾u[羃���I�$1ݾ"�˾�%���웾���O�R��=(�l���佲ڽ ������`��C���쾣)(�K�g����1ſ7x�~~���(�L�>�"�P�8\]��b���]�$�Q�4�?�p�)������|ſ8����   �   p䀿�:�N���5���Uo���!���佼)���C�����T �Z��q/�FS�Nv��Ɗ�T������'����I��]���J���V�z���W� r4��^��@VŽ1���ս�Q�&��t� ϴ��2� j<�*Ձ��M��B)ܿl�� �"�D�=�6�W�N�m��}�GX����}�b�n�bHX��>�N�"���nCۿ�R���   �   2w���1J��^�Jο���~�n�'�����r��!���Ċ�Pt����ƽ+W��b����,��DC�CU�I�`��Je�b�	�W���F���0��_�����MCнf몽���\���"������v,�Y��h�¾�8��lL�̌�����$4���l�0��'O���l�kS��7���r���X��z����l�Z�N��
0�@G���f���   �   :1��<T�R8�u�Ⱦ"Y���+��5߽���=k�(�\��.v�`������p��e�E��ì"���+��S/��,���$������\轓���2���:y��3�o���}���������0��J���̾�T��V��Γ���ÿ��� R�d�9�n�Z� U{��ы�Ð��@�����ǋ���z�"Z���8��)���������   �   ���[zW�[��+�˾@��1-��޽|����^�(%J��#]�����bR����Ƚ������g������*��p��n������н~��0掽�o��]�ӛq�_����Y�2��!��$EϾM���;Z��7����ƿ����^��j=���^��;���׎�?��Ey��>ޘ�����F����]���;���WS��s�Ŀ�   �   �0��]T��7���Ⱦ�X��3�+��4߽����k���\�4.v�F������v��e�H��Ƭ"���+��S/��,���$������\�|������y����o���}�������?�0�0J���̾�S�1�V�Γ���ÿ����Q���9�f�Z��S{��Ћ��e��F���MƋ���z�&Z�
�8�F)��������   �   v���/J�p]��̿���~��'��བq��j����Ê�
t��j�ƽW��^����,��DC�LU�O�`��Je�b�
�W���F���0��_�����
Cн몽b������狼��
꽌u,�F����¾�7�7kL��ʌ����;2����0��%O�d�l�R���5��Wq��^W��'y����l���N�^	0�F�������   �   �‿��:�����3���Ro�ޟ!�)��,(���B��������D��q/�ES�Rv��Ɗ�T������*����I��\���F���H�z���W�r4�����UŽ0���ӽ�{N�&��t��̴�1��g<��Ӂ��K���&ܿ����"���=�4�W���m�
}�KV��"�}��n�pEX�R>�\�"�T���@ۿ�P���   �   j�f�P'�͖� E����\��\��`�_ҽ�3ܽ6|��G#��M�x~�����v���@ɾ�t۾|[羉��J�$1ݾ�˾�%���웾����R�9=(�����佰
ڽ
���/��`�&A������&(�s�g� 
���-ſZt�*|�"�(���>�Z�P�X]���a���]�`�Q��?���)�|��Q��d�Ŀ���   �   ��G�����̾Ū��+XI�=a�{G��������{4�>g��ƒ��8��M�۾> �y�>��Q&�I?)���&����9�������޾�n��F���I7l�&9����UU�����[��(L�V����;�p��=H�QL����ݐӿ5����P�Z$��3�|=�4�@��=�|/4���%��X��F��enԿIl��jW���   �   ��'� ��&	��~x�p 7�D;�&s�2�R>��u�� ����̾
���o���g3�SQJ��\�^h��l��0i�>^�BL�Y�5�d���U���ϾP����^z�G�A�V	�z��`�7�8��|y��}��'��"�'��7_���������%տg����;
�t*��
��� ����*��c�������ֿFF��HN��o�_��   �   p����Ǿ����%�U��(��-�`�ʡ>���w��7���ؾ�
�=-���P���s�7��%=��`�����!����>���^��v0v��xS��j/������ھ'P���z���@�E���k�L�(��U������KǾ�����4��i���������\�ɿ�3������Bs����>���6�)�˿���g=����j�P 6��   �   ��׾Y矾�rm���7�x@�"����6�v�k�"����"־^����6�r�c�;��Ċ��@��{�¿]�̿U�п;�Ϳ�Ŀgⴿ�5�������mf�:�8��@���׾�韾�um�|�7�7A����l�6���k�Ⱎ�L־'����6���c��8��D���8=��p�¿)�̿�п��Ϳ�Ŀ{ߴ�3��H���jf��8��>��   �   M����z���@����$k���(���U�����vNǾ���F�4��i�����1���ɿ�6�A�����u�ԕ��A��':��˿�����?���j�	6�y����Ǿ�␾x�U��(��-�5�i�>��w�=5���ؾ��
��9-���P�6|s����y:��������F����;��\���+v��tS�Rg/�ީ�v�ھ�   �   �Yz�إA�!�V���_��8��~y�����)���'�':_�-������U(տ8���r=
�8,���� !����,��e�����]�ֿ|H��P��Q�_���'���?��x��!7�z;�Xr�V�F>���u�������̾����[���c3�?MJ�z�\�VYh�A�l��+i��^��=L���5�#��$S���Ͼ�����   �   S�8����S����\��)L�g��z�;r��?H��M�����֒ӿ�����Q��[$��3�|=�F�@�(�=�d14�r�%�Z�UI���pԿn���X����G�[��C�̾ ����YI��a��F��0���^���w4��	g��Ò��4����۾p ��u���&��;)��&������
����޾�j��� 2l��   �   ����8ڽ����`��`�#B�����((�)�g�C��L/ſ%v�B}�v�(���>�2�P�Z]��b���]�L�Q���?��)����S��ſ���w�f��'�ߘ�sF���\�;]�+`�tҽ0ܽ�y�QD#�J�M�?r~�C���r��(<ɾ�o۾V���뾇D��+ݾL�˾w!���蛾���'�R�`9(��   �   pQŽ(-��(ҽ��M�L&��t��ʹ��1��h<�>ԁ��L���'ܿ���
�"���=���W���m��}�HW���}���n��FX��>�f�"�0��GBۿ�Q���〿�:�����4��5To�~�!�&���&��z@��\������m/�iS��v��Ê��P��ԇ��_���F��ȵ������a�z���W��m4�n	�m���   �   �������ã��N
꽧u,����L�¾�7��kL�eˌ�����	3�L���0�x&O�z�l��R��Q6��r��!X���y����l���N�*
0��F� ������v���0J�$^��Ϳ�Ξ~���'����p�����o����p��j�ƽR��[��`�,��@C��U���`��Ee��b��{W���F�+�0��\�����>н�窽�   �   �o���}�E���5�1�0�<J���̾ T�n�V�-Γ���ÿq����Q���9���Z�DT{�/ы�R�����������Ƌ�D�z��Z���8��)���������1���T�(8�<�Ⱦ�X����+�55߽���~k��\�|+v�z����󸽨�Xd�q��ª"���+�bQ/���,���$����Q��Y�������Gw���   �   �x��������'� �RE�&��*����(��p��K���wڿ�U���,�N�Q�Lz�K@��oڢ��ͮ����"Ȯ�0���'��<y�̨P��+��9
�1�ؿeУ��<n���&���� �}VA��`��|��4���t*m�܀��(����⽏C��P�#�"�8�+��/�Nu,�bJ$��D�������r���q���⍆��   �   dd���F�����0
�zFC�["���	�n�%��l�����׿�$	�f�)�N� u��'��b;��Nߪ�������*0��<���Wt��M��(�P"��Rտ�F���zj��$�/a޾����7�?�v���������l���D{��d]����ѽ��������%�Ի4��x>��B�D?�p86�j�'�ej��� �?׽���l;���   �   �T�����B��L���c>��Z����־����ia�����ͿV��z�!�0|C��Cg��t��������0���ٟ��+���~����f���B�!���q�˿����Í_�|���ԾFe��.;�I-���C��zN��F���X?��f�ོ�	�b%�ޅ@���X��6l��x��}}���y�d�m��([��=C�dT(����:��f-���   �   �۽�Pǽ>�ҽBx�f7�̔���oǾ����O�e���������X���3���R�Nwq�v��c8��)���vw���c��6r��#S���3�B�;񿧦��@���uN����kvž�䄾}e4�� ��yͽ����x1ս�l �,%��C�ÿj�����OÙ�Zz���h��w������х��:*���,��A-n��G��r"���   �   f������M��`�/��w��$����@�9�y��
�����ؿ���R) ���:�J�S��ri��Cx���}���x�Hnj�P�T��n;��� �d���ؿ�?����~�$�8�D�������0u��T-��;������l_�/[6�
�d��M��Lʩ�ӵž��޾?������@�,@ �B�����ĿǾ�᫾�Q��j�h���9��   �   :L��K$��A������)�O�a�����r\�I� �]�q����G����"�
��#!�"�5�yF�V�Q��=V���R���G�n�6�`"�����b�p�������\�89 ��e⾂�����_�&�'���J����!��I��e���ۢ���ɾL;�������5.�܉7���:��
8�)!/�O
!�%������l̾����<���   �   ��b�U�&�-�?���&���L�׉�����T���#9��pv�K��Ŀ�i������r%�"L.�p�1���.�Zc&��1������뿍ſ�ힿ�w�r^9�����r���R��F@K��
%���ݤ+��RS�9���{e��o�⾕(��3*�]pF�ț_�g�s�c:���������k�t�r;a�7/H���+����O�Wh���   �   ����[��&NU�'�0���'���:��l������bܾ+K���G����ݟ���C�ݿ�����������y�0\����-�����߿�������jq���H�>���ܾ�"���`l�.g:���&���/���S��6���뵾�Kﾬ���?�3�f��v���A��'������-��<����_���Y��Ú��pi��vA��0��q��   �   i����3��8gK�qa.�2.���J�������������:J���{��m��Mկ��Wſ�Hֿ�@�MD����(w׿��ƿHI��[���E�}���K�P�~e�C���.2���eK�a.��2.���J�����a���"����.>J���{�xp��.د��Zſ>Lֿ]D��G�y�ῇz׿��ƿL��¹��D�}�/�K����   �   ?����ܾ�$���bl��g:�Z�&�ŷ/�~�S� 4��x赾bGﾸ��h�?���f�t��?��'}��g���)������\��W��T���?i�1sA��-�\m��|���Y���KU���0�~�'���:���l������eܾtM���G����hߟ�����h�ݿv����������{�(^�x��������߿ �����,s����H��   �   �`9�n���t���S��9AK�t
%����b�+�OS�|}���a����⾘%��/*�6lF�$�_�c�s��7�����i���z�t��6a�.+H��+���HK��d����� �U��-�+>�J�&�&�L��؉�������&9��sv�M���Ŀ�l꿪��� ��t%�RN.���1��.�Ze&�R3����p���ſY�w��   �   !�\��: ��g⾭�����_�0�'�5��d����!�I� c��Eآ�^�ɾ�5���T��1.���7�`�:��8�G/��!���)���8h̾����9��.6L��H$�@�e��&�)��a������^�� ��]�����I��|�返�
�D%!��5�X{F���Q�J@V� �R��G�L�6��"�ܨ�e�0���Q���   �   f�~�y�8�(��ҧ��
2u�&U-�;�K��J���<\��V6���d�UJ��5Ʃ��ž��޾n�������=�%= ����S��"�Ǿޫ�BN��?�h���9�*c����u�����/���w�\&��!����9�ʛ�������ؿ����* �H�:�J�S�ui�0Fx�R�}��x�zpj�.�T�tp;�Ē �^����ؿ�@���   �   �@���vN�E��Nwž儾�e4��� � xͽ}����,ս�i �S!�b�C��j�]�������]v���d��9�������ၨ��&��_)���'n�VG�Uo"�����۽YNǽ��ҽEx��f7�����,qǾ�����O�f���]��Y�̋3�t�R�.yq�����9��]����x���d���r�@%S���3��񿣧���   �   zᙿz�_����|�Ծ�e��N;��,��sB��_L��N���x;��y�ཻ�	�~^%�Ɓ@�e�X��1l���x�Rx}�ݶy���m�$[��9C�Q(��������)��WR��o�����l���d>��[����־W ��ja�q���Ϳ���>�!�(}C�Eg��u���������!����ٟ�P,��N����f���B��!���˿�   �   �F���zj�$�^a޾����,�?����D��w��ঀ�Dy���Z����ѽ.�������%�p�4�dv>�'B��A?�!66�O�'��h�� �b<׽����9��Hc��KF�����_
��FC��"��p
���%���l�����׿%	���)��N�� u�(���;���ߪ�-�����0�����BXt�M�F�(��"��Rտ�   �   DУ�<n�ҽ&�X����=VA�L`���{��켁��)m��ۀ��~(��~��vC��P��"�'�+��/�Gu,�bJ$��D����罂����������^�x�܈�����]� ��E�J&��o���(�J�p��K���wڿV���,�l�Q�lz�Z@��zڢ��ͮ����Ȯ�'�����"y���P��+��9
��ؿ�   �   F���yj�o$�t`޾���c�?� ������������y���Z����ѽ/�������%�u�4�iv>�+B��A?�"66�M�'��h�� �L<׽~���9���b���E�����	�,FC�1"��~	�B�%���l�q����
׿�$	�"�)��N��u�J'���:���ު�,�����/�����Wt�4M���(��!�Rտ�   �   ?�����_������Ծid���;��*��@A���K��چ��3;��Q�ུ�	��^%�Ɂ@�l�X��1l���x�Zx}��y���m�$[��9C��P(������潒)���Q�����N
��r��c>�UZ���־���ha�-��Ϳ�����!�n{C��Bg�1t��N������C���3؟��*���}����f��B�X!����˿�   �   !?�� tN�|���tž�ㄾ�c4�V� �Qvͽr���N,ս`i �:!�U�C��j�^�������bv���d��=�������と��&��Z)���'n�=G�.o"���۽9Mǽ)�ҽ�v��d7������nǾ����O��������|���W���3���R��uq�q��?7������Kv���b��`r�l"S�X3�N��	�g����   �   B�~�o�8���󤲾A.u��R-��9�J������[��V6�u�d�NJ��4Ʃ��ž��޾w�������=�(= ����R���Ǿ�ݫ�2N���h�H�9��b����]��z����/���w�n#������9����̛���ؿ���( ��:�l�S��pi�<Ax�6�}�(�x��kj�V�T�Jm;�2� �H��M�ؿ>���   �   ��\�e7 �c⾓�����_���'�|��Q��V�!�I��b��6آ�X�ɾ�5���X�� 1.���7�d�:��8�G/��!������&h̾�����9���5L�4H$��>����i�)�׃a�\���?Z��� ��]����F������
� "!�H�5��vF� �Q�h;V�B�R���G�x�6��"����`�v���[ ���   �   �[9�!��0p���P��=K��%�օ�L�+�]NS�L}���a����⾕%��/*�8lF�)�_�h�s��7�����k���z�t��6a�++H��+���0K��d��N��C�U��-�]<��~&��L�eՉ�U������k!9��mv�AI���ĿUg�v��,��p%��I.�<�1���.�La&��/�T�����ſ�랿{w��   �   �����ܾm ���\l��c:���&��/�w�S��3��N赾KGﾳ��g�?���f�t��?��*}��i���)��!����\��W��R���;i�)sA��-�:m�|��,Y��sJU�0�0���'���:���l������_ܾI���G�Y����ڟ�_���O�ݿ�����������w�8Z��������Ӳ߿�������|o����H��   �   Ra�&����/���aK��].��/.��J�6���C��������:J���{��m��Oկ��Wſ�Hֿ�@�QD����)w׿��ƿHI��Y���>�}���K�B�Pe�󎰾�1��dK��^.�R/.�T�J�����ȡ��`�쾟��7J���{��k���ү��Tſ�EֿN=Ό@�a�῾s׿��ƿeF��Ӵ����}�{�K����   �   5y���V��dGU���0�b�'���:�l�b���WbܾK�|�G����ݟ��E�ݿ�����������y�2\����/�����߿�������fq����H�*����ܾ�"��t_l�e:���&�ִ/�ܞS��1��D嵾!C������?���f��q��n<��=z��U	���&������Y��ST��Ε���i�oA��*��h��   �   ���|�U���-�;�^~&��L��։�I���?���#9��pv�K��Ŀ�i������r%�$L.�r�1���.�Zc&��1������뿊ſ�ힿ�w�c^9�����r��R���>K� %����B�+�KS��z��P^��)���"��,*�>hF���_���s�35��m���ώ��z�t�C2a�'H�x�+���lF�a���   �   �1L�EE$�
=�����)��a�����8\�;� �]�q����G����"�
��#!�"�5� yF�X�Q��=V���R���G�n�6�`"�����b�n�������\�%9 �ze����>�_��'�������Ƙ!�LI�H`���Ԣ� �ɾs0������H-.���7�>�:��8�Z/�!��������c̾D����6���   �   �_�2{���������/��w��$��ޢ�8�9�u�������ؿ���R) ���:�J�S��ri��Cx���}���x�Hnj�R�T��n;��� �d���ؿ�?����~��8�-��k����/u�WS-�Q9�<��Q���Y��R6�a�d�G��R©���žj�޾ж�����:� : ���� ��_�Ǿ�٫��J����h��9��   �   `۽JǽB�ҽ�v��d7�n����oǾ����O�e���������X���3���R�Nwq�w��c8��)���ww���c��4r��#S���3�B�<񿧦��@���uN�}��2vžL䄾Vd4�T� �uͽ���f(ս�f ����C���j�@�������r���`��������}���"��&��""n��G�ak"�Ć��   �   �N�����		��*��5c>��Z����־���ia�����ͿX��|�!�0|C��Cg��t��������2���ٟ��+���~����f���B�!���p�˿������_�s��ŒԾe��p;�+���@��J��w����7�������	�0[%��}@��X�	-l���x�7s}�αy���m��[��5C�sM(��������%���   �   �a���D��Y���	�FC�@"���	�l�%��l�����׿�$	�f�)�N� u��'��b;��Nߪ�������*0��<���Wt��M��(�R"��Rտ�F���zj��$�a޾����۬?�\�������~�������w���X���ѽ��������%�?�4�t>��B�,??��36�'�'��f�f� �n9׽���7���   �   ����o��������	�p*R�������H�3�]��Dͯ�
���(R8�P\a�i[���F������|��y���C�����+�������}`�s7��W����Fή���~��n2�H��*���P���Bp���Q�����FU���Ĩ��̽E��ħ�� ���.���7��?;�`8��/�ݯ!�����'����Ͻ�ҫ��b���   �   �9��,���t���
��RP�O�g�ﾰ�0��|�����������>5�H4]����4͚������պ�T��-ں�&��������L���v\�
y4���S����Ҝz�*�/�+�����8N��?��1��Fs��0&��Q����9��H��2.��K��2���A�|�K�t�O��`L��B��B3�խ���	���潡[���֟��   �   ��~��$ͽp�
�E*K��И��!�vk(�@&p�����EڿT�hq,��sQ��y����%������cͲ�ѥ��������jey��	Q���+�B�
��ٿ�4����n��v'�(��ס��5I�����ɽ�d��LǮ�J�Ƚ������2���N��uh���|��	���i��TP��?�}�/�i�VP�L�3�c��T���/̽�   �   :����ս�F⽪����C�����ؤԾ6��̎]��U��ޔɿړ ����?�8�b����������֟��B��<���	߂���b�^�?�J��M �5 ɿi͗�(�\�m��WjӾ��$B��t<߽�ҽa��n�
�*�+��YR���{��S��旤��������俾༾�ó�t���N��U�}��ZT�ft-�����   �   X��	��ލ��9���;�J=��X$��2[��E��5��^���(��&`���*�:�G�d��H|��{��F������}���d�P|H��"+�Fu�f��W��뇿9fE���
�08��vm��1`:���� ��!�M��9D���u�^����⵾�ӾQ�����q�P��3�duﾙ�Ծs-��l���7�w�e.F��   �   t�Y���/�E9����P5�$�p�������:s+���k�q���z~ȿ����� ,��TB��U�$�a��uf�><b���U�:$C�*�,�����$��ҹȿ������k��.+���<��3�o�S#4�������-�VX�����*����PؾD-���]�*�0(:�;D��G��VD�p�:���+��������پHد��׊��   �   �D��]Ad���9��((�
	2�}�Z��1��"�; �i�E��}���Ĩ��п������Z@"��0��C:��=��:��W1�6#��0�q���l�ѿC3������r�E����;�ᒾ��Y��/1�",'��g8�D�b�M����������6��$T���n�6 ���̈�~8�����dl����o��JU��'7��Xh��?���   �   ��þ������c�T*=�W�3���G���|���Ä뾒� �̏U�F`������MA̿�r�Jw�8���$����$t��O�4�����CͿiF��)㉿�2V�V� ���G��u�|�|�G�m3��u<�4�b��풾Y�¾� �@�$���L���v�P����b���`��y_�������������,���X��Ax�l#N��l%��� ��   �   �X��#p������vY��:���:��Y�:ċ�ڻ��h��[�'�&X�R������������Iҿ�2����5���3�h��Eӿ?}���z��4��]*Y�I�(��T��xm����uY���:���:�QY�<Ƌ�"ݻ�m��>�'��)X�����2��������Lҿ_6������7���/Iӿ.���}��;6���-Y��(��   �   {� ���7����|�=�G��3��s<���b�a뒾��¾$ �~$���L���v������_���]��'\��7���Ѱ������I��,V���<x��N��i%��� �M�þ������c��(=�N�3��G�x�|�P���9���� ��U�Qb�����9D̿!v�(y�>���&���@v��Q�����FͿ�H��剿|5V��   �   ��E���	�;%㒾��Y��/1��*'�+e8�.�b�3J���������n�A6�d T���n����� ʈ��5������i����o�yFU�$7�x��c��c;��(B���=d���9��'(�Z	2��Z��3����;���E�����ƨ���п)���r��`B"�0�0�&F:���=�J�:�Z1�(#��2�I���˕ѿ25������   �   Ӭk��0+���|��]�o�c#4��������-��X�����7����KؾK*����|�*��#:���C���G��RD�M�:�-�+�*��� ���پ�ԯ��Ԋ�Z�Y�ƃ/��7�A���P5���p�����5��!u+���k�%�����ȿ�������,��VB�U���a��xf��>b�,�U�H&C��,�"��1'����ȿ�����   �   쇿�gE���
�[9��n��h`:�s��r ������z4D���u�����޵�֞ӾHK��O��%���0��oﾪ�Ծ<)��������w�0*F�S�� ��Č�P9�c�;�8>���%��t\���E�7��󖴿!��^a�(�*��G�Jd�FK|��|������s����}�
�d��}H�6$+�Tv���jX���   �   5Η�N�\�4��KkӾ���`B���c:߽��ҽ���8�
��+��TR���{�sP�������������E࿾�ۼ�����Bp��{K����}�VT��p-���� ��:�սgE⽫��[�C�����J�ԾR��`�]�W��9�ɿ�� ���^�?��b�����������yן��C��c����߂��b���?�*���M �Bɿ�   �   95��Z�n�vw'�Ƥ�%����5I�|����ɽsb��.Į�*�ȽO��|���2�[�N��ph���|�����f���M���}�q�i��QP���3�b��BO��P,̽q걽
}��Q#ͽ��
��*K��ј��"�Sl(�w'p�R���Oڿ��:r,��tQ�P�y�e�����!���lβ�̦��a����	���fy��
Q���+���
�cٿ�   �   ���z�Y�/�G+�+����8N��?��0��r���$��5����6�� ��T,��I�m2�m�A���K�ǎO��]L�q�B��@3�׫��	�ӱ�fY���ԟ��8�������s��!
�SP���%��<�0�[|�~�����L��
?5��4]������͚�$���ֺ��T���ں����������L��8w\�Ry4�:�ET��   �   #ή���~��n2��������P�x��o���Q��؂��U��xĨ���̽�D������ ���.���7��?;�`8��/��!�����'����Ͻ�ҫ��b�����Bo��躽���	��*R���?��x�3�}��iͯ�7���DR8�n\a�{[��	G���������{���=������������}`��r7��W�����   �   m���z���/�K*����7N��>�0���q��F$������6����T,��I�m2�r�A���K�̎O��]L�r�B��@3�֫��	�ű�DY���ԟ�D8�����;s���
�CRP�!�'�ﾀ�0�Q|������俶��D>5��3]�ԕ���̚�!����Ժ�~S���ٺ����"���EL��6v\��x4���aS��   �   �3��f�n�v'���렗�4I�{��X�ɽ�a���î���Ƚ%��p���2�^�N��ph���|� ���f���M���}�s�i��QP���3�U��O���+̽�鱽2|��"ͽ��
�])K�CИ�� ��j(�}%p������ڿ�
��p,��rQ�̗y�� ��C������\̲�̤��������dy��Q�2�+���
��ٿ�   �   `̗���\�K���hӾ�}��0	B�1��8߽��ҽ���
���+�uTR���{�uP�������������K࿾�ۼ�����Cp��xK��|�}�VT�sp-�|��C���ս�C�?��#�C�䁏���Ծd����]�-U��Гɿ,� �����?���b���������u���ԟ�GA������݂���b��?�B��4L ���ȿ�   �   �釿fdE�v�
�I6��l���]:����d ������C4D���u�����޵�ڞӾPK��T��*���0��oﾦ�Ծ7)��鸘���w��)F���P������7���;�,<���"��(Z���E��4�����}��_�T�*���G��d�0F|�(z��ԉ��������|���d�|zH�j!+�t�u�濌U���   �   �k�
-+���,�� �o�� 4�K�����8�-�gX����(����KؾJ*������*�$:���C���G��RD�P�:�,�+�(��� ���پyԯ��Ԋ���Y��/�|6�g���M5���p�`���C��q+���k������|ȿ�����
�6�+��RB�@U���a�sf��9b�R�U�"C�V�,�0��W"����ȿѫ���   �   ��E�� �;�ߒ�y�Y��,1��('�d8�}�b�J������{��j�A6�f T���n�����ʈ��5������i����o�xFU�$7�r�wc��?;���A��=d�c�9�&(�t2��~Z�-0����;U��E�L|���¨���пG����n>"�ʪ0�hA:���=���:��U1�2 #�4/�f���אѿ#1��ೃ��   �   �� �r�뾔��S�|��G�*3� r<���b�뒾��¾ �~$���L���v������_���]��*\��;���԰������J��+V���<x��N��i%�p� ��þ(�����c�4'=���3���G�%�|��񪾍��`� ��U�i^��Q����>̿�o쿄u�D���"����r��M�Z�/��AͿ�C��ቿX/V��   �   RP��)j�����4qY�:�:�6�:�gY��Ë��ٻ��h��R�'�
&X�R������������Iҿ�2����9���3�j��Eӿ?}���z��4��V*Y�<�(��T��+m�����sY��:�Ǌ:��Y��,׻��d����'��"X�7�������}��OFҿ7/�A��i��#0���俆Bӿ2z���w���1���&Y�_�(��   �   ��þ����_�c�h%=�
�3���G�S�|��󪾈�뾃� �ďU�C`������MA̿�r�Lw�:���$����&t��O�4�����CͿgF��%㉿�2V�C� ��������|�N�G�3��p<�
�b��蒾S�¾� �*{$�B�L�t�v�����\���Z���X��卻�������S��S���7x��N�jf%�� ��   �   ?��9d�ϓ9��$(�H2��Z�c1����;��^�E��}���Ĩ��п������Z@"���0��C:��=��:��W1�8#��0�q���k�ѿB3������f�E�����;]ᒾ	�Y��,1�('��a8��b�dG���������m
��6�)T���n�����Eǈ��2��&��g���o�BU�; 7�D��a^��Y7���   �   n�Y��/��4�}���M5���p�����Z��+s+���k�p���y~ȿ���
�� ,��TB��U�(�a��uf�B<b���U�:$C�*�,�����$��ѹȿ~�����k��.+������ďo�!4�ĩ�����-�\
X�����~~���Fؾx'�Z����*��:���C�&|G�*ND�!�:�R�+��������پ�Я��ъ��   �   ������@���6���;��<��$��[���E��5��^���)��&`���*�:�G�d��H|��{��G������}���d�P|H��"+�Fu�f��W��뇿,fE���
��7���l���^:����M ������$0D�V�u�L|��hڵ���Ӿ�E��"��������,�"jﾙ�Ծ�$��N�����w�r%F��   �   �����ս�A�ڨ�^�C�`�����Ծ)��ǎ]��U��ޔɿۓ ����?�:�b���������֟��B��<���	߂���b�^�?�J��M �5 ɿh͗�"�\�^�� jӾ�~���	B�4�D7߽��ҽǁ�*�
�;�+��OR�+�{�!M��8���n��H}���ۿ�D׼�V���bl��H����}�QT�jl-�T���   �   �汽z��� ͽD�
�})K��И��!�nk(�=&p�����FڿT�jq,��sQ��y����%������cͲ�Х��~������ley��	Q���+�B�
��ٿ�4����n��v'��㾚����4I������ɽ`��(���T�Ƚ�����t�1�H�N�Rlh���|�R�� d���J����}���i��MP��3�6���I���'̽�   �   �6��錙�tr��[
�2RP�2�V�ﾬ�0��|����������>5�F4]����4͚������պ�	T��-ں�&��������L���v\�
y4���S����Ҝz�'�/�+�����G8N�,?��/��q��,#��u����4��l�㽲*��G�G2��A�]�K�;�O�c[L� �B�t>3�ȩ��	�����V���ҟ��   �   `狽1���vĽ�l��X� 륾������8��Ѓ�д���4W�H�=��+i�Z������������E������tD������s��z���H�h�R�=�v�{;�+���ʖ����8��P������VX�N��#�ý.0����@"���?��B@ֽ���DY�h�&�R5�?f>���A��>��[5���&�d��OA ��׽��������   �   �Ֆ�a��KȽH��%�V�>���/���5���������"�������:���d�r���+T������0�����������m���H�������d�܏:�̼���꿟�������O�5�W����Z��m&V�4
�p^ǽ��������綠�;Ľ�����v$�W�8��H�e�R���V�(S�h�H�Y9��$�Y9����#!Ž�ѥ��   �   �`��-䵽�NԽ7;��|Q�)t���	�2y-�Dw�]©�!<࿶��1��X����=������)��Q���S2��׭��)
�������iX��1�����߿ч��f�v�b1-���뾾���P����DhӽX���z��4aҽS������V�8��jV�Q�p��ӂ�K���������������/q�{�V��h9�lf�O���;Pӽ�   �   0��Tݽ�
꽴K�(�I��꓾�۾zF ��;d�uٜ�HuϿ U��#��BF�pk�"݇��ۗ��ʢ������٢���4���~k��AF�z�#�"@�IϿ����c�7 ���ھG����sI����E-齛qܽ-�����^2��SZ��������zN��e1��4�¾6ƾ�¾�b�������җ�:܂���Z��2��I��   �   �$�^-������-�A�M]��gƾ��nL�\Y�������~�,��>S0���N�ܚl��!������������?����l�>O��k0�Ȼ�x�^칿�C����K�_����ž�!���oA����V�L��YI$��K���~�����Q����ھ~p����`�t���.�y<������^۾���[Y������ZL��   �   �`��)5�dE�^��!5;��jx�_��]I���0��0s�!{��T�ο�4��ε���1�HI���\�8j���n��9j�$�\��TI���1�����a����ο2���&s�k�0���hծ��x���:�!�������4�#)`����^�����߾������0��L@�gYJ�l�M�WsJ�|@��0�8�$��_�.$������   �   �Η��tk��?���-�3�7���a�>񗾵~ԾX���L��������d׿�� �����'���6�lu@�Z�C�z�@���6��'��U�2� ���׿�9��o���L�;��6qԾ|ۗ�Lma�{�7��p-��E?�2k�M���J�ľ�F��9E��D<�)F[���v��5���"������S5��BW��vw�q�[�t�<���^����ž�   �   ��ɾ�C���$k�&oC�F�9�m�N����������E��%�\�\��Ս�� ����ҿ��
��N���������Vy�����U���ӿ�=��1���<�\�U&�Zc�С�������N��k9�:C�0�j�����oɾ�l��*���S���O�����,���/B��/��.���Ԧ�����܈�{AT�Ae*�Z���   �   3�mc¾"����`�@A��A��`�H����2¾K��6�-��Z_�t�>⦿�����ؿ�P뿓���)���6��}���Cٿ�����'���+�� �_�p�-�6��`¾b����`��A��A�N�`�W����5¾���0�-��^_�����妿������ؿ?T�}���-��h:��)��UGٿ����%*���-����_�&�-��   �   �&�rf�ң��������N�kk9�68C���j��
���kɾj��*���S�(�ML������괿<���>���+������Ѧ�����I���=T�9b*�	��4�ɾ\A���!k��mC�:�9���N�%��� ����I�3�%���\��׍�e����ҿ������0P����:�����b{����!Y���ӿ�?����:�\��   �   \L�߹�_sԾ�ܗ�]na�L�7�Mo-��B?���j�L���9�ľAA���A��@<��A[���v�3���������{2���T��w��[���<����l���	ž�˗��pk��?���-���7�F�a���P�ԾF��D
L�����C��Og׿{� ���،'���6��w@���C���@��6�"�'�FW��� ��׿�;�������   �   2)s��0�: ���֮�x���:�'��z��O�4�|$`�����J�����߾���<���0��H@��TJ���M��nJ��w@��0���3��8Z�X �������`��&5��C�����5;��lx���L����0��3s��|����ο;7��h����1��I�R�\�j���n�~<j���\��VI�f�1�.���c��m�ο�����   �   �D��P�K�]����ž�"���oA����}�ڸ��E$�f�K���~�����L��B�ھ�j�������o+�R9� ����Y۾ï���U�����VL���$�F+��������A�@^��ƾe��IL��Z���������l���T0���N�<�l�7#��a���G��7���@����l�O��l0����y���   �   䱜�L�c� ���ھȠ��tI�W��*+�*nܽ@������Z2��NZ�ꋂ�����lJ���,����¾�ƾ~�¾�^�����qϗ�>ق��Z�#�2��F�ݿ�BQݽk	꽴K���I��듾!۾�G �X=d��ڜ��vϿ V�(�#��CF�@k�Aއ�ݗ�7̢����Yۢ�F��9��k��BF�d�#��@�/JϿ�   �   [���/�v��1-�>����+�P�G���fӽ
 ���w���\ҽ�������m�8�JfV�L�p��Ђ�r���ދ�2���=����*q�)�V��d9�Uc�g���sLӽ6^��x⵽,NԽV;�W}Q��t���
�z-�GEw�/é�.=�^��1�2�X�ҋ��"������*��e���Z3��Ů���
��%����jX���1� ����߿�   �   ״�������5������Z��`&V��	��]ǽ�~��!�����9Ľ�������t$��8�J�H���R���V�xS���H�	9��$��7�ˉ��ŽХ�~Ԗ�R`���JȽz����V����������5�丁�������<��8�:���d�Ὁ��T��E�������O���j���熵��H��������d�(�:������   �   �������ϑ8��P��N���X���ɇý�/���
���!��e?���?ֽ����&Y�M�&�:5�+f>�~�A��>��[5���&�j��VA ��׽��������狽p��*wĽ�l�h�X�X륾�����8��Ѓ�,д����NW�f�=��+i�m�����������E������nD������d��i���(�h�6�=�^�S;��   �   !���8�����5�����TZ���%V�h	��\ǽ+~��������9Ľ�������t$��8�Q�H���R���V�|S���H�9��$��7���Ž�ϥ�8Ԗ��_��2JȽ�����V���������5�\���S�����꿤��l�:�h�d�&����S��9�������.���O���܅���G��D���t�d�\�:�j�����   �    ���+�v�{0-�M�������P�<���eӽ5���:w���\ҽΗ�����j�8�KfV�R�p��Ђ�w���ދ�7���@����*q�)�V��d9�Kc�2���"Lӽ�]���ᵽ�LԽJ:��{Q��s���쾦x-�?Cw�����j;�<�n�1�4�X�����v��!����(��@���B1��լ��F	��Ղ���hX�>�1� ��	�߿�   �    ���}�c�
 ���ھ����qI����S)�mܽ�����|Z2�vNZ�苂�����pJ��-����¾�ƾ��¾�^�����pϗ�:ق���Z��2��F�"��Pݽ��AJ���I��链e۾�E ��:d��؜�5tϿnT�&�#�RAF��k�܇��ڗ�tɢ�4����آ�������k�<@F�f�#�F?��GϿ�   �   �B����K�����ž� ��mA�Z���|�0��tE$�'�K���~������L��D�ھ�j����	���t+�V9�����Y۾�����U��Ј�IVL�v�$��*�~����8�A�(\���ƾ	���L�WX�������|����Q0�(�N���l�� ��g��3��> ��5>��,�l�RO�
j0����v��깿�   �   <$s�l�0�(��JӮ��x���:�H��M����4�$`�׻��8�����߾���>���0��H@��TJ���M��nJ��w@��0���0��-Z�D �����8�`�'&5��B�����2;�-hx������F��U�0��.s��y��k�ο92��Z���1�"I�6�\�tj���n��6j���\�FRI���1�"���^��Y�οv}���   �   XL�;��LnԾSٗ��ia�W�7�dm-��A?�F�j�����ľ/A���A��@<��A[���v�"3���������~2���T���w��[���<���[����ž�˗�pk���?�ö-���7���a�m;|Ծ���?L�i�����9b׿r� ����'�V�6��r@���C���@�h�6��'��S��� ��׿}7�������   �   ��%��_�
���f���`�N��h9�k6C���j��
���kɾj��*���S�'�NL������괿@���>���+������Ѧ�����H���=T�0b*������ɾA��� k��kC�h�9�p�N�枂�7����B�q�%�\�\��Ӎ�}�����ҿ���4��L�z���}�t��Bw���nR���ӿ�:������\��   �   ��H]¾מ���`�XA�lA�K�`�ȅ��O2¾6��,�-��Z_�t�?⦿�����ؿ�P뿘���)���6������Cٿ�����'���+����_�f�-� �``¾ࠐ�j�`�CA��A�t�`�����/¾>��}�-�NW_�H򊿨ߦ�������ؿ�L�����%���2��Ǎ뿁@ٿb����$��A)��2�_�r�-��   �   M�ɾn>��rk�jC��9�9�N����2����E��%�S�\��Ս�� ����ҿ��
��N���������Xy�����U���ӿ=��0���3�\�D&�c�d���ѝ����N��h9�	5C���j�T��Qhɾ�g��*���S����I������紿���Q;��O(������Φ�3������9T��^*�z���   �   �ȗ��kk��?�d�-�a�7�Ǡa���`~ԾB���L��������d׿�� �����'���6�nu@�\�C�|�@���6� �'��U�4� ���׿�9��m����L�#���pԾ�ڗ�vka���7�wl-�i??���j�e~��d�ľJ<���>�=<�:=[���v�t0����΄���/���Q��qw�}�[���<��������ž�   �   ��`��"5��@�����2;�eix�� ��I����0��0s� {��S�ο�4��ε���1�HI���\�:j���n��9j�&�\��TI���1�����a����ο1���&s�Z�0�����Ԯ�Vx�f�:�������̯4��`�����o�����߾�����;�0�LD@�lPJ�K�M�\jJ�|s@�"�0�8�$��U�;��|���   �   �$�6(���F�r�A��\��ƾ��eL�[Y�������~�,��@S0���N�ޚl��!������������?����l�@O��k0�ʻ�x�]칿�C����K�I��O�žn!���mA�"���{�&��aB$��K��~�v���OH��;�ھ�d��l������ (�*6�+���ST۾H���	R��؂��QL��   �   L��Lݽ���I���I�x꓾_۾kF ��;d�tٜ�JuϿ"U��#��BF�pk�#݇��ۗ��ʢ������٢���5����k��AF�|�#�"@�IϿ����c�( �]�ھ埓��rI�����'�;jܽH�����V2��IZ����������F���(���¾�ƾ��¾@Z������˗�(ւ���Z���2��C��   �   �Z��rߵ�xKԽ:��{Q��s��k	�,y-�Dw�\©�"<࿶��1��X����=������)��S���S2��׭��*
�������iX��1�����߿χ��c�v�X1-�v�뾀��<�P�^���dӽ�����t��Yҽ	��������8�bV���p�B΂�����Kۋ�l�����&q���V�a9�`�����Hӽ�   �   �Җ��^��hIȽ�����V�!������5���������!�������:���d�s���*T������0�����������m���H�������d�܏:�̼���꿟�������L�5�I����Z��&V��	��\ǽ�}�����뤽�6Ľݡ����r$���8��H��R�X�V��S�^�H��	9���$��5����&Ž�ͥ��   �   ޗ��+�����ý^����W�40������8�*��M곿�n�z���=��g����D!���˸�N^������`��rظ��>������]h��l=������cb��ڄ���8��o���ȥ�G�X�{���8ŽV̌�Zܗ�g貽t�׽�� ����#'��s5�Α>��A��b>��5�ۭ&��g�������ֽ����W����   �   �z��S�����ǽ��^�U�T�����n5�\��4���鿘9�l�9�\�c�<��뉠�x���k��6���� ���������~0��p	d�Z@:�V���[�Ᏹ�{m��֛5����������V�����	ɽ�9��沗�8�����Ž,｣w��%��'9���H�LS�m�V�9�R�'�H�Ϫ8��v$�������ƜĽ�h���   �   r䷽Wm����ӽ���f�P��Ϝ��뾔�,�7!v�1���;߿�k��0�ؘW������_��#���]��j���R��5ܨ��]��?���W��-1� ��Q�߿�X����v�� -����.V��y�Q��|�ս�����&��YԽJ �r����9���V��q��傾�������b��|���H�p��=V���8���q�����ҽ�   �   ��#�ܽ�o�'���HI�_���?ھʛ��Fc�?4��9�ο����D#���E�6j�[c���K��!�����P���+���H�� j�6�E�f^#����(�ο�u���c�G��u�ھ�ѓ��J�����V�ݽK`�\��^3�H�Z��΂�����_���!���¾K�žm¾�ڸ�� ���H���`���Z��I2�_���   �   �B$�`��d����QA��Pež�"�dPK�ً�^��?��6K�D�/�p]N���k������n��G|��hS��˒����k�8N�Ⱦ/�vC�^���}������t�K��a���ž�J����A��=�,�Fl���$�lL�2z�q8���y���	۾FZ���������:������������|ھ�뻾.���h�~�(�K��   �   ��_�O�4��������:�b�w�����h���`L0�Pxr��	��"ο����n��]1��H��=\�(`i�2�m��)i���[�SH��1�t7�n��9ο����r�o0�����,ˮ��Rx�_M;�-*��s��G5�U�`�$����﴾6	���\��%�0�
@�0�I�xPM�`�I�s�?�*0��o��V�l`߾�_��6����   �   �E��.�j��2?�Po-���7�HAa������Ծ�]���K�Eb������׿� �����O'�p36�x�?�LSC���?�x�5���&����nW ��ֿE���|K��ԀK�|b��!Ծ|ɗ�ĕa��8���-�.�?��dk������ľ�S���A�}3<�� [�?�v�� ��.֌�S%��'���YЅ�C
v�h�Z�`�;������uAľ�   �   �ɾ�ӗ�æj��,C��h9�jN�K~��0[��P�򾝟%��4\������ʯ���ҿ^��V��N�
���tZ�>��\6�A)�ҿu���i����[�@z%���S��;�����N��9�TvC��k�/���oɾdc��	*�|�S���~��/��j�����8�����������`����!ؓ�KP~�JCS�ͣ)����   �   ������8[��|y`�
A��A�{�`�R{���¾&���[-��$_�Պ�m���*]����ؿz�꿚���%o���Q��ؓ�Dؿ���[������v�^��-��������xY���w`��A��A�ޛ`�`}���¾Z���^-�(_�k׊�/���O`���ؿ7�꿀���s���U��~��]Gؿ����]��&�����^�t-��   �   v|%�)��U��\���Q�N���9�vtC�`
k�����kɾ�`��*�u�S���~��,���f��͡��ϧ��v���\���U]����}Փ��K~��?S�Ƞ)�@�dɾ@ї��j�p+C��h9���N�����]������%�#8\�Ӥ��4ͯ���ҿϹ�B��f�>��$��\�H��48��,�kҿrw���k����[��   �   (�K�"d��#Ծ�ʗ�ؖa�~8�F�-�~�?��`k������ľjN���>��/<�?[�'�v�:���Rӌ�o"��R����ͅ�Rv��Z���;���������=ľ�B��z�j��0?�^n-��7��Ba�2���=Ծ�_�2�K�d��ĭ��׿�� ����R'��56���?��UC��?���5���&�N���X �^�ֿ?���	M���   �   b�r��p0�����y̮��Sx�sM;�5)��q��D5���`�����봾�ް����$~0��@���I��KM���I�7�?�&0�(l��S��[߾�[��P�����_�z�4�������:�8�w�A������RN0��zr�^��M!ο;����o��_1�2�H�d@\��bi��m�^,i��[�BUH�|1��8�wp��$	οu
���   �   �����K��b��žAK���A�4=��*��i��$�qgL�(t��4��Fu���۾^T��p��,���7�n�����8����wھ�绾����Ņ~�ݗK��?$�J��@��Ԧ��QA���fž2$�;RK�Qڋ��_��@��rL���/�^_N�@�k����>p���}���T�����ʩk�� N�,�/��D���U���   �   pv��C�c���t�ھzғ��J����ʫ���ݽ`[���(3��Z��˂����
[�����n�¾��ž�h¾7ָ������E���]���Z��E2�b���	�L�ܽtn�&���II��_��Aھ��[Hc�Q5����ο����E#��E��7j�vd���L��u"��%�����0-���I���j�l�E�R_#�8��A�ο�   �   kY��z�v�!-�?�뾂V����Q��|��ս@���x#�� �ӽ� �,����9�8�V��q��₾�}������_��֫��j�p�y9V��8���������ҽ�᷽�k��ʷӽ����P��М���v�,�s"v����&<߿ll���0��W�g����`��%���^��|���S��#ݨ��^����� �W��.1�����߿�   �   ����m���5�D��������V�p��%	ɽX8��/������@�Ž�(ｶu��%�`%9�K�H��S��~V���R���H���8��t$�������x�Ľ�f���y��������ǽ���U���������5�����������9���9��c����n���	������Ǜ��L������s����0���	d��@:�����[��   �   ?b��������8�Oo���ȥ� �X�D��s8Ž�̌�ܗ�-貽.�׽q� �����#'��s5���>��A��b>��5�ڭ&��g������ֽ����|������b�����ý�����W�i0��O����8�/*��s곿 o����=�"�g����W!���˸�U^������`��hظ�|>������]h��l=�������   �   e���m��F�5�>���e����V����mɽ�7��갗�ߡ��(�Ž�(ｴu��%�b%9�O�H��S��~V���R���H���8��t$�������^�Ľ�f��Ry��3���Դǽ���U�"������=5�8�������d9�$�9���c������������������1 ��������0���d��?:���[��   �   X��t�v��-�N��=U����Q��{�Cսj����"����ӽ� �����9�7�V��q�ゾ�}������_��ګ��m�p�x9V��8����a�����ҽ?᷽�j��y�ӽ���x�P�VϜ�� ��,�q v�����e:߿Lk�z�0���W����6_��9���\��Z���	Q��3ۨ��\������W�-1�z��K�߿�   �   �t��t�c�����ھ�Г��J����꽼�ݽ�Z�؃�3��Z��˂����[�����t�¾��ž�h¾<ָ������E���]���Z��E2�.����&�ܽ�l齶���GI�3^��p>ھ���Ec�p3��(�ο���C#�z�E�~4j�Yb��_J�����P���	���*���G��8j�ԖE�R]#������ο�   �   ������K��`���ž,I��`�A�x;��)�+i���$�/gL�t��4��@u���۾dT��s��0���7�s�����<����wھ�绾������~���K�[?$����+����$OA��퇾�cž�!��NK�؋��\�����"J���/��[N���k�e���Jm���z���Q��m���>�k�NN�>�/�:B�_��`|���   �   n�r�m0�����ɮ�FOx��J;�T'��p��C5�<�`������봾�۰����(~0��@���I��KM���I�:�?�"&0�*l��S��[߾�[��/���F�_���4����,����:���w�؁������J0�	vr�$��<ο?����l��[1�ʰH�P;\�f]i�T�m��&i���[��PH��1��5�wk��ο7���   �   &~K��`��ԾTǗ�O�a���7�]�-�L�?��_k�թ����ľVN���>��/<�?[�+�v�;���Tӌ�q"��T����ͅ�Vv��Z���;��������=ľ�B����j�`/?�{l-���7�`>a�ȡ��/Ծ\�3�K��`��쿭��
׿�� �>���M'�016��?��PC� �?�&�5���&�Ĝ��U �K�ֿ����I���   �   �w%�Q���P�� ����N���9��rC�=	k�=���kɾ�`��*�q�S���~��,���f��ϡ��ҧ��y���_���V]����Փ��K~�~?S���)�4�2ɾ�З�Ƣj��)C�f9�p|N�||���X����\�%��1\�Ѡ��Lȯ�+�ҿ!��~�J��|���FX�.��v4��%�ҿ�r���g��o�[��   �   ��������V���s`�$A�A�ܗ`��z��?¾���[-��$_�Պ�m���+]����ؿ}�꿞���*o���Q��ۓ�Dؿ���[������p�^��-��������X��v`�A��A��`�y���¾���X-�2!_��Ҋ�ֻ��/Z��>�ؿ���ǃ��?k���M��&�꿑@ؿ����[X��������^��-��   �   ��ȾWΗ�l�j��'C��e9�3}N��}���Z���򾌟%��4\������ʯ���ҿ_��V��P����xZ�@��^6�D)�ҿu���i����[�0z%����*S������R�N���9�HqC�ik����Qhɾ�^��*���S�f�~�_*��d������y�������}��Z��	���ғ��F~��;S���)����   �   �?����j��,?�k-�ǣ7�o?a����PԾ�]��K�Ab������׿� �����O'�r36�z�?�NSC���?�z�5���&����pW ��ֿE���zK��ʀK�gb�+!Ծ�ȗ��a���7�t�-��?�N\k�&����ľrI��l;��+<��[�B{v������Ќ��������ʅ�L v���Z���;���������9ľ�   �   ��_���4����;����:���w����'���PL0�Hxr��	�� ο����n��]1��H��=\�*`i�4�m��)i���[�SH��1�v7�n��:ο����r��n0�����ʮ�Qx�K;��&�o�A5��`� ����紾L�߾��a��Lz0�y@�:�I�_GM�n�I��?�/"0��h��P��V߾�W�����   �   �;$�B�����~��\OA�N�dž�"�XPK�ً�^��>��6K�B�/�r]N���k������n��G|��iS��̒����k�:N�ʾ/�xC�`���}������k�K��a���žJ���A�D;�l(�"g���$��bL�qn�$1���p����ھ�N��W�����54�#��}��m���irھ-㻾櫜��~��K��   �   ��ӷܽ�j�N���GI��^��g?ھ����Fc�>4��9�ο����D#���E�6j�Zc���K��!�����P���+���H��j�8�E�h^#����(�ο�u���c�9��>�ھ�ѓ�`J��������ݽgV���-
3�,�Z��Ȃ�����*W��`����¾�ž	d¾�Ѹ������A���Z���Z�kA2�����   �   %޷��h���ӽt����P��Ϝ�f뾌�,�5!v�1���;߿�k��0�ؘW������_��$���]��j���R��6ܨ��]��?���W��-1�"��T�߿�X����v�� -�w���U����Q��{�� սȧ��X ��-�ӽ  �"���9��V��q�g����z��E���]��3�����p�5V�6�8����5�����ҽ�   �   �w������ǽR���U�5�����j5�\��4���鿘9�n�9�\�c�<��뉠�x���i��7���� ���������}0��p	d�\@:�V���[�㏱�zm��ӛ5�����ޙ����V���LɽG7��Я��A�����Ž�%�t��%�+#9���H�S�|V���R� �H�1�8��r$�������ΗĽ�d���   �   `���U;�����s�ڧO�����P3�_1��r|��A��;��x����5���]�SN������t���|��L��2���p���^/��J���$�^��6�n���1濲b��-~��S2��-򾭄���R�j�
�ұ��4Ô�����x����ﭽ�ѽ<�����"��/��8��S;�Z8�
�.��� ����W��Dνz|���E���   �   ���cM��䭿�^���M��Ꜿ����<.�yx������H�B��*�2�RZ���������7����L������+H��ĝ���Ę�����B�Z�N�3�����񢫿�z��|/����f���IP�&�
�cý�ӛ���������O��_O�
I
�6 ��x3�z�B��PL�~rO���K�q�A��$2�!�������TƼ�Ë���   �   �l��v���\˽
V	�u�H�Z����/�-&�H�l��Ģ��(׿�C	��D*���N��sv��,�������D��b[��)���g��>&��>�v��IO���*�d�	��4ؿţ��8On��D'�]��ZT��P,K�mI�0�ν���R���&ν��������3�zGP���i�X]}������	��ު��8|�f�g��}N�d2�s����Xʽ�   �   ����%Խ@u��p���A���~%Ҿ����Z��~���<ǿJP���Z�D�=��u`� M�����G3������C ��Vӏ����;`��>�̕�������ǿy����[�>��~�Ӿ����C��=���㽱�׽e^콲E���-�iDT��s}��ܒ�/Ҥ�����@����񾾰���}@���ۣ�gÑ�T){�.R���+�FJ��   �   �f���� ��#��J:����.���	�
�C��Ɔ��ɲ�˂俦0�^�)�xF��Kb�z����~Շ��ф��Dy���a�B�E�:)����	����߁D��x
��>��	���b�;���W8�I�� �>8F�4�w�h>�� b���Ӿ��f����x*
�.���� ����OeҾ��l���Lu�hD��   �   ��W��.�}(�����%4�X�n��C����Z�)�R�i��\���ǿ���~6�+��:A��S��_��c��F_�N�R�@W@�NX*���?m��[�ƿ�W����i��9*�=8�����\p�(~5�cT�F����/�F�Y�bz����e�ؾ�9����|*�ge9�j�B�Z�E�HB��8�(�)���K�׾i����>���   �   ����Lb�c8�iU'��B1��qY�ZX��]�̾x��SD�⣂�|˧���Ͽ������"�!�J�/�*�8���;��k8�$�.�Զ �P-�n���ϿuT��Qi��-D�����̾Z���xNZ��:2��r(�۹9���c�^ϒ��[������B�5�8�S�:n�kc���쇿���n���W뀿��l�<lR�6�4�f��|?�?����   �   ���Ja���hb��r<��3���G��#|��M��:t� ����T��ǈ�\ߩ���˿P�������r��j����w�$E��V�uʿ����8����S�|t�[�5���F|��G�ˬ3�#<=�ˀc�i&���¾�����H$�
�L��Tv��2���Π�E���9)�����k˶��ݭ�&����Z��H�t��OK�HE#��]���   �   �����麾#S����X�՛:���:�!9Y�����󅻾���*h'���W�9"���*�����ѿ�o'�������~0�9oпz۹��5���_��TfV�ģ&������溾tQ��(�X�c�:���:�k;Y�����򈻾A���k'�f�W�{$��/-������}�ѿ��2+�񿳨�4�xrп`޹�G8���a���iV�^�&��   �   �v�W��6��I|���G�I�3�W:=��}c��#��`�¾�����E$�&�L�4Pv�90��̠�����%������'ȶ��ڭ�L����W����t�SLK�`B#�/Y�����_���eb�`q<��3�ψG��&|� P���w�e��؏T��Ɉ��᩿��˿��뿜�������l�����x��F�Z��wʿA���:����S��   �   ^/D�\���̾�����OZ��:2��q(�F�9���c�{̒��W�����q�5�έS�Nn��`��#ꇿ �������耿�l�hR���4�i���:�������� Ib��`8�{T'��B1�6sY��Y��ى̾O�0VD������ͧ�P�ϿŜ�����"�!���/���8��;�$n8�J�.��� ��.��p���	Ͽ_V���j���   �   �i� ;*�V:�T����]p�<~5�vS�M����/�ʺY�[w��+��}�ؾ�6�~��0x*�:a9��B���E��zB�Ե8�j�)����BH�w�־�����;��v�W�.��&�i��h&4� o��E�����8�)���i�G^���ǿ2��8��+��<A���S���_���c�*I_���R�HY@� Z*�N���o��7�ƿfY���   �   ��N�D��y
��?��������;�~���6��F�g	 ��3F�b�w��:���]����Ӿ1�c����3'
������ �b��p`Ҿ�촾ݖ��u�?D��b��� ��#��K:����0��Q�	���C��ǆ�i˲�����1�Ԋ)��yF��Mb��z�-���և�"ӄ��Fy�
�a���E�X;)�����[���   �   G���[���t�Ӿ��R�C�X=����Z�׽�Y콂B�~�-�`?T��m}�Oْ�GΤ����������P���X<���ף�����#{�r�Q���+�`G����/#Խ�s��p���A�{��&Ҿ�� �Z����F>ǿ�Q���[���=��w`�'N������4���������yԏ�u���<`�
	>����������ǿ�   �   O����On�E'���㾫T��s,K�$I���νҐ��2��� ν�������3� CP��i�X}�A������)����2|���g��yN��2���[���hTʽAj�����\˽&V	�!�H�����0��-&�v�l�nŢ��)׿:D	�XE*���N�2uv��-�������E��g\��*���h���&��^�v��JO� �*���	�V5ؿ�   �   )���z��|/�A��g���IP��
�4bý�қ������
��M��3L�+G
� ��v3��B�ANL��oO�Y�K� �A��"2�(����2��ļ��������L�����������M�`뜾m��L=.��yx����&Iῢ����2��Z�Z����������5M��<����H��9���CŘ������Z���3�T��i���   �   �b���,~��S2��-�|���yR�4�
�{���������5����ﭽ��ѽ����ʄ��"���/��8��S;�Q8��.��� ����W��Dν�|���E�������;��8����s�#�O�����3�1��r|��A��e�俐����5���]�cN�����t���|��L��,���f���P/��;����^���6�X���1��   �   w���z�%|/�D�]f���HP�c�
��aý9қ������
���L��!L�(G
� ��v3���B�FNL��oO�]�K��A��"2�)����&��ļ�ꉞ�\��FL���������M��Ꜿs�쾔<.��xx�U���DH����2��Z�����E���ǒ��'L��(����G��;���hĘ�c�����Z�֊3��������   �   ����Nn��C'���pS���*K�H���ν����������ͽy�������3� CP��i�"X}�F������.��� 3|���g��yN��2�v�0���"Tʽ�i�����Z˽&U	���H������.�~,&���l�!Ģ�/(׿(C	��C*���N��rv�,��ᅠ��C��_Z��(���f��k%���v��HO���*���	��3ؿ�   �   o��W�[���ތӾl���C��;����2�׽�X�GB�Z�-�L?T�tm}�Lْ�HΤ����������U���]<���ף�����#{�d�Q���+�0G���"Խrཌྷo�z�A�����X$Ҿ��q�Z��}���;ǿ�N��Z�(�=��t`�1L�����2��R�������"ҏ�y��h9`��>������e�ǿ�   �   ����D�Bw
��<�����;�̽��5�F�� �v3F�9�w��:���]����Ӿ4�c����8'
� ���� �h��r`Ҿ�촾�ܖ��u�	D������Ԕ ��!� I:�����-���	���C��ņ��Ȳ�'�俞/��)�bvF��Ib��z�m��ԇ�aЄ� By��a�t�E��8)������|���   �   8�i��7*�r5����lYp�a{5��Q�!��۾/�U�Y�5w����n�ؾ�6�}��2x*�<a9��B���E��zB�׵8�m�)����BH�o�־�����;���W�g.��%�����#4���n�RB�����)�"�i�*[���ǿe ��5�p+��8A�ƒS���_�l�c��C_��R�$U@��V*�d���j��E�ƿBV���   �   �*D�����̾E���!KZ��72��o(��9�1�c�@̒��W������m�5�έS�Pn��`��&ꇿ#�������耿�l�hR���4�g���:����K���pHb��_8��R'�@1��nY��V����̾��_QD�d����ɧ�g�Ͽ���p��:�!�&�/���8�6�;�xi8���.�ش ��+�k��ϿYR���g���   �   r���a2���B|���G���3��8=�h|c��#��+�¾�����E$� �L�0Pv�80�� ̠�����%������+ȶ��ڭ�N����W����t�QLK�ZB#�Y�������^���db��o<�3���G�V |�hK��
q����ĉT��ň�ݩ��˿,�������`��h����u�RC��S�4rʿ�	���6����S��   �   l����㺾O��O�X�
�:�C�:��7Y������������h'���W�7"���*���� �ѿ"�q'���� ��0�=oп}۹��5���_��QfV���&������溾�P����X��:�ܵ:��5Y�_����������e'�X�W�  ��(���ﺿ�ѿ�㿻#�%��B���,��kп|ع�"3���]���bV��&��   �   '���B\���ab��m<�{3�f�G�t"|�MM���s������T��ǈ�Zߩ���˿O�������t��j����w�&E��V�uʿ����8����S�nt�"꾤4���E|���G���3�A7=��yc�_!����¾h����B$�~�L��Kv��-��)ɠ����"��r����Ķ�w׭�d���[U��S�t�xHK�A?#�NT���   �   r���uDb�.]8�XQ'��?1��oY��W���̾_��SD�ޣ��y˧���Ͽ������"�!�H�/�,�8���;��k8�&�.�ֶ �P-�n���ϿuT��Pi��-D���7�̾ж���LZ��72��n(���9���c��ɒ�	T��:������5���S��n�0^��n燿^������"怿*�l��cR�֜4�F���5���   �   ��W�T.��#�����#4���n��C��΁�I�)�K�i��\���ǿ���|6� +��:A��S��_��c��F_�P�R�BW@�NX*���Am��]�ƿ�W����i��9*� 8����2[p��{5�Q����,�/�R�Y�rt��p��Ӫؾ4�2��wt*�*]9���B���E��vB���8���)�]��XE���־О���8���   �   p�s��k� �Z!�4I:�� ��5.����	���C��Ɔ��ɲ�ɂ俤0�^�)�xF��Kb�z����~Շ��ф��Dy���a�D�E�:)��������؁D�}x
�u>�����;�����4�D� �`/F�لw�Y7���Y���Ӿ�
�`�~���#
�в��� ����z[Ҿe贾nٖ�
u���C��   �   @���Խp�(o���A�F�F%Ҿ����Z��~���<ǿIP���Z�F�=��u`�M�����F3������D ��Vӏ����;`��>�̕�������ǿy����[�0��H�ӾB����C��;�g�㽉�׽�T�p?���-��:T��g}��Ւ��ʤ��񲾃񻾠达����78��ԣ������{�~�Q���+�D��   �   �f���
��vY˽�T	���H����w/��,&�D�l��Ģ��(׿�C	��D*���N��sv��,�������D��b[��)���g��?&��>�v��IO���*�f�	��4ؿƣ��5On��D'�>��T���+K�@H���νl���'���7�ͽݽ��� ���3�?P�"{i�S}���"�������-|��g�juN�) 2�d�0���.Pʽ�   �   ���#K��=���Ι���M��Ꜿ����<.�yx������H�B��*�2�RZ���������7����L������+H��ŝ���Ę�����B�Z�P�3� ����򢫿�z��|/����f��hIP���
�_aý�ћ�����	���J��{I轌E
�/ �vt3���B��KL�SmO���K���A�r 2�%��$��-�佈�����   �   snt��3��FX�����VA��򓾟w߾��$�>�j�y���uտ�)��(��M��7t�&ލ����ת�����>ݪ�~>���/���;u�BN� *�4R	��h׿�	��Eim�M�&�l⾝S��{E����쳽�����z�������B����ĽDS�@�����$�n�,��S/�~,��K#���Q�,��,׾�����[���   �   T&���ߋ��ް�&S��s?�z��� ܾ|"��Fg�M���:ҿ�7&�D�I�ҥo�~������������	��c���0��Fup��J��X'�(*��Կar��0�i���#���޾�W��0\C��%��c���2��#m��d�������ڽ���L5��Q(�'z6��Z?��B���>�H�4��&����h���.�ӽC���ȑ��   �   𖢽c����������:�����Ҿٝ��\�ӳ��
�ȿ|# �x��ަ?�F�b�r̂�����S��"���0���ґ��Â��c��@@�t^��� ��9ʿ�阿��^��3�LվH�����>���B½�����騽|e�����0��o�(��OC���Z�(Dm�Q�x�"�|���w��rk��[X�5b@�;�%��y
����B��   �   *u׽AĽ��Ͻ�w��b4�W0���þ��K��C������G���� �0�pxO��m����8u��|���5���O���l�,O��0�P!��f�*޺�Z���:M��E�K�ž0��O�7�/����սbeʽd�ݽ���*
#� G���m������@��$`������$Q����*D�����ч�4�i��jC��x�|9��   �   ��?���ؾ�m���w-�a)t��1���c ��a6��;{��ܦ���տ.��!��f8��6Q�`f�nt��x��vs��e�d4P���7������[�տUB���0|�nW7�H��β�xw��=0����[������4.���9��h�����F���-ƾ:�޾J��O���� ���mB𾌘ܾL�þ{���w���d�`Q6��   �   ��H���!� ��d�R�'��^�z霾r'�>N�	�Y�����������	�,��J�3�f/D���N��|R�MN��C���2��������B�柹��򐿑.Z���C4������a��*��������$��"L�X���~�l�ʾ�q󾣌�t.��-�]�5���8�;@5�_,�����'����Ⱦ֨�����   �   ����R���+�_�2d%�V�J������Ͼ��i��7�J�s�H����U¿��迺�����(�#�D,�v�.�Ԍ+�V�"���������"@��=��� s�c�6��t�,4��b.��_L���&�V���.���U�su��b���(㾦���)�0�E�7S^�?�q���}�Qπ���|�,Bp�,�\���C�^(�+��R�������   �   n���|���@S� �/�XN'��v:���k����ھ�zRF�8l��Þ�'m��=�ܿ����x���F��W������������ڿ�弿���?�}� VE����Jھ>Ꞿ��k�P;��9(��71��U�Ų��v��5ﾍm��?�f��ʅ�#G��{���"��浭����!0���#��������c�45=��������   �   ��꾟L��e��p�J��{.��.�#;K�:���Q>���
��D��2I��z������֮�YĿoԿ��޿Z��u޿+6ӿ��¿CU���M��1mx�h�G��%����'J�������J�7{.���.�C=K����A���쾇G�$6I��z�+����ٮ��Ŀ�rԿ�޿���	޿y9ӿ�¿�W��=P��qx���G�m(��   �   ��eMھ잾��k�;�T9(�M61��U�p���"���ﾢj�[?��f�eȅ�^D��������Ʋ������<-��@!��L�����c��1=�.�����k���z��&>S���/�DN'�x:��k�(��:�ھ@ �tUF�p�ƞ��o��]�ܿ���X���H��Y����^������ڿ{輿������}��XE��   �   ~�6�7v�6���/��`L���&���].��U��r�����$㾱�V�)��E��N^�I�q�d�}��̀���|�Q=p���\���C��(�d����e�U�����R�t�+�}�rd%�� K�읈��Ѿ�^k�,7�n�s�C���YX¿x��\�����0�#�j ,���.��+�L�"����"��.�YB��
���#s��   �   �0Z����86�+����a��*�϶�&���$�\L������죾ٮʾ l�m���*��-�H�5���8�5<5��,�j���$�M��hȾl��������H�V�!�����c���'��^��Ꜿ�)��O�n�Y�^�������m濆�	�ԧ�6�3��1D��N��~R�LON��!C�X�2�4��$��E忤������   �   b2|��X7��H��ϲ��w�)>0����BY��T���+�F�9�nh�G���6���tƾ�z޾���J���� ����<�j�ܾ��þ1w��Ut���d�~M6�A��u���ż�6��Zx-�+t�t3��e ��c6�>{�ަ�i�տF��X"��h8��8Q��f��t�~�x�Pys��e�66P��7�"������տ�C���   �   ���;M��F�1�ž�����7�·���ս7bʽ��ݽ���Z#�KG��m�����!=��1\�������L�����L@������·���i�;fC�_u��6�7q׽�>Ľ^�Ͻ�w��c4�1��i�þ��K��D������Ό����L�0��yO��m����\v��1}���6���P����l�n-O�$�0�""��g�-ߺ��   �   3꘿r�^�R4��վ����Ӌ>�ǹ��@½ޡ���樽�a�����4����(�tKC�<�Z�B?m�0�x���|���w�.nk�dWX�W^@��%�w
�a���캽z���ma���컽���9�:���(�Ҿ����\�������ȿ$ �.��Ƨ?�n�b�(͂�~���dT��	���1��Jӑ�LĂ��c��A@�_�$� ��:ʿ�   �   �r��x�i�	�#��޾�W��&\C��%�c���1���k��f������ڽ;��P3��O(��w6�aX?�%B�9~>���4�y&����5�����ӽ�@��Ǒ�6%���ދ��ް�|S���s?�����!ܾ�"�aGg������:ҿd��7&�̌I���o�����{���n��/���	��ɺ��o0���up�v�J��X'�Z*�/	Կ�   �   �	��im�$�&��k�nS��:E�Q��쳽J����z��q���mB��E�ĽS� ������$�X�,�wS/�s,��K#���R�7��8׾�����[���nt�.4���X�����A�"��w߾��$�w�j��y���uտ�)�,�(�M��7t�4ލ����#ת�����9ݪ�u>���/���;u��AN��*� R	��h׿�   �   �q����i�Z�#�+�޾RW��][C�9%�Vb��;1��Rk��6��a����ڽ4��J3��O(��w6�eX?�)B�;~>��4�{&����6���|�ӽ�@���Ƒ��$���ދ�ް��R���r?�P��� ܾP"�pFg�����9ҿ���6&��I�^�o�/�������|��3�����繛��/���tp���J�2X'��)�UԿ�   �   �蘿��^�3�!վk���Q�>�ʸ�v?½���o樽Ga��p��"����(�nKC�=�Z�G?m�8�x���|���w�5nk�jWX�V^@��%�w
�9�⽐캽����`���뻽B�����:�����pҾ\��6�\�W���e�ȿ# ���(�?�R�b��˂������R��:��0���ё���jc��?@��]�� �9ʿ�   �   a��E9M��D���ž��v�7�v���սaʽ,�ݽh��0#�.G� �m����� =��2\�������L�����R@������·���i�-fC�Gu��6��p׽{=Ľ��ϽNv��a4��/���þD���K�C������:�� �0�(wO�x~m����t���z��]4���N��6�l��*O��0�Z ��d��ܺ��   �   =.|��U7��F�Ͳ��w��;0���(W�������*� �9�Dh�8���,���pƾ�z޾���P���� �!���<�p�ܾ��þ0w��Qt��md�KM6����8���˺���u-�P't��0��c ��`6��9{�mۦ��տ:����ne8��4Q�Bf�t���x��ts��e�t2P���7���������տ�@���   �   %,Z�D���1�����a��*�����$��L�]����죾Ȯʾ�k�l���*��-�K�5���8�7<5��,�l���$�L��bȾ^��������H���!�����a�0�'��^��眾M%྿L���Y�v���3���Ԝ	����x�3�P-D�n�N�2zR��JN��C���2� ��n��}@�𝹿��   �   ��6��r��1��k,���[L���&�N��8.�2�U��r������#㾨�R�)��E��N^�K�q�h�}��̀���|�V=p���\���C��(�c��݄�J�%�����R�`�+����a%���J�ۚ��a;� h��7�~�s�����S¿��2��:��6�#�*,�N�.���+�V�"�������翾=��C���s��   �   ���<Gھ�瞾��k�	;��6(��41�� U��������ﾖj�R?��f�dȅ�]D��������ɲ�����=-��B!��N�����c��1=�*��~���j��Iz��=S�3�/��K'�2t:�A�k�����ھ���OF��h������j��L�ܿL�������D��U�����������ڿ=㼿4���{�}�SE��   �   ��G������J�x.���.��9K�����>���
��D��2I�ޒz������֮�YĿ!oԿ��޿]��x޿/6ӿ��¿EU���M��1mx�f�G��%�Ӌ��I��\��E�J��x.�2�.��7K�6����;���hB��/I���z�P���9Ԯ�Q Ŀ�kԿ�޿����޿�2ӿ�¿sR��mK��ix��G�T#��   �   �g���w��:S���/�9K'��t:�8�k������ھ��oRF�.l��Þ�%m��<�ܿ����x���F��W������������ڿ�弿����?�}��UE�܎�fJھ�鞾N�k�L
;��6(�d31��T�������y��g��?��f�ƅ��A�����|������󚪿N*�����ٕ��j�c�9.=�H�����   �   ~���8�R���+����a%���J�����DϾ��i��7�@�s�D����U¿��迸�����(�#�F,�x�.�Ԍ+�X�"���������$@��>��� s�\�6��t��3���-��l]L�G�&�~��>.��U�p��D��������)��E�,J^�t�q�Q�}�ʀ�o�|�q8p�6�\���C��(�y��5�ླ�   �   y�H���!����a�=�'��^�霾0'�,N���Y�����������	�*��H�3�d/D���N��|R�MN��C���2��������B�矹��򐿌.Z���	4ᾕ���ra��*��������$�&L�ʷ��W飾~�ʾ�f�Y��`'��,�K�5���8�285��,�����!����Ⱦơ������   �   �������"����v-�\(t��1���c ��a6��;{��ܦ���տ,��!��f8��6Q�^f�nt� �x��vs��e�d4P���7������_�տWB���0|�fW7� H��β�ww�Z<0����,U��T����'�.�9�>h����V����ƾ�u޾���j���� �4��/7�>�ܾ'�þ8s��q��d�,I6��   �   Bl׽o:Ľ��Ͻ�u��a4��/���þ��
�K��C������F�� �� �0�pxO��m����9u��|���5���O���l�,O��0�R!��f�+޺�[���:M��E��ž���*�7�{����ս�^ʽT�ݽ����#��G���m������9��cX�������H���	��v<������wˇ�c�i��aC��q��3��   �   4����^���껽������:�戌��Ҿѝ��\�ѳ��	�ȿ|# �x��ަ?�F�b�ŝ������S��!���0���ґ��Â��c��@@�v^��� �:ʿ�阿��^��3�,վ�����>����>½����䨽�]����r����(��GC���Z��:m�G�x��||���w�uik�	SX�iZ@�z�%�6t
�����躽�   �   �#��v݋�jݰ�R���r?�_��� ܾx"��Fg�L���:ҿ�7&�B�I�ҥo�~��� ���������	��a���0��Fup��J��X'�**��Կar��0�i���#���޾�W���[C�g%�8b���0��Pj�����g���ڽ����1��M(��u6�V?��B��{>���4�d&�ʎ�������ӽ�>��ő��   �   N�T�:i�3��d�὎P-����xɾ��H}S�ߚ��m���Z;��VB���7�jX���x�铊�NH��G����M������f{y��dY�X�8����ת����¿�Z��vQV��a�l�̾HL���3�p�콵���F�}�I�i��|�5�������սb����
�P��Ѹ����[���]�������rN̽,������Q�g��   �   �2g��Nu�t��c!�Y�+�p`���ƾ;��f+P�Y������������4���T�)t��Ç�3%��x��k���·�d�t�nU���5�>������꿿f���}�R�����ɾR��C�1���콈Ц�J����{��R���C���pƽ�콑�������%��x-�G�/�=B,�I#�H������&�=ʼ�n7��d���   �   �v���z��񩦽	����'���|�s����p�F�uň��i��_�翐>�\+,���I���f���aO��F���.��8a���f�L7J���,����t鿽����!��V�H��������U��J-�t��N���x�������������ԽX� ��v�Uc1���F��W�Zma���d�6`�֚T�kC�+,-��������Jʽ�����   �   �ȿ��[���
����F"��n�}1��y� ��j7�@�|�H�����ֿ����/��9���R� Ph�d�v��{�"4v�d�g�4aR��x9�^<���)�׿�����~� )9�6C�-첾s���&�u���s½���J�ɽ�F�D��4�)�W�bzy�ο�����9ޞ�v#������
��V���^�t��~R�;�/�������   �   ���P߽\lսt,�j��c�[�$���F�2<$�^lb�3���S��K��F��T&�hO;�f�L�0wX��R\���W�T�K�&O:��?%��}�[�N����� �c��]%��w龌ơ�{`�n���b��m	޽}�����(�5�R�0]��*����G��0-ɾ�Zھ,+�;��k5�E�ؾ�ƾ�}��������|�bM���#��   �   Y�4��p���������(�I�ފ��]ʾ���Y]D��Ђ�����;п[,��6P�b"��60�_9��T<���8��&/�~� ��K������aϿ���UȂ� �D��,��`˾�����L�Z��_�^������X9�Bik�M���y���ܾ~���l��h!���#��l&�:T#�����0��R����ؾ�!��\�����e��   �   8�t��=�:�������@7���v��5��1��x%���[�ˍ���ȯ���ҿ���N��V
��L���������j����(�пU���Ԍ��"[���$����Z���Ax�x+9��g�,6����D�A��3y��>���o;�����]��s2���H��Z�.�d��_h�.d��X�@�F�vK0�l?���7ʾ�q���   �   ���.(v���>�Q������(��U��Ï��ž���^�2�r�f�9u���F����ǿ�߿kP�����8� �5���W�𿆲ݿf�ſ񗪿W+��V�d��1������ľ挏��QU�$W)��d�˝ ��A��sy������ؾa�
��{,�.�O��q�%ć�}a��󥚿�𜿌���^�� |��8�n�~'M��C*�t��C:վ�   �   BXӾy:����j�<7�0������7�zl��x��6վ.��5��8b����1��"]���G��C�ɿl�̿��ȿW���칯�gn��k����_��3����UӾ=8����j��7��������7�c}l�{���9վ����5��<b�������`���J��x�ɿ��̿��ȿY��������p��������_��3�ұ��   �   ���s�ľ�����SU��W)�Xd�I� �@A��oy�ྤ��ؾ��
�rx,�B�O�g�q������^��"�������[���y����n��#M��@*����6վV���j$v�/�>�$�����(� U�tŏ���ž����2�ߋf�Sw��I��]�ǿ'�߿�S�W����� ������𿇵ݿ�ſB���J-��z�d�R�1��   �   s�$�M�����Cx�^,9�xg�5�s����A��.y��;���k;����rZ��o2��H�R Z�}�d�([h��d�!{X�:�F��G0�d<���=ʾ�n��ǉt�
�=�]��J���1B7��v� 8��B��%�z�[������ʯ�2�ҿ������"��N����`�����k�\���пY����Ռ��%[��   �   �D�S.�[b˾����L�2Z��^������)U9�(dk������t���ܾ����.������#�i&��P#�X���-�hM��>�ؾ���F�����e��4��n�0������R)�yI�6���~ʾ���_D��т�E��>п�.���Q�"�t80��`9��V<�v�8��(/�� �0M�����cϿ�����ɂ��   �   Ԅc��^%�zy龌ǡ�|`�����a���޽ y�0����(�H�R�#Z�������C��k(ɾ�Uھ�%徿��0�6�ؾb�ƾ�y��C�����|��M��#�����L߽pjս,������[�u���H羭=$�dnb��������F��t���&�Q;�B�L�4yX�
U\���W��K��P:�DA%��~�$��P������   �   g�~��)9��C��첾�s���&����&r½���5�ɽA�A���4��W��ty�����=|���ڞ����,��(��'�����t�zR�8�/��������Ŀ�BY��p	�����"�5n��2��`� �5l7���|�e�����ֿ����0�J�9��R��Qh�B�v��{��5v��g��bR��y9�H=�|�U�׿y����   �   "����H�	�'���V��k-����$����������	����Խ�� �Ws��_1���F�.W��ha��d��`���T�uC��(-��������zFʽ����mt��ry��@���3�㽌�'���|�t��c�m�F�ƈ��j��i��2?�$,,���I���f�`��P���F���/��zb���f�"8J���,�H��u�\����   �   ������R�4��)�ɾc��7�1�z���Ϧ�8�{�Q��MA��nƽ�콾�����y�%�[v-��/�@,��F#�b��0��$��Ǽ��5������0g�ZMu�Rt���!���+��`���ƾ���,P�sY������\�����t�4���T��)t�ć��%��zx������·��t��nU�ث5�z������꿿�   �   �Z��FQV�ta�5�̾L���3���g�����}�Ři�|�����j��Sս$����
�8��������P���]�������qN̽,���$���}�g���T��i�K3������P-�����ɾ��}}S����������;��lB���7� jX��x���UH��G���M������R{y�~dY�D�8����������¿�   �   ������R����R�ɾ�~��~1����6Ϧ����{��P��0A��nƽ�콺�����x�%�\v-��/�@,��F#�d��/��$㽹Ǽ�p5�����T0g��Lu��s��� ��+�H`���ƾ��,+P��X����m��`����4���T��(t�WÇ��$���w����0·���t��mU��5�������0꿿�   �   � ��T�H�������U��-�%��񧰽ȇ��z�������ЄԽ�� �Fs��_1�~�F�-W��ha��d��`���T�xC��(-��������VFʽP����s���x��.������7�'���|�xr��>�΃F�ň�]i�����>��*,���I���f�Ъ��N��WE��0.���_�d�f�P6J��,���s������   �   B�~��'9�AB��겾�r��&�F��~p½���t�ɽ�@��@���4���W�wty�����=|���ڞ����.��*��*�����t�zR�/�/����V��`Ŀ�NX��������"�_n��0��˸ ��i7���|�i�o�ֿ���.���9�F�R�hNh���v� �{�D2v���g��_R�nw9�T;�����׿l��   �   �c�,\%��u��ġ�`�U���^���޽�w����(��R�Z��t����C��h(ɾ�Uھ�%�ĉ�0�>�ؾg�ƾ�y��C�����|��M�Ӫ#����pK߽�hս2)�����[�歟�ND��:$��jb����������:��&��M;���L�>uX��P\���W�z�K��M:��>%��|�Z���L��{���   �   аD�^+�8^˾2�<�K��W�P]����6���T9��ck�䍔��t���ܾ����,������#�i&��P#�[���-�jM��<�ؾ���8�����e���4�n�.�������&���H�t���nʾ3��[D�Qς����:п*���N��"��40�]9��R<���8�%/��� �XJ�����_ϿR����Ƃ��   �   ^�$�c������u=x��(9��d�^3�Y��$�A�@.y�};��yk;v���jZ��o2�~�H�R Z�~�d�*[h��d�&{X�>�F��G0�d<� ��4ʾhn��o�t�m�=�`���}�T�x>7���v��3��j��%��[�-����Ư�=�ҿ�󿾍����J�̖����*�lh�����п(���;Ҍ� [��   �   �����ľ����pNU�0T)��a��� �3A�oy�����nؾ��
�gx,�9�O�a�q������^��#�������[���y����n��#M��@*����u6վ-����#v�<�>����K�x�(��U�����6�ž�����2�L�f�Gs��RD��ڳǿ�߿'M�`���v� �������p�ݿ��ſ���B)���d�2�1��   �   dQӾ5����j�^7������2�7�$yl�7x���5վ�ܐ5��8b����.��!]���G��D�ɿn�̿��ȿ\���﹯�in��m����_�
�3�����TӾ�7����j�T7����w���7�cvl�v���2վ��
�5�.5b�������\Z���D���ɿ8̿��ȿO�����k��0���.�_���3�:���   �   7����v�|�>������(��U�'Ï���žy��N�2�g�f�4u���F����ǿ�߿jP�����8� �8���Z�𿈲ݿh�ſ򗪿W+��S�d�޹1������ľ�����PU�HU)��a��� ��A�Yky������ؾH�
�Zu,���O��q�4���&\��^���D뜿���8Y��w��z�n��M�e=*�g��u2վ�   �   ��t��=�1���|�(�J?7���v��5�����g%���[�ȍ���ȯ���ҿ���N��V
��L���������j����)�пW���Ԍ��"[���$�z�����@x��)9�5e��2����0�A��)y��8���g;}���cW�Dl2�|�H���Y���d�zVh��d��vX�'�F�BD0�>9����ʾ.k���   �   Ӏ4�jk���� ����&�� I�v���ʾ{��N]D��Ђ�{���;пW,��4P�`"��60�_9��T<���8��&/��� ��K������aϿ���UȂ���D��,�^`˾����� L�/X��\�M����SQ9�4_k�֊��
q���ܾ'�����y�\�#�je&��L#�����*��G��`�ؾ����|����e��   �   ד��G߽4fս(����l�[�֮���E�%<$�Vlb�0���Q��I��D��T&�fO;�f�L�2wX��R\���W�V�K�&O:��?%��}�]�N������c��]%��w�Gơ��`�����^��-޽�t�@��=�(���R�8W�� ����?���#ɾ�Pھx �]���*�*�ؾ��ƾiu��������|��M��#��   �   a����U��3����;"�&n�E1��j� ��j7�:�|�G�����ֿ����/��9���R� Ph�d�v��{�"4v�f�g�6aR��x9�`<���,�׿�����~��(9�+C��벾l s���&�J��co½�����ɽ�;��=���4�9�W��ny�]����x���֞��������������t�uR��/�l�����   �   nq���v�������O�'�4�|��r����k�F�sň��i��_�翐>�\+,���I���f���aO��F���.��:a���f�N7J���,����t鿾����!��U�H��������U���-�d��d���p���Y������Խ� �Up�+\1���F��W�Hda�x{d�.`�A�T��C�%-�������Bʽ�����   �   �-g��Ju�s��e ��+�U`���ƾ7��d+P�Y���������� �4���T�)t��Ç�3%��x��k���·�d�t�nU���5�>������꿿g���}�R����ɾ8���1����Ϧ�P��{�}O��d?���kƽ��$�������%�Kt-��/��=,��D#�������!�>ż�W3��"���   �   j�.�u�@�t����J�����Tg��߮�� �[8���}�����b�׿�M�J����:�^_T��@j��+y�z~�3y��oj�b�T�Ά;�r� ��p��ٿ_���$����;�B\�ri���o�� ��ѽ�����eb���P���`�;��J���I���/�ٽ�t󽎠�@�	�t����nm �_K�;νF'�������Kh��?��   �   �?�1�K��䃽�����Mad��M�����*)5���y����ڃԿPO��j�D�7��P�Z�e��Zt��uy��Pt�l�e��Q�nX8�\O�$S���ֿ=���B}���7�zD� ���.�l�Y��R�ѽ2J��q�l���`��v������A�н��v��Ĩ�&R��
�����j�h��m��Wý� ��>��kU��   �   Z�p��cm��"���4ý
D���[��㤾���,��un�����M˿���R�v/�*6F�p�Y�`�f��Uk�:�f�roY�t&F�&D/���7e��*�̿����/q�>4/�~k��ۨ�Bzc�K���rҽ�Ϝ��Ɔ�d���Tp�������Y����'f�O�.��
=���E��7H��
D�.�9�L�)��n��� ��Fս�����$���   �   i�����ɳ���ǽ>b�[O�6t��)#�6��4b\�����)��g�迲H�ؼ!��d6�iG�$�R���V��LR�*�F�$�5��{!�FS�tR���᭓�FU^�͆!����V̜��U�Z���Խ ;���8������ս.�H��e	>��o[��ru�xۄ�B&��w���c/������Jp��"U�U�6���j���7�Ž�   �   	�⽐����.���ϽTE�0�?�|3��H�ɾ@��JE�~������Nѿ_{����R#�$s1���:���=�HN:���0�."��v�s���_ѿ�#��D샿fhF�2@�#̾�ˍ���D�r���3۽�4Ľ�ͽ�q�C���9�>�c�hڇ��6���)������!AȾ�˾E$Ǿi༾�C��H�������[�?�1�&���   �   3��}���ߓ۽�`ݽ�M�'2/��w�TC�������+� 6d�咿WX��pڿ����̹�����l!�<�#�R� ���ȴ����	ٿ����O����%d��t+�M����̱��z��:3����z罌����f#�BO�֐��� ����߾���EH�x����Y���۩��̭۾����Ŝ�G.}�9�G��   �   &�T��)%�j�0��������ܝW��o����Ѿ���T�?��%w�븙��|��`�տ�pￒ�����2�	��v��� �b��ӿ�㶿�����u�$�>�����
ҾU��M�Y�&�"�J�����l ���*�A[�3���������޾������/��4>�`�G�̣J��F���<��-�Cp����^�ھ�课���   �   ش��m�V��)&�h
�����K��t:�ԙ{�����|��� I���z�𧖿�ޮ�8
ĿanԿ>�޿��$�ݿ�ҿ-¿� ������w��CG�}���K�0۫�|{�t�:��f�_����T�)�p�Z��n������"�}��&H5���R�Ym�y������%��挆��t��j��"P�y�2�'�v����   �   �:���:���:M�� ���	��a
��D!�cQO�I̊��s���V��vp��iE���m�D/���%��RL�������Xͯ�b
��a���	����j���B�i��G�8���8��18M�a ���	�-b
��F!�FTO�vΊ��v���Z��&s�&mE���m��1��U(��O���������%Я�	��ғ��7���ʫj���B�k��K��   �   �N�aݫ�Z{��:�4g���I��)���Z�Bl����򾤑��D5���R��m����~�����s���"p��~j�%P�<�2�W$�6 �T���v����V��'&��f
�����L��v:�!�{�u������e	�"I�R�z�!���ᮿ�ĿYqԿU�޿<��/�ݿ��ҿ�/¿�� ��x��FG�����   �   6��Ҿ���!�Y��"�1������
��*�[�Y��K�Z�޾L�����B/��0>�D�G���J��F�'�<�,-�*m�Y��}ھJ対2F�T�+'%�ph�����������W�mq����Ѿ���ͼ?�)w�ٺ���~����տ�s� ��$����	��x�&� ��d��ӿ�嶿����̷u�a�>��   �   7v+�����<α�Ǡz��;3�����x罜���
�Cc#��=O�����>렾з���߾"��6E�F�x�~V���f�����۾���������(}��G�(��R���k�۽�_ݽ�M�f3/�w�+E��3����+��8d��撿;Z��Grڿ���<��L���n!���#��� ����$��A"��ٿa��������'d��   �   �iF�AA��̾�̍���D�����2۽�2Ľ��ͽ�l�"@�h�9��c�8ׇ�3���%��4���j<Ⱦ�˾�Ǿܼ�{?�����������[�6�1�
��t��w���	-��?Ͻ�E�z�?��4���ɾ���LE�-�������Oѿl}��!��#��t1�,�:�j�=��O:��0�j/"��w�T����ѿ0%��D탿�   �   |V^���!����͜�ƫU����Խu9��v6����I�ս+�����>��j[�8mu�]؄�#��/���.,��� ���Dp�U��6��������Ž�e����������ǽ�b��O�9u���$�T���c\�{����*����迒I��!��e6�tjG���R� �V�`NR�t�F�D�5��|!�T��S��������   �   V0q��4/�Cl���ۨ��zc�g��4rҽ�Μ�ņ����4m�������T�&���b���.��=�{�E��3H��D�d�9���)��k�߮ �QBս����!��A�p�am�2"���4ý�D���[�c䤾����,�wn�����9˿5���S�>	/�7F�z�Y���f��Vk�R�f�lpY�J'F��D/����f��ߖ̿7���   �   fB}��7��D�)���P�l�T����ѽ�I����l�(�`���v�������i�н�
񽯳�ݦ�+P���ˢ��h����j�AUý�������`hU�?��K��䃽$���O���ad�TN��֡���)5���y����e�Կ�O�@k���7�z�P���e�f[t�"vy�xQt���e�0Q��X8��O�XS�ڋֿy����   �   
����;�#\�Ei����o�� ���ѽ����deb�J�P�_�`��:����������ٽ�t�x��(�	�b����bm �RK�;νF'�������Kh�-�?���.�Ʀ@�����&K��Q��Ug��߮�'� ��8�0�}�������׿�M�^��ƹ:�r_T��@j��+y�z~� 3y��oj�T�T���;�`� ��p��ٿA����   �   YA}�@�7�D�n���S�l���� �ѽ�H����l���`�D�v�|�����V�н�
񽨳�ܦ�*P���̢� i����j�=Uý����o��$hU��?�e�K�6䃽Y������ad��M��ˠ���(5�~�y�U����Կ"O��j���7���P���e�0Zt��ty�>Pt���e�:Q��W8��N��R���ֿ���   �   V.q�]3/�4j��3ڨ��xc�)���pҽ�͜�UĆ�z����l��s����T����b���.��=�z�E��3H��D�e�9���)��k�ܮ �<Bս謬��!��~�p��_m�8!��m3ýVC�)�[�㤾���,�,un�z����˿J��rR��/�^5F�~�Y�N�f�|Tk��f�bnY��%F�XC/�^��d��;�̿����   �   �S^���!���!˜�1�U�����Խ�7��j5��F ����ս�*�d���>��j[�,mu�Z؄�#��/���.,��� ���Dp�U��6������}�ŽPe�����H����ǽ a�O�[s���!�^��
a\������(��/���G��!�pc6��gG���R��V��KR���F���5��z!�bR��P�� ��ଓ��   �   �fF��>�4	̾=ʍ���D����"0۽�0ĽY�ͽ�k��?�1�9���c�&ׇ�3���%��0���j<Ⱦ�˾�Ǿܼ�|?�����������[��1�ܔ�Ծ�p���e+���Ͻ�C��?�a2��Ɓɾ1�zIE�}��P󨿙Lѿ�y����#��q1���:�&�=��L:�"�0��,"�fu�]����ѿu"��냿�   �   �r+�w����ʱ�ћz�H83�}���u网��
��b#�G=O�Ս��$렾������߾��5E�E�y��V���i�����۾���������(}���G�ѕ�3�����۽]ݽ�K�(0/�:
w��A��$��� +��3d��㒿�V��nڿ/���t��<��Tk!���#��� ����\��N���ٿ��������#d��   �   ����Ҿ?��"�Y���"�������{�
��~*��[�.��+�@�޾B�����>/��0>�E�G���J��F�(�<�0-�+m�X���|ھ@対��T��&%��g�������Y��0�W��m����Ѿ?���?�#w�)����z����տn��������	�Tu�� �=_��ӿWᶿ���±u���>��   �   H龆ث�~{�W�:��c�է����)��Z�l������򾗑��D5���R��m����~�����u���&p��~j�'P�<�2�T$�, �@���Q�����V��&&��e
�����I�r:�X�{�����G����^I�5�z�㥖�#ܮ��Ŀ�kԿ9�޿	���ݿ�ҿ_*¿C�������w��@G�#���   �   �4��[6���4M�m ���	��_
��C!��PO��ˊ�hs���V��jp��iE���m�A/���%��QL�������[ͯ�e
��c������
�j���B��h��G��7���8��m7M�% ���	�F_
�UB!�NO�ʊ��p���R���m��fE���m�-��Y#���I��}��9���ʯ����㎙�ʆ���j���B�Uf��C��   �   �����V�c$&�?d
�J��,J��s:��{�����Q���I���z�맖�}ޮ�7
Ŀ`nԿ?�޿ ��%�ݿ�ҿ-¿� ������w��CG�w���K�۫��{�f�:��d�ԧ�� ���)���Z��i���������wA5��R��m�Ƶ����*�����uk�jzj�DP���2��!����ì���   �   ��T��#%��e����~�����W�Po����Ѿ���G�?��%w�渙��|��\�տ�pￒ�����4�	��v��� �b��ӿ�㶿�����u�!�>�����
Ҿ��l�Y���"�$�������
�_|*��[��|�����޾�������/�	->�>�G���J��F�J�<���,��i����txھ�᯾J쉾�   �   ���������۽�[ݽ�K��0/��w�C��X����+�6d�咿RX��pڿ����̹�����l!�>�#�P� ���ȴ����	ٿ����O����%d��t+�4���|̱�5�z��93�����t�I����_#�<9O�.����砾����0�߾���<B�" �F�ZS��������۾Z���*���"#}���G��   �   ������8)���Ͻ�C�I�?�03���ɾ1��JE�~������Nѿ\{����R#�$s1���:���=�HN:���0� ."��v�s���_ѿ�#��E샿ehF�)@� ̾hˍ��D����/۽$/Ľr�ͽwg��<�>�9�ǭc�&ԇ��/���!�����7Ⱦ˾Ǿ�׼�o;����������[���1�����   �   �a��-��¯��ǽDa��O�t��
#�+��-b\�}����)��e�迲H�ؼ!��d6�iG�$�R���V��LR�,�F�&�5��{!�HS�vR���⭓�DU^�Ȇ!�}��*̜�n�U�f���Խ�6��p3��=�����ս(���� >��e[��gu�^Մ��������)������b?p�U���6�k�������Ž�   �   ��p��\m�7 ���2ýjC���[�v㤾��	�,��un�����M˿���R�v/�(6F�n�Y�`�f��Uk�<�f�roY�t&F�&D/���7e��+�̿����/q�<4/�pk��ۨ��yc�����pҽ͜�'Æ�����9j�����<P佂���_�L�.�>=���E��/H�D���9�\�)��h�&� ��=ս&�������   �   T?���K��ヽ������ad��M�����')5���y����كԿPO��j�D�7��P�\�e��Zt��uy��Pt�n�e��Q�nX8�\O�$S���ֿ=���B}���7�vD�������l���h�ѽ�H����l�
�`���v���������н����&��]N�����<g���g彥RýO������3eU��   �   ]Q�%���vL�؝��a���B�=��ϰؾ����V�9���G����q����^��u1�.B�~%M��Q��)M��/B���1����$Q��?俽Ӹ�[���JY���bi޾����O�M����|����i���L��0=���J� l��@��ä�\���s�ѽ�jὌ�꽞/콾����׽��ý佪��H��
�g��6�K��   �   C��N��G�Q�6D��7^���?��~`վ�o��R�Bb���3���߿�}���J�.���>�t�I��[M���I��>��.��k�,���]嵿q���U��Q���ھ#f��k�J����g���������T�V�J��>]��Ɓ��������1zн��mL��n��"�������ｺ�ٽ �������`���I�N��
&��   �   ��=�)#;��7b��۟����{�8�"Ŋ���˾�i���H�p������'տY#������q&���5�2r?���B�^L?��V5�pe&���E���gDֿb`���H��v�K����<�оD�����B�t�����Lu��y�o��s�j����ѥ�-ǽ������j��Vx!��m(�D*��&�S����������ս|���E���`��   �   �R��Y�n����8������$�-�}A��sμ�Sp���9�Y�w��Q���ſ}�쿴
	�|���_'��%0��3�n�/�"�&��}�d��k�쿷ƿ�
��2yy�[�;��`����C{���7�8����5��<���t���zl���"��VC�Z0
�ن#��<���Q��>b��nl�[o���i��n]���J��83�8��z����˽r���   �   h ��K@���8�����9�ὸ!�6�j���|
�}:&��]��Ꮏ�r���Կ�Z��
�j���i�b���	��D��q	��Q��7Կ�D���
��l�^��R'���㬾�fq�X�(������������\��C�ѽJ�5E ��C��Sh�����ɺ������$���Pī�LI���w���#��D����^�[o8���7X��   �   &��=@ѽ�����:�۽���u�P������Ѿ6;��n@�Q x��X��C���ֿ���h�z����
��^�H����DGտf)��I���Z~w��]@�����
Ӿx���h@U�&���UZǽ*Hǽ��w��22���_��C��zޣ�������Ծ�h�]��h���!𾕤��о�������������T��~'��   �   ��2���
����DK̽�ٽZ���i6�`�~�jn��l��U�!�P�}恿s/���D���9˿�Bܿ���]K�V�1�ڿ�ɿo���=Κ��߀�&-O��� �V,򾂅��d����8��
��c���׽x��gF�(�;��q��!��%2�����������Q� �6o(���*��'�������c'�%�ݾ�㷾����!h��   �   ��n�k�4�����齗?޽�����EnU��M����ƾ�����)�<|S���~�j���5��� ���弿���/���ٲ�S~��,U���{��Q�m�'��f���ľ�F��g�T�	x�1��ɖ㽟�����;�:��v�����;������2�@H�*TY�Vd�Uwg�"c��uW�f�E�"E/��I�9X��GaȾ�r���   �   �n����g�:�-��a�֝�����	��c0���k��#��tsо6���&�K�H� ii��"���Z��0]������l��?��j���P\f�6�E�s	$�`����̾`l��^�g��-��`�&�����>	�f0�>�k�C&���vоx����&���H��li��$���\���_������Ĕ��A�����`f�e�E�$�x��6�̾�   �   ��ľeH��ݦT�yy�#2��B��r�����'�:�^�u�"����;W�����\2��H� PY�d�sg��c��qW�ʟE��A/�G��S���]Ⱦ:p����n���4������a?޽i!��~�qU��O����ƾ���)�)�]S�;�~��������t#��輿+����1��ܲ�����4W��d�{��Q���'�|h��   �   $/�|������g�8�
��c�c�׽H���C���;�R�q����F.����=�����~ ��k(��*���'�N��Į��$��{ݾ෾�
��h�;�2���
�����I̽H�ٽF���k6�a�~��p�����j�!�o�P�"聿e1��G��<˿gEܿj��#N�"���ڿ=�ɿ����К�ဿ�/O�g� ��   �   !���Ӿɳ��BU�����>Yǽ�Eǽ�佫��n2�Ă_��@���ڣ�����ɃԾ�c���������𾎟㾆�о����"����݃�i�T�-{'�����<ѽg��2����۽ă�g�P�#┾(�Ѿ�<��p@��"x�eZ��E��=�ֿ���i���� �
�`������QIտ++��ƪ����w��_@��   �   �S'�����䬾hq�$�(���J���ȣ��l���ѽ3G��A �z{C�[Nh�����K�������.���M���aE���s��C ��C���u^�k8�����R�u���=��#7����� ���	!��j�-󩾣��;&���]��⎿t��ܬԿ�\��6
�����j����@��E��r	�wS���Կ�E���� �^��   �   b�;��a�����{��|7������5������W���si�����)>�,-
��#�I <���Q��9b�il��o�N�i��i]��J��43�g4��t����˽� ��*P����n���������� �-�TB���ϼ�Bq� �9��w��R��_�ſ��쿎	�r���`'��&0��3���/�&�&��~�,������ƿ����zy��   �   (�K�H���о����^�B���4���qt����o��s������Υ��(ǽ ��8��X��u!�Hj(�� *��&����������X�ս�����A��`�V�=�� ;��6b�ܟ����N�8��Ŋ���˾;j���H��������(տs$��j���r&�p�5�s?�^�B�4M?��W5�f&�D�3���*Eֿ�`��]I���   �   f�U��Q�9�ھGf����J����$���;��� �T�5�J��;]��ā�弚�����hwн��(I�����l�����������ٽ����I���}���=�N�Z&����?���Q�eD���^����?��$aվ&p���R��b��4��߿0~�z����.�0�>��I�Z\M�*�I���>�X�.��k�F,�=�࿢嵿����   �   `JY����/i޾�����M����7����i��lL��0=���J���k��@���¤� ���9�ѽ�j�^��x/콝����׽�ýܽ���H����g���6�i��Q�j��RwL�\؝�Sb��	B�i��
�ؾ����V�T���f����q����^�v1�:B��%M��Q��)M��/B���1����Q��?信Ӹ��Z���   �   ��U�XQ�N�ھ�e����J�e��V�������L�T���J�^;]��ā�����v���Pwн��I�����j�����������ٽ����A���n����N�&�@����	�Q��C���]��ٓ?�\C`վ�o���R�b��O3��6߿�}������.�`�>��I�l[M�B�I���>���.�Tk��+�W���䵿���   �   v�K���&�о|�����B�w�����`s���o��s�R���JΥ��(ǽ���"��F���t!�@j(�� *��&����������N�ս�����A���`���=��;��4b��ڟ����ǌ8��Ċ��˾
i�W�H����y��H'տ{"��B��:q&��5�fq?���B��K?�V5��d&��&���rCֿ�_��?H���   �   
�;��_�����;z��=7�����q3��~���G����h��1���=��,
��#�* <���Q�{9b�il��o�I�i��i]���J��43�^4��t����˽V ���O���n�;��B��������-��@��oͼ��o���9��w�Q���ſ:���		�����^'��$0��3�P�/��&��|������m ƿ�	��ywy��   �   Q'�����ᬾ)dq�p(�2�򽺽�����&���ѽ�F�IA �@{C�/Nh�����?�������)���L���`E���s��A ��B���o^� k8�v���R�����<���5��M�����8!�Q�j�j𩾲�B9&�c�]�����7q����Կ�X��
�B��ph�����NC�|p	��O��qԿC���	��m�^��   �    ��GӾ�����=U����rVǽ�Cǽ=�+��2�y�_�t@���ڣ�r�����Ծ�c���������𾏟㾆�о��������݃�P�T��z'�:���;ѽ����	���۽���H�P�#ߔ��Ѿ�9��l@��x�RW��\A���ֿ?��Tg�(��b�
�b]����+ �Eտ|'�������{w��[@��   �    )����:���8�ȃ
��_㽋�׽I��4C��;��q����$.�����4������} ��k(��*���'�P��Ʈ��$��{ݾ�߷��
���h���2��
�]��wG̽{�ٽl��Xg6�S�~�Xl�����t�!�V�P��䁿�-���B��77˿6@ܿ��濠H꿟濖�ڿt�ɿ<���O̚��݀�x*O�e� ��   �   ��ľED����T�Wu�e,��P�㽵����~�:���u������;9�����R2�~H�PY�d�sg��c��qW�̟E��A/�G��S���]Ⱦ&p��Z�n��4�%��齸;޽���|�BkU��K����ƾ��N�)�TyS��~�c������r��C㼿ݣ��q,��ײ��{��S��3�{��Q���'��d��   �   �i��A�g��}-��]�����꽛	��b0��k�z#��Msо'��ޞ&�@�H��hi��"���Z��0]������m��?��k���R\f�8�E�r	$�\����̾Bl����g�^�-�j_�̙齺�꽐	��`0���k�4!��.pо��F�&��H�Kei�� ��TX���Z��,������6=��H���}Xf��E��$���u�̾�   �   ��n���4��� ��:޽������mU�JM����ƾ�����)�0|S�v�~�e���2��� ���弿����/���ٲ�T~��-U���{��Q�j�'��f���ľ\F��ϣT�w�.��[��*��c����:��u�L���!;ʒ����&2��H�1LY��d��ng��c�nW��E��>/�AD��N���YȾ7m���   �   \�2��
�	�ཪE̽#�ٽ����h6�~�5n��F��F�!���P�x恿o/���D���9˿�Bܿ���_K�Y�3�ڿ�ɿq���>Κ��߀�$-O�}� �D,�a���(���8�Є
�%`㽇�׽���A���;���q�����*����⾜������z �Zh(���*�>�'���ǫ�"�wݾ-ܷ����h��   �   l���7ѽ=��|��
�۽�����P�Z�����Ѿ);��n@�G x��X��C���ֿ���h�|����
��^�J����DGտf)��I���Z~w��]@�����
ӾI����?U�)����Uǽ�Aǽ�	佴���2�~_��=��Zף�p���0Ծ�^澵�����r𾇚��о���������ڃ���T�Cw'��   �   ����9���3��n
������!���j���]
�r:&���]��Ꮏ�r���Կ�Z��
�j���i�d���	��D��q	��Q��7Կ�D���
��l�^��R'���r㬾!fq���(�.�򽌽���������g�ѽRD��= �wC�%Ih���賕�6���O���]���A��,p�����9���.^��f8����L��   �   �L����n���������齋�-�JA��Sμ�Hp���9�R�w��Q���ſ{�쿴
	�|���_'��%0��3�n�/�"�&��}�d��k�쿷ƿ�
��0yy�Y�;��`�����{��L7������3����������f�����9�*
�m#��;���Q�x4b��cl�co���i�vd]�K�J�Y03��0��n����˽T����   �   ��=��;�$3b�Pڟ�����8�Ŋ���˾zi���H�o������'տX#������q&���5�4r?���B�`L?��V5�ne&���F���gDֿa`���H��v�K����-�о,�����B���踷��r��*�o�Ĥs����g˥�%ǽr�꽜��p���q!��f(�m�)�F�%������I�����ս�|���>���`��   �   G��<~��Q�hC���]���?�vt`վ�o��R�Bb���3���߿�}���H�.���>�t�I��[M���I� �>��.��k�,���]嵿r���U��Q���ھf��@�J��������������T�V�J�w9]�XÁ� ���{����tн@��<F��2�����v�������ٽ���
���������N��&��   �   �İ��,˼����s�psƽ���Io�.W������U.���h���s(��X߿HS��;�& �nU&��;)��W&���&u����:࿴���@l����k��q1�p@�P@���H~�*�-�Sr�4���0�o��D�PD8��C���\�b�J��xݣ�P�����©ý�ý�&��\���᜽�Ԇ�У]��	.����ʼ�   �   ^ɼJ�ۼT�yt�q�Ľ}��H�k�_���F%����+��?e�/���T��O�ۿ����$�\��J�#��}&���#�n���'��b���ܿj�������0h�~�.�HU��E\���pz��i+��&K��w�r���J���B���Q�#�o��[��+������9Ž��ѽ�Nؽ�ؽ��нf�½ J���k����z�H�F�65�`��   �   �	��u��(���w������9���a��������L�#�}�Z��猿�����ѿ�\�r��\�������:���=�@��C���ҿ=믿W���Z�\��.&�H>����eWo���$��k�]���8�|��_�Wc���~�X1������c˽�潛�������:^��M����+��mCʽ�ɩ�����JV��_&��   �   �I���3��}B�F�J������>�R������ ۾}H��J��N������}¿��Z���B	��,�T~����`��I`��77�و¿)k��r炿��K�#�8n߾����3^��T���ٽv���V[���#��荽d����ǽ�RE�Ċ�\S/��<�(�C�&�D��@��,5�7 %�qN�����	8ʽꊠ���z��   �   �撽�tt��i�԰��״����7�?��Ҋ�ٵľ����4��si�,W��򝮿��ʿ,�Sj���N��O���l����?⿘�ɿM&���1��^�i�1�5�
���Ǿw���j�H�����&Ͻ����� ��(ɝ�������߽R.	�o�%��C�;x_��Zx��ą�m���6���䉾'n��*�n���R�rD4����ެ������   �   �wѽj��O��9����ڰ����*�i�s�W���t|����`�J��g|��З��M���ſ�ֿd�5u�w��տa�Ŀ�1���𖿰@{�&�I�����1����P�x�e!1��_ ��Ž�몽૽XpĽ��)��5<��oe���������,%��\�ž\Ⱦ�9ľrڹ�$9���Ɩ�F0���IV��O,����   �   �����߽]��?z������4ܽL��;"Q�|���ϭƾ��W0*��'T��s��}�������紿0̽�����2���س��m���-��6#}�\SR�p�(�J9�%�ž����r�R��6���=5��Ժ���sʽ`���:���?J��~�����sѺ��&ؾ %��9�x�	�[s�������j�aҾ�X��-�����p���<��   �   �B�$X�1��/���QX���c̽jB��0��q����_�׾b�
��,���O���q��釿֎���ښ�)��FJ��c��������o��FM��X*�?����Ծ�㠾�1n�?�.����ѽk����cɽ����L��L����K/��v*Ѿ����^��r#��k1��,:��<�D?9���/�!�~�������˾�;�����   �   ��}�\�=��:޽0(��s����n�Xw�!�C�ޤ������d~۾L���#���>�D:V���h�N3t���w�*-s�оf���S�"�;�r!����־I5����}���=�J�޽�'��,���q�Fy��C�񦂾�����۾KN���#�Ӡ>��=V�Ԫh�P7t���w� 1s���f��S�.�;�
!���`�־�7���   �   栾
5n�P�.�D���ѽ���0bɽr��NJ���L�P��7,���&Ѿ�������o#��h1�{):���<��;9�F�/�!��������ʾ�8��\���B��U��㽌���X���d̽�C��0�q�����׾m�
�t�,���O�;�q��뇿󐓿ݚ�G+��qL��s�������o��IM� [*�(����Ծ�   �   p�žU�����R�W8��C5������pqʽ]���]��<J� �~������ͺ��"ؾ �7���	��p�������e��\Ҿ_U��,�����p�Е<�.����߽���y�������5ܽȢ��$Q�G���Q�ƾ���2*�v*T�w��������$괿yν�^����4���ڳ��o���/��;&}��UR�q�(��:��   �   �3쾛
����x��"1��` �5�Ž6몽ޫ�8mĽx�&��1<��je�0������H���!����ž�WȾ85ľ[ֹ�e5��NÖ�p-��8EV��K,��2sѽ�f��1M��s���۰���｣�*���s�,���뾊����J�Ej|�+җ��O���ſ=�ֿ��zw�Ey���տL�Ŀ_3���'C{�"�I�j���   �   ����Ǿx�����H�A��C'Ͻ;���P����Ɲ�������߽\+	�ǚ%��C�$s_�NUx�����3�������ቾk����n���R�/@4�����M���?㒽(pt�i�i�l����״�a����?��ӊ���ľ��P�4�vi�kX��h���[�ʿ�-�Rl���O� Q���W����A�(�ɿ�'��3��,�i���5��   �   �#�mo߾����	5^�3U��ٽ9���bZ���!���卽�`����ǽ�MB�4��^O/�:<���C���D�@�d(5�O%��J������2ʽˆ��7�z�I�d�3��{B��E�ﳺ������R����� "۾�I��J��O������~¿m�������B	��-�8�^��.���a���8��¿l��/肿�K��   �   $/&�?�7���Xo���$��k�3����|�ƕ_��Sc�g�~��.�����_˽潇������X[��J�����.���>ʽ�ũ�\���EV��[&��	��s��(���w�!���::���a���������#���Z�S茿�����ѿ�]����\�V �V�����>�Ɓ�,��łҿ�믿����!�\��   �   ��.��U��|\���pz�j+���J����r�Q�J��B�V�Q�F�o�*Z�� )�����X7Ž˸ѽ�Kؽؽ��н��½�G��Qi����z��F��2��[�bɼt�ۼ�S�myt���Ľ�����k�䯭� &��0�+��@e������T��־ۿ���v������#��}&��#����(�3c��y�ܿ���������h��   �   �q1�V@�*@���H~��-�r�������o��D��C8��C� �\�����>ݣ��������ý�ý�&��<���᜽�Ԇ���]��	.����ʼ�İ�-˼G���s��sƽ����o�_W��*��V.���h��󕿍(��s߿US��;�0 �rU&��;)��W&���u�ع�v:࿛���+l��r�k��   �    �.��T���[���oz�Xi+��?J����r�t�J�k�B���Q���o��Y���(��c��>7Ž��ѽ�Kؽؽ��н��½�G��Ni����z���F�n2��[��ɼ��ۼ�R�8xt��ĽG���k�-����$��|�+��?e������S����ۿ���� �����#�:}&�`�#���z'�,b����ܿ����B����h��   �   �-&�=�����Vo���$��i�ȕ��Ҕ|�-�_��Rc�P�~�$.��Y���R_˽��R������K[��J�����"���>ʽ�ũ�J��FEV�[&�m�	��r���(�z�w�l����8��a�h������­#�¬Z�3猿G��0�ѿ\����[���
������<����7���ҿp꯿�J�\��   �   �!��l߾����E2^�FS�X�ٽ<����X��� ���䍽�_���ǽ.M�jB���9O/�<���C���D�@�\(5�J%��J�p����2ʽ������z�5I��3��yB��B����������R�����l۾�G�~J�N������|¿�~�����PA	��+�v}��������^���5Ῑ�¿j���悿W�K��   �   ̠�@�Ǿ���b�H�����#Ͻֹ������{ŝ������߽�*	�u�%�@C��r_�$Ux�����)�������ቾk����n���R�$@4���ߦ������Ⓗ�nt��i������Դ�>����?��ъ�_�ľ��\�4�?ri�V������/�ʿM*�th���M��N���u���>���ɿ�$���0��N�i���5��   �   �.���f�x�+1��] ���Ž�誽.ܫ��kĽM�&�S1<�Mje�������2���� ����ž�WȾ35ľWֹ�a5��JÖ�j-��(EV��K,��
��rѽf���K��Z����װ���9�*���s�����3z�V��p�J�,e|�"ϗ�GL��-�ſ�ֿ7��r��t࿿�տb�Ŀ�/����={���I�%���   �   ��ž����|�R��4��罍1��𶶽uoʽ�������;J���~�X����ͺ�t"ؾ��7���	�p�������e��\ҾXU��#�����p���<����ʟ߽u���v��t����0ܽM���Q�Ɔ��|�ƾU
�Z.*�J%T��p�?|�������崿�ɽ�ʟ��L0��jֳ��k���+�� }��PR�<�(��7��   �   ]ᠾ6.n�`�.�����ѽ�����_ɽ���I���L���,��q&Ѿ�������
o#��h1�x):���<��;9�E�/�!��������ʾ�8��7�b�B�VU����}����T��:`̽_@��0�W	q���h�׾y�
���,���O�[�q��燿ʌ���ؚ��&��H��N���ј��Do��CM�V*�/����Ծ�   �   K�}�*�=����޽�#��%���zl�{v�}�C���������:~۾�K���#���>�=:V���h�M3t���w�,-s�Ծf���S�"�;�q!����־:5����}�4�=���?޽�$�������j��t���C�΢������z۾�I�9�#���>��6V�B�h�_/t���w�4)s��f��S���;��!����E�־f2���   �   ɳB��R�A��r���8T���`̽^A��0�)q����4�׾P�
�ڮ,���O���q��釿Ԏ���ښ�)��FJ��e������o��FM��X*�<����Ծ�㠾�1n���.�8��ѽ����p^ɽ��|G���L����7)���"Ѿf���	��l#�le1�&:� �<�r89��/� !�4�����,�ʾs5��j�~��   �   �����߽����`u������1ܽl���!Q�C�����ƾ��H0*��'T��s��}�������紿0̽�����2���س��m���-��6#}�YSR�l�(�E9��ž�����R�M6���	2��4���tmʽw���B��*8J��~�v����ɺ�Kؾ;�z4��	��m�X��T��a�kXҾ�Q��	�����p���<��   �   �mѽ�b���I��<����װ�	��`�*���s�+���S|����T�J��g|��З��M���ſ�ֿc�8u�w��տc�Ŀ�1���𖿰@{�$�I�����1������x�� 1��^ �R�Ž>誽�ګ�'iĽd	�d#��-<��ee�O��]����������žTSȾ�0ľDҹ��1��𿖾�*��T@V��G,����   �   2ߒ�zit���i������Դ������?�|Ҋ���ľ܅���4��si�)W�����ʿ,�Uj���N��O���n����?⿚�ɿN&���1��^�i�.�5����ǾY����H�����$Ͻɹ�������Ý������߽X(	��%�1C�0n_��Ox�������������މ�h��
�n���R��;4�d����K��   �   I�j�3�rwB��A�����N��؍R������ ۾rH��J��N������}¿��Z���B	��,�V~����`��J`��67�و¿)k��r炿��K� #�-n߾�����3^�(T�<�ٽ`���]X������⍽*]��-�ǽ�H?�����K/�<�H�C�'�D��@�4$5�q%�wG�f����-ʽf�����z��   �   �	��p��(���w�}���89���a��������F�#�v�Z��猿�����ѿ�\�r��\�������8���=�@��B���ҿ=믿X���Z�\��.&�B>����;Wo�K�$��j����T�|���_�"Pc���~��+��v����[˽�潷��|����X��G�m���U�罒:ʽ©����?V��V&��   �   |	ɼ��ۼR��wt���ĽQ��*�k�S���<%����+��?e�/���T��O�ۿ����$�\��J�#��}&���#�n���'��b���ܿj�������0h�}�.�DU��?\���pz��i+���xJ����r���J�n�B�C�Q���o��X��@'�����$5Žd�ѽTIؽzؽ,�нH�½@E��@g���z��F��/�VW��   �   J7��ec����xc.����8I󽻜;�p⊾L�ƾ�X	�>�7��7m�`���כ���7ο@��ۇ��b1��h��2��������@�ο�d����ҟo�0�:���C_ξ�9��x�Q�f���ҽn�����u��U�RM���T���f���|����������������.Ѣ������� u���q��I�H��f%�h0����a��   �   `����ɼ�t/�zᔽ�T�o9��׈���þ�6��4�~�i��w��s⮿u˿���I���h$��O�� �����0�,�˿���o`����k�y7��Y
�˾Z摾��N�~��*�н~ؚ�8w�YZ�*�T�Y�_���t�H������2k���T�������E��گ�(���n��\k����d��V7��
�T�Ƽ2݋��   �   ���xH���I�c 3�l쑽n��~v1�=肾�ź���Dz,���^�SΊ�d񦿢����ٿ�j��b��u���A��0B쿝�ٿ�¿Y���r��6z`�9�.�h���w���&����E�a��p�ɽPӘ��{�ݱg���k�]��������a��`���ȽWb׽F��E��#r�k5ڽwhʽ� ������P���H����L�ݼ�   �   a� �������:�b
���F۽��%��Qs����:��j��M�V��7r��ix���ɿ��ڿ����|�3���kڿu)ɿ�D���y��d�����N�b� �������ɣ��\F7�����1��L�������	*��9>���R��3�ӽe��Y���:��&��$��t���������⽜@��i��6n�Ԓ4��   �   HY�߬1��)���H�̅��w(̽@H�0 \�����/4־9��pR8���e�Nj����sȴ��IĿpο�Xѿ��ͿC�ÿ�"��yc������e��8�܌���ؾ����h�f�Z%��ｵ�� ��E���EM�����֨Ƚ���˭���#���8��5K���X�ݺ`�+�a��[�wO�֍<��%�z����1ζ�)匽�   �   �*����{��UY��^��ֈ�Ρ���e��B��U�������;�����0pG��@p���!��#�������޵�����F٩�2��;芿��n�leF��]�y���z���\���H�Rq��׽ׁ��%H���ޙ��ݮ��6ӽ/�������>��_���~�w'����������g������c-��,�����m�-9K�:�'�@C�i�н�   �   ��Jr��H닽V$�pl��Į��Iｄ�'�`�h�~F����Ѿ����'�5�I���j�����v������C�a1�����������h���G���%��=�d�Ͼo(��мh��#*�"a���9���K���m���宽�PԽ"��[�(�R�M<�0���?y���S��)�о�;ھ�ܾj(ؾ��̾�a��쥾�����k�%O=����   �   �|�F
转@��迕�dr��V��8�ҽx��zB�d��E���oܾ���R{$��>?�f�V��vi�u���x��3t�J�g�2�T���<��!�xG�w�׾�@��or��>�np��Խ��������K���˽@M�m7)�f�Y�*��6+��UkȾ.�羯���o�s+�
*�>3���
�����{�ྋ������|���� I��   �   g=I����4���������~����꺽������/T�>I��wǯ�v'پ��d���h)���7���@��C�,@�6�;�&����������ҾaQ���1��@:I�n����������⒞�}캽������!3T�fK��Fʯ��*پ������k)���7���@�&�C�R@�6���&���������ҾT���3���   �   �u�
>�(r��Խ��������,����˽eK��4)���Y����9(���gȾ���L��Zm��(�I'��0���
����\��������&���I��y�S�>��l���r���V��"�ҽ&�� }B�0�FH���rܾ����}$��A?���V�^zi��!u�L�x�t7t���g�:�T���<�R�!�\I�z�׾BC���   �   C*��u�h��%*�~c���:���K��?m���㮽�MԽ���e�(�<R�x7�B����u���O����о'7ھ��ܾ$ؾ��̾�]���襾�����k�EK=����o��"鋽("�^l��Ů�0L�]�'�"�h�nH��5�Ѿ����'���I���j����bx��m��� ���33��n��������h�%�G���%�G?�؄Ͼ�   �   �{���]����H��r�l�׽K����G��Aݙ�@ۮ�$3ӽ�������>���_���~�w$��q���z����c��E���'*��4���=�m��4K�p�'�,@���н�&��U�{�^RY�y�^��ֈ�����f��B�fW������{>��U��RrG�ZCp�ċ����ᓪ�����ൿ����ک��3���銿8�n�fgF�9_������   �   ~�ؾ̞���f�.[%�m��B���~��a����K������Z�Ƚ����?�#��8�1K���X�ĵ`���a��[���N�b�<�	�%�	��F��tɶ�nጽ�Y��1���)�ĖH�*����)̽kI�\�%Û�6־{��T8���e�}k�����ɴ�{KĿο?ZѿW�Ϳεÿ"$���d�������e�X�8�����   �   �����v���EG7�D��=2��J����߂��(��o<��m����� �ӽ���V���Ќ���������\��|�W�⽺;���d��4/n�c�4�_�t���0���:��
���G۽��%�NSs����۶�/k�h�M��V��7s���y��Q�ɿ&�ڿa��E~鿑��/mڿ�*ɿ�E��}z��!�����N�L� ��   �   ܻ�Dx��8'��9�E������ɽTӘ�a�{�[�g�*�k���������-_��2����Ƚ@^׽߃Ὣ��wm��0ڽdʽ����
~�������H�8��@�ݼ����D���G�R 3��쑽m��Rw1��肾�ƺ�>�{,��^��Ί�"�y����ٿ�k��c��v���B��C�r�ٿ�¿�Y��xs��{`�ت.��   �   �Y
�O˾�摾��N����N�нtؚ��7w�uZ���T���_�e�t�����&��Mi���R�������C���ׯ��%���l��Ri���d�MS7�_�
���Ƽ�ً��`����T�ɼ�t/��ᔽ\U��9��׈�P�þB7���4��i�Zx���⮿�˿ �ҩ���$��O�� �Y���i1俇�˿V����`���k�dy7��   �   ��_ξ�9��Q�Q�J���ҽL�����u�ͳU��QM�[�T���f���|�G��J���|��������Т����S����t��Gq��I�!��$%�F0��l�a�8J7�,fc�~����c.�F����I���;��⊾~�ƾ�X	�d�7��7m�v����8οS�����f1��h��2��������1�ο~d������o��:��   �   lY
�v˾�呾�N���Z�н�ך�k6w�~Z�
�T���_���t��������i��vR��^���pC���ׯ��%���l��Ii����d�ES7�2�
���ƼZً��`����ɼ�s/�ᔽDT�39�c׈���þ�6���4�,�i��w��1⮿"˿,��٨��*$�lO�^ �[���}0俳�˿����`���k��x7��   �   º��v��&����E������ɽ�ј��{���g���k���������^��������Ƚ�]׽���v��Nm㽶0ڽ�cʽ�����}��Ͷ�k�H�����ݼ`��RC��bE�l3�t둽Y���u1��炾 ź�0��y,�5�^��͊�������;�ٿj��a��t���@��9A쿳�ٿ¿[X��Qr��(y`�b�.��   �   ���Մ��ڢ���D7�����/��U���hނ��'��N;��t���0��`�ӽ��V������l��g��Έ�K��p�;�⽚;���d���.n�݌4������e���:�����D۽o�%�HPs������;i���M�WU��]q��lw���ɿ��ڿ���~{�ԋ忓jڿ5(ɿ�C���x������A�N�G� ��   �   ��ؾ$���6�f�fX%�Y��1��}|������J��7���)�Ƚ��}����#���8��0K���X���`���a��[���N�S�<���%������Bɶ� ጽ�Y�{�1���)���H�̃��=&̽�F�j�[������2־%��Q8��e�Bi��d�Ǵ�aHĿ�ο�Vѿ�Ϳ��ÿ<!��!b������e�D�8�����   �   �w��[����H�vo��׽�~��$E��.ۙ��ٮ��1ӽ;��5����>��_�B�~�T$��V���e����c��9���*��.���0�m��4K�Z�'�@�:�н~&��ò{�PY���^�;Ԉ�*���d��B��T��診�p9����CnG�}>p�;������z���;��ݵ�ꫲ��ש�q0���抿M�n�FcF��[������   �   Y&����h��!*�>]��^6���H���j���ᮽ�KԽ6����(�� R��6�����u���O��ݺо7ھ��ܾ�#ؾ��̾�]���襾����k�,K=������7n���狽���i��*����F�[�'���h��D��"�ѾY���'���I�(�j�k���t��ɡ��m𘿏/������X
����h�.�G���%��;��Ͼ�   �   xn��>�n��Խ"���-��������˽�J�4)�%�Y�����'���gȾʜ�<��Nm��(�D'��0���
����X�������������I��y����<������ho���R����ҽJ}��wB��wC���lܾ���	y$�P<?�e�V��si��u�5�x�|0t��g��T�7�<���!�tE�3�׾^>���   �   �6I�������P������b����躽˞����R/T��H��;ǯ�C'پ��S���h)���7���@��C�*@�6�;�&��������}�ҾVQ���1��:I�����y������\���o纽x�����,T�G���į�$پ�����&f)���7���@���C��?�6�t�&���V����ҾxN��d/���   �   �v�Y��9����n��AS���ҽ�~��yB�񂾜E���oܾ���@{$��>?�\�V��vi�u���x��3t�K�g�2�T���<��!�tG�l�׾�@��Ar�?>��o�TԽz���v��������˽�H��1)��Y�`��C%��&dȾϘ�����j�&��$��-�m�
�\���$��a�����������&I��   �   �⽻j���勽��Hi������2H�ԋ'�׾h�DF��h�Ѿگ��'�(�I���j�����v������D�a1�����������h���G���%��=�Y�Ͼ^(����h��#*��_���7��I��/j��X஽]IԽT��"�(�-�Q��2�T�pr��L��Ҷо�2ھ%�ܾ�ؾ^�̾)Z��A奾����k�,G=�ƽ��   �   �"��<�{�LLY���^�Ԉ�⟼��d�SB��U�������;�����#pG��@p��� ��#�������޵�����G٩�2��;芿��n�keF��]�p����y��~\����H��p���׽���E��;ڙ��׮��.ӽ2�����>�߈_�J�~�!��9������(`��⯛��&��:�����m��/K�~�'��<�8�н�   �   ��X�H�1���)�/�H�̃���&̽�G���[�����4־,��fR8���e�Kj����qȴ��IĿqο�Xѿ��ͿE�ÿ�"��yc������e��8�ڌ���ؾ����0�f��Y%������|��屢��H�����-�Ƚ�������#��8��,K���X�İ`��a� �[���N��<��%����K��yĶ�Q݌��   �   U����m���:�����E۽�%�`Qs�c�� ��j���M�	V��5r��jx���ɿ��ڿ����|�4���kڿu)ɿ�D���y��d�����N�a� �����������F7�T���0������ ނ��&���9��a���g ��Զӽ��,T���t�������b����b����⽿6���`���'n�n�4��   �   ����\?���B��3�x둽���:v1�$肾�ź���>z,���^�QΊ�c񦿢����ٿ�j��b��u���A��1B쿝�ٿ�¿Y���r��5z`�8�.�e���w���&��u�E�$����ɽ4Ҙ���{���g���k�Ƌ��D���{\�������Ƚ^Z׽��M��i�u,ڽ�_ʽ����}z�����,�H�����yݼ�   �   �`������ɼXs/�����ST�N9��׈���þ�6���4�{�i��w��s⮿t˿���I���h$��O�� �����0�+�˿
���n`����k�y7��Y
�˾T摾��N�_��Ӌн�ך�z6w�.Z�d�T���_�T�t���������g���P�������A���կ��#���j��~g����d�dP7���
�f�Ƽ�Ջ��   �    -�����D�p�߼P�T�/c�������S�i���j�Ѿ�%�>(5�z1b��W�����色�' ¿�̿H�Ͽ�̿C/¿���s��!��c��t7�>�5�پMj���io�On0����k,̽%����t��>���d���m��@q������"������۔��(��`������s	q�#T�~2����D�м0C���(��倻�   �   ��z�@���<�R��X⼯nS�\���/�P��f��	tξ��	�
S2���^��6��B��0į�����ȿ�F̿��ȿ��g䯿"���=����-`��x4�i��
[־�ӟ�ѩk���-��� �ɽ�2�����`x�� c��|Ċ�^=��r
��t��5n��U���y����4���	��Zl���m�5�I�d#��N��4ѩ�<�N�p�ػ�   �   �!%�ذ"������4EP��������H��玾5ž>��!*��YT����.��#���#S��������¿̒��R7��릧�-���S���uU�`�+��*��*̾eR����`���%����E½R2���W���������)�����0���9J���G��\���F½˿����)�������["d��4�(\��й�Hhq��   �   z쩼�C������|�����L����Q�����:�nτ�	Ӷ����A��=D��l�zǉ�[��1��� %��T
�������E������������l�ܹD��P��N���I��\���M�O�#��s轴[��֬�����`����V�������#����˽W�ݽw�����j� �p�D����u�ڬ޽�Uƽ���������Z��M#�"��   �   s���fR�(�7�J��9���*轝�)��9p�������ھq����/���S���v�̊�m薿헞�a%���X���{���N��:�u��1S��|/�&7���ܾ],��@~{��&:�[R
��ӽHk����,���v"��Ὣ���ýa�Ǧ���Y�+�Q�'���/��A3�4�1�nq+�� ����_�����ӽCͪ�;�����F��   �   �Gh��3������!�eM������=ҽ<!�E�S�pt���-��z������7��U�жp��ւ�Qz��r���*���F���Jo�szT��m6�b����󼾾����1�Y�4�!��/���@B������.������ƽ�������"���9���O��b�dep�5�w��Wx��'q���b�GhN���5�2N�1!��dxȽ_ؙ��   �   F���RZ��x�P���@�h�U�!��2���z�#37�~w������ϾF� �r���3�,2J�"�[��f�:Fj���e�QJZ��RH���1�O���c���̾���V�s��6�o�D�ν@W�������/��Ą��R|��#�����/�HQ�Ws�%找���٢�7���q���K��H������A�}�X�X�kL3����-�޽�   �   �a꽬���C���j��&f��ք��	��B~� ���O��t��vϫ���Ӿ�Y�����ʮ$�c�2��~;�7;>��:�� 1��Q"��������,;�I���q��&�E����*�߽����Đ�
#��J�������n�߽pY�{3�?^�I2�������X&ɾ��ؾy`⾇����߾��Ӿ�	¾٫�fE��Hft�+�D�݋��   �   *�o��i��Q���3��j���ZE���ɽ<��?�,��]��!�����l-ʾX0龥T�L���)�����V�`������1���p젾ܡ����J�~'�����������n��b���7F��pɽ�����,�;�]�$������0ʾ4��V������������
��������X�������	 K��   �   ��E�����߽����Ő�\#��ɫ��@�����߽�W�dx3��^�0��������"ɾ��ؾ^\�[�侼�߾��Ӿ1¾�ի��B���at���D����']�h}������j��%f��ք��
�������>�O��v���ѫ���Ӿz]�����+�$���2���;��=>���:�e1�2T"���������/;�K���s���   �   8�s�D�6��p�g�ν�X��,����/��Ƀ��dz��)����P�/��DQ��Rs��㉾�	���բ��3��on��0H��
������}���X��H3��}�X�޽�|���W����P���@�؜U��!���3��4|�#57��w������Ͼ�� �`��O�3��4J�߱[�˽f�Ij���e��LZ�
UH���1�*���f��
̾�����   �   ���L�Y���!��1����B�����.��������ƽ��Ȍ��"���9���O���b�{`p��w�JRx�["q���b��cN��5��J�6��}sȽrԙ��Ah���3�����!�KM�f���K?ҽ�"�U�S��u���/���|�������7�F�U�V�p�N؂��{��ߧ��{+��HH��3Mo��|T��o6������Ҿ���   �   �-��*�{�0(:�ZS
��	ӽl��X���ߑ��!��C�����ý�]འ���W�(��'��/��=3�<�1��m+�$
 �H��$�����ӽ�Ȫ�n����F�����N�.�z�J�y:��n,���)��;p�
�����ھ���t�/�b�S���v�3͊��閿<����&���Y��'}���O��0�u�x3S�<~/�B8�w�ܾ�   �   �J��%���p�O������h\��'������̃���U��K���L!����˽��ݽ9��A���ʱ �Xm�����p񽆧޽�Pƽe �����4�Z��G#�:��婼�>������T���!�L����Х���:�MЄ�@Զ�����B��>D���l�]ȉ�W��?���6&��n�������F������R����l��D��Q�
P���   �   k+̾�R��t�`�;�%����jF½�2���W��(��ζ��(��V��8����G�� E��2����B½oǿ�e��������ܦ���d��4��W�^ɹ�`\q�%���"�L��Z�꼺EP�6�������H�1莾6žޭ��*��ZT������ݱ���S��^���c�¿����
8�������-��RT���vU��+�I+��   �   \[־4ԟ�-�k�ż-���f�ɽ�2�����,x���b���Ê��<��\	��&���l�����������2�����|j��#m���I�d#��I���̩�ЄN���ػ�uz�X�����R��X�)oS��\��|���P�g���tξH�	��S2� �^��6��cB���į�����ȿNG̿G�ȿ{���䯿i���w���.`�'y4�����   �   �پ7j���io�<n0����Z,̽���kt��"����c���m��
q��b����!��`��D۔��(�����I��	q��"T��}2����ހм�B��(� 倻�,����TD���߼��T�qc����:�S�������Ѿ�%�^(5��1b��W���������3 ¿�̿K�Ͽ�̿=/¿���h����c��t7��=��   �   wZ־�ӟ�-�k��-�%�s�ɽ 2��>���w��.b��XÊ�<��������`l��a���w����2�����^j���m���I�F#��I��f̩�<�N���ػ�qz�0�����R��V��mS��[������P�uf���sξ��	��R2�8�^�o6���A���ï�Y����ȿ{F̿y�ȿ���䯿Ŏ��鹆�0-`�gx4�	���   �   �)̾�Q����`���%�����D½1��V���������'��l��c���G��dD������1B½ǿ����T�ߨ������Qd���4�zW��ȹ��Zq��%�ħ"� ��>��}CP�����u���H�玾i4žʬ��*�8YT����������sR��է����¿����6��3���c,��BS���tU���+�**��   �   BH��b�����O�������Y��������#���T��鬧�	 ����˽��ݽ[������� �m�E����o�K�޽�Pƽ8 ������Z��G#�(�J䩼�<�����������L�D��|�����:��΄�Ҷ�·�A�w<D�ʚl��Ɖ�x��6���$��A	�������D�����������l���D��O��L���   �   �*���{{�	%:��P
�"ӽ
i������ݑ����r�����ý=\�<���mV��'���'���/��=3��1�]m+�
 �.������[�ӽvȪ�3���G�F��
�\�xJ㼏���J��7��o(�!�)��7p�^���6�ھ]����/���S���v��ʊ�?疿����$��;W���z���M��"�u��/S�N{/��5�Ȯܾ�   �   ������Y�G�!�,�����?������+��������ƽ�����"���9�(�O��b�`p���w�Rx�0"q���b��cN�ӓ5��J���@sȽ ԙ��@h�4�3����'�!�M�R����:ҽ���S� s���+���w��n����7���U�r�p��Ղ��x��	����(���E��FHo�1xT��k6����p��ں���   �   �s���6�m���νXT�������,��G���.x��#�����y�/��CQ�Rs�R㉾�	���բ��3��Vn��H��
����� �}���X��H3��}� �޽|���V����P���@�x�U�`���.��y��07�{w�����Ͼ�� ������3��/J�~�[�$�f�`Cj���e��GZ�PH�q�1�[���`���̾�����   �   
�E�}��<�߽@������ �� ���������߽�V��w3��^��/�����W𴾒"ɾ��ؾ@\�E�侪�߾��Ӿ&¾�ի��B���at�i�D�Ԉ��\꽼|������j�k!f��ӄ����yz潰����O��r��ͫ� �ӾZV��y��z�$�ޭ2�:|;��8>�>�:�K�0��O"�l��W����);!G���o���   �   �$�$����_���}��N����B��WɽC��_�,�O�]��!�����'-ʾ 0龏T�=�s��!�����R�Y������)���f젾Ρ����J�I'������H����������1B���ɽ���o,���]����D��;*ʾ�,龏R���������
�"���-������頾����#�J��   �   X�Vy���
���j��f��ӄ�z��N|�.����O�tt��*ϫ���Ӿ�Y��o����$�X�2��~;�1;>��:�� 1��Q"���������,;�I���q����E����d�߽g��Ð�� ������������߽�T�;u3��^��-��*��g�4ɾ��ؾIX�2�侠�߾��Ӿ�¾�ҫ��?��]t���D�څ��   �   >x��T����P�^�@�y�U����0��z�p27�j}w�����L�Ͼ*� �\����3�!2J��[��f�8Fj���e�PJZ��RH���1�L���c���̾
���4�s���6��n�R�ν�U��z����,�������v��������/��@Q�!Ns���������Ң�t0��k���D������|��Ӥ}�P�X��D3��z��޽�   �   �:h���3�t��U�!�{M�����<ҽ� ���S�0t���-���y��׳���7���U�ɶp��ւ�Pz��r���*���F���Jo�qzT��m6�^����缾������Y���!��.�|���@��)��H+��x���ܷƽ�
�����"���9���O��{b��[p���w�Mx�'q���b�_N�ʏ5�G���MnȽ*Й��   �   >��켺E�6�]�J�8���)��)�,9p�t�����ھa����/���S���v�̊�l薿헞�c%���X���{���N��9�u��1S��|/�#7���ܾT,��"~{��&:�R
��ӽ�i��1���ݑ����0�����ý�Y཭���2T��$�r�'�E�/��93�J�1��i+�p ��~�����
�ӽ�ê�p|��4�F��   �   �ݩ��7��^���D���ײL����f���^�:�Eτ��Ҷ�����A��=D��l�xǉ�Z��0���%��U
�������E������������l�ڹD��P��N���I��P���*�O������Z��y������́��YS������2���˽��ݽ���U���&� ��j�����j�I�޽�Kƽ����"���h�Z�0B#�j���   �   <%�8�"������hCP�͚�����UH�h玾�4ž5��*��YT����-��$���#S��������¿Β��S7��릧�
-���S���uU�`�+��*��*̾]R����`���%����PE½s1���V�����N���N&��Z
������GE��+B�����P?½Ŀ�񲸽ꬽ¥��̣���d��4�fS�¹��Oq��   �   �`z�𥲻d�R�.V��mS��[�����P��f���sξ��	�S2���^��6��B��/į�����ȿ�F̿��ȿ��h䯿"���<����-`��x4�g��[־�ӟ�ũk�q�-�o�ܖɽ^2��Z���w��b��Ê��;��_����rk��M���6���&1��L���h��"m��I��#�E���ȩ��}N�h~ػ�   �   ���;�'�;�D���k�}
���}���νjV��`��\���^Ͼ\��%-'�$�I��ak�����h��������:����r��{Ä���k���J�`�(�
����׾92�������G��`��p��J�3ͽ�sĽ&���i���ɋ���ܿ��������"����࠽J����pl��K��'����\b����k��Kػ ��;�   �   hL�; �I; hA��5r��E
���{�d9̽�L��]�����B̾��>�$��F�%�g�X���������n��↕��!��ğ��+h�@�G��;&�Nt�3Ծ����*}���C� ��� ��A)ݽ߽ʽ��½!������P�½�½�6��Sع���� 5���a���ю��d�S4^�G`:�����ݼ�$�����+6�`�;�   �   @W2�@gB�x�������
�qu��\Ž u��T�ܚ��YFþ���x��p=���\���x�.{��'���d�y���e��J�x��]��
>��C� �vʾ?��Pq���:����x��c/ԽZ�ýPώ�W��Z����ƽ!$ɽ�.ʽ��Ƚ?Ž�ƾ���������m����b��G�s�~�J��X �$ 켪���<.0�8����   �   �]���P?#�����&U�f�l�U�����F������_���K��K�D/�)L���e�J+z�'���u���*p��׽y�Bee���K��/����?��_��������^��,����;L��ƽ������u����ý~1ͽ_Xֽ� ޽"��{�sQ�Ƙ���ڽ_Ͻ^���"������u�HB��N�:Ǽ<m|��   �   �a���ȉ�v]��4�������%d���2� ���5��x�����"Ҿ@������6���M�߷_��5k�Po���j���^��L���5��7��� �Ҿlm���:���&G��b��_��`̽�õ�B���a�������Ƚi�ٽ���a������i�޿�5���U���^����.,ؽ"��(#���To�qX3��P ��   �   S��d�򼺍Ӽ��漰�c^�lR꽙0#���\�����c����0��R��h2���A�x�K�:�N�VK���@���0���Q��R��
���鏾W�_��R,�Լ���ս$��D٣�*���0����ѻ��	ӽ7+�V�������"���/���9���@�W�B��?�k8�23+�oB��c�����������}�V��   �   I u�/�;��`�X��9')�Y]�У��T�ӽ6��U�@��pz��1��mT¾��a��<�c�"���*��_-�p*��U!�n��Y������Y����p��;�&0�e>ཞ���v}��H��������p��Ե½����)����6�2�IxI�=�^�WHp��#}��ׁ�7~��۽z�]k���U�C<�=0 �����ѽ�ҡ��   �   q�������*V�6�<��A�c�"����+��� ��M'��U�e��t;��x�����ܾ6��t�#8�I���
�����Y�Ծ^춾�c���v���B��0�o���ȵ�r���2��� Ճ�F+��N��QнS������܊9�(-Z� /{�:��|ǚ�N��^誾.����H��֝�,/����~��IZ���4��|�˜��   �   �뽵ƴ��=��Bo��1a�$4q�����D�����t-��5���^�Tz���(���豾�ž��Ӿ��ܾ�޾
�پY'ξǼ�9Q��������n�A�j��뽊ô��;���>o�=/a�3q�����E��M���.�,�5�P�^�$|���*��p뱾�	ž�Ӿ�ܾ��޾��پ�*ξ#ʼ��S��Y�����n�;A����   �   3���轐˵�m��������Ճ��+�����н���E����9�&*Z�B+{��7���Ě����e媾"����E��*ӝ��,��J�~��EZ�%�4� z�@��آ��	���&V�=�<��A�~c�����$-��� �LO'�n�U��f���=�����ܾ�9��V�:�N��� 
����C�d�Ծ��e����v���B��   �   �;��1�"Aེ�����P�������p���½�你(�����2�JuI��~^�6Dp�@}�"Ձ��{����z�TXk�^�U�!?<��, �ʾ�$�ѽ�Ρ�*u�r�;�T]� ��
&)�`]�������ӽ}��;�@�*sz�|3���V¾�����>�g�"���*��a-��*��W!�@�}[����J���[����p��   �   ��_��T,�-����ս���jڣ�䰡�f����ѻ��ӽg)�������g�"��/�j�9�~@���B�'�?��8��/+��>��`�.��R ��Φ��4�V�M����� �Ӽ�����^�P��1#���\���d��侙������i2���A���K�_�N�pK���@���0�7����������c돾�   �   �;��9(G��c��a���a̽�ĵ�����������Ƚ,�ٽ��뽰�����g�r������R���p��G���&ؽX������SMo�[R3�L ��Y����LY��Μ��T��U&d���� ��5�� x�����#ҾZ����6�~�M���_��7k�Lo���j���^���L�b�5��8�����Ҿ�n���   �   b�����^��,�U���M��ƽƊ��<��������ý�0ͽ	Wֽ�ݽ���x��M�����ڽ Ͻ$�������"�u�"B�7I�4Ǽ�^|��R�h�9#�t���'U�H�l�B��ӎ�D�F������`��dM��L�i/�}L��e��,z�����J����p��\�y��fe���K�
!/�������`���   �   ���Qq�[�:����t��*0Խ��ý�ώX��.���Zƽ<#ɽa-ʽ>�Ƚ@Žgľ� ����������_���s�m�J� T ��켖ٜ�P"0�ȑ����1��B�0������
��qu��]Ž�u��T�����?Gþ8���2��q=���\���x��{�����𐿥y��ff��G�x�_]��>�BD�� �9ʾ�   �    ����*}�
�C�q��C���)ݽ6�ʽ��½2��������½t½!6��\׹�����3��`��*Ў��a�T1^�h]:���
ݼ< ��x�P6�P�;�T�; �I;�aA�45r��E
�G�{��9̽:M���]���7C̾d����$���F���g����� ��U������1����!�����z+h���G�I<&��t�b3Ծ�   �   *2������zG��`��p��J�3ͽ�sĽ���F��������ܿ�\����������R࠽���z�col�K���'�Q���a����k�@Iػ ��x�;� �;(�;�D���k�C}
�7�}���ν�V�H�`��\���^Ͼu��@-'�@�I��ak������h����󋚿:����r��vÄ���k���J�Q�(������׾�   �   Q���s)}�4�C���� ���(ݽL�ʽڴ½Y������:�½�½s5���ֹ���@3���_���ώ�{a��0^�]:�϶��ݼ������6� �;pV�;`�I;�ZA��2r�E
��{�9̽�L���]�g��aB̾����$���F�ūg� ����������"������:!��z����*h�ŚG��;&��s�2Ծ�   �   �����Oq���:�8��H��<.Խ.�ý�߽�zV�������ƽ�!ɽ,ʽ�ȽEŽ�þ�r�i���.����_��]�s���J��S �`��؜�� 0����� �1� �A��	�������
�Xou��[Ž^t�B�T�U����Eþ,�����6p=��\���x��z�������yx��Je��8�x��]�
>��B�p ��ʾ�   �   ����'�^���,�����J�Y�ƽH������F���j�ý�.ͽUֽA�ݽ�㽥v��L�����ڽ�Ͻ���*��� ����u��B��H�dǼ�\|��O���4#�
}���R���l����	����F�ב���^���J�"K�C/��L�N�e��)z�]�������[o��F�y��ce�0�K��/����� 쾤^���   �   �9���$G�Da��]���]̽�������������i�Ƚ��ٽ��뽔�����f�ļ�����R����+����&ؽ�������Lo��Q3�wK �JX������TV������K���!d� ��� ��5��x�~���\ Ҿ<�����6� �M��_��3k�_o��j���^�4�L�[�5�(6���&�Ҿ�k���   �   ܒ_��P,�>���ս����֣�����B����λ��ӽ�&�����b�"��/���9��}@��B���?�F8�I/+��>��`���� ��������V���\��քӼ`�漞�^��뢽U��.#�`�\����7a��s	�ָ����Qf2���A�h�K��N�>	K���@��0�����������`菾�   �    ;�%.�;�Ĕ���z����������Tm���½��B'������2�CtI��}^�~Cp��}��ԁ��{����z�Xk�3�U��><��, ����ݛѽ]Ρ�Ju�E�;��[�����")�h
]����
�ӽ9����@�pmz��/��R¾N����;�l�"���*��]-�T*��S!����6X� �ᾖ���W��s�p��   �   y.���轢ŵ�����r���P҃�3(���
��#нS������Z�9�)Z�J*{�u7���Ě�:��.媾�����E��ӝ�w,��)�~��EZ��4��y���p������%V���<��	A��c�-���{(��� �K'���U�(c��39�������ܾ�2���	�(6�F���
�.��R �6�Ծ�鶾9a��P�v���B��   �   N	�ڿ��h8���8o��)a�\-q����B��ݤ�.,��5�l�^��y��+(��m豾yž��Ӿ[�ܾ��޾��پD'ξǼ�+Q��򛏾��n��A�E�n�ô��:��r<o�#,a��.q����vA�����+�3�5��^�>x��(&���屾�ža�Ӿ��ܾk�޾z�پ�#ξ�ü�jN��������n��A����   �   Ӟ������ V���<��A��c�`���^)��x �{L'���U��d��;�������ܾ�5��\�8�=���
�����M�ԾR춾uc����v���B��0����Hȵ�����ԃ��(Ӄ��(��~
��6н�������b�9�o&Z��&{�m5��<�����X⪾����B��EН��)��~�~��AZ���4�w�]���   �   9u���;�2X�<��A!)�
]�w���)�ӽ6��d�@��oz�U1��T¾���C��<�S�"���*��_-�j*��U!�i��Y�۹�����Y����p��;��/��=�ٖ��S|������<���hm����½ϙ�>&�O����2��qI��z^��?p�t}��ҁ�6y����z��Sk���U�*;<�f) �ѻ�"�ѽ�ʡ��   �   �����RӼʯ漭�
^�|좽���/#���\�6����b��o���>��	h2���A�o�K�4�N�RK���@���0���N��H��
���鏾9�_��R,������ս<���ף�H�������zλ��ӽU%����n�"���/���9�Oz@���B�*�?���7��++��;��]���Ὄ�������X�V��   �   �P��躉�(R��ޕ�����+"d������ ��5�hx������!Ҿ(����u�6���M�ط_��5k�Mo���j���^��L���5��7�����Ҿcm���:���&G��b�y_��R_̽�µ�э��\������Ƚ��ٽJ�뽇�����e��������O���z�����!ؽ��������Eo�L3��F ��   �   4E�h�.#�,{��ER���l�4�������F�q���k_���K��K�6/� L���e�G+z�&���t���*p��׽y�Aee���K��/����:��_��������^�Ď,�X���K�H�ƽ����W������X�ý7.ͽFTֽ��ݽL��Yt�J�ː⽔�ڽ�Ͻ�
�����\���N�u�B��C�$Ǽ�N|��   �    R1� �A����x����
��ou� \Ž�t�ȺT�����<Fþ����o��p=���\���x�.{��'���c�y���e��J�x�]��
>��C� �rʾ9��Pq���:����)���.Խ��ý_ཽ�V�������ƽy!ɽr+ʽ#�Ƚ�Ž������R�������J]��߄s���J��O �8��Ҝ��0��}���   �   x\�;P�I;@SA�X1r��D
�߰{�9̽�L��]�����B̾��8�$���F�"�g�X���������n��㆕��!��ğ��+h�@�G��;&�Mt�3Ծ����*}���C���� ��	)ݽ��ʽ�½����6���C�½�½N5��~ֹ�����2��
_��ώ��_�/^�0[:����(ݼ���p���5���;�   �   ��G<��.<���;�]���d��_�(����E�߽�8"��[`��`���G����qi�
k(�t�=��N�&�Y�̅]���Y���N�0$>��)�������FjȾ�ڡ�J���KT�V'2��h�9��|������L��Z���{�>���|G��C�ὦ*Ƚ���<(����r�S�A�$��T�ͼ|�y��Ի��~:`��;HS/<�   �   L�0<`�<X�;�ҝ��b���5(�򞏽i�ݽU ��}]�}U��؂������2�4�%���:�K�K�IV�[�Y�~AV�T�K�8;��Z&��p�P��a0ž�C���7��6�P��W/�������jg
���v��
��~��F��]��B��r���γ�t7̽����|�����G�N�� �vZ�.��������� ��;\�<�   �   e�;�(�;�[
;��ջBI����'�;����E׽o��jDU�t��ƈ��y�����M0�812��B�r,L���O��L���A�x2�c�����ջ�h����bt��%G��('�-�����a�g_�#���z�.��T���߷��; �P���ؽ�T½����%^��v}w�F�H����4|޼����P�@ҿ�0�u;�   �    YD� B�9�"���ln��0(��و��ν��� �H�u���F����ѾE���qg��$�,3�wj<�\�?�>&<�n�2��&$�"��\���08Ӿ�=������a�J�7� N�����������1���B� �t��x 
�
]��k��
�ڳ�! ���ｏ޽��ʽ:��F���m��e^��.�؆���ܪ��vD����   �   ��7��`���m� �μ�+�&O����ý�Z	�Q�9���r���0佾�㾡�����k ��~(��+��(�؁��}��C��ྜྷ�������,%z��sI�N$$�y�	����&U⽔�޽X�dVｱ���ڪ�P�	��{��/���#��	� �����E��#ӽ(���q��z�����Q������ݼB����   �   ��ͼ�����󒼚I��RH���)4�����>I���L����)���Z��������#�ǾK��� ��r�u+�B9��b���	��I���6��E¾���s̅�BX��.����
�n>ҽَŽ|
Ž�ͽ�ܽ���Z �e	�D��+]����V!���"�c�!�<��k%��=�� ��⽠���֟�L[}��@�ԛ��   �   �,.���	�`���������C��ф�����;�ԃ���C��7r�P4������~�ľ��ھ��뾦t��+R��^"��`�IԾ������������_�%�4�/��	�a\ƽ?���駽 ��'z����ʽ�D����x�+���'��63�,�=�~[E�4�I���I�03E�l�;�{�-��V�r(�Љ彽'���ғ���c��   �   �ǁ���O�2�1���)�X�7���[��`��K���������;/��DT���{�'���0������h�¾S|ʾ�̾�<Ǿ�q�������E�����9]���4�$����鼽���i��w�����N��Gͼ��۽�/��1�'�V<��P��c�lKr�6�|�J�gi��Kv�ٚf��lQ�U\8�HR�^>���ѽ1����   �   e߲�rS��'-t�:`��c���|��̔�����\۽�������;�S�X�HWv�������p蝾�Ȣ�����n���L���^���xq�yaO��-����ܲ��P��s(t�6`�ޣc�1�|��˔����]۽"�����#
;���X�)Zv�y���	���Ꝿoˢ�(	��iq��TO��a���|q��dO��-����9"��   �   v�켽0�������y��*��u���ͼ�@�۽ /��z��}'�LT<���P��
c�Hr�d�|�:���$e��Gv�ǖf��hQ��X8�JO��;�=�ѽ�����ā���O��1�K�)���7��[�X`��^��i������</��FT���{�����2��,����¾ʾ�̾�?Ǿ@t�������G���	���<]�b�4�Z���   �   �0���_ƽbA���맽9"���{����ʽbE�����U��d'�&53��=��XE��I�t�I��/E���;��-��S��%�Ƅ�[#��=ϓ�u�c��'.���	�R�X�����@�C��ф������<�݄�a�C�:r��5��Z�����ľ0�ھ��뾠w��6U��X%���b羟KԾ�������̉��b�_�n�4��   �   U.�G���@ҽ�ŽHŽ}�ͽ0ܽ����Z ��d	���@\���� U!���"���!�����"�:;�T� ���� ���ҟ�T}��@�����ͼ����>HE��dE���(4�Ȁ���I��N����)�_�Z��������Ǿ[M�E� �0t��,��:�%d�I�	�,L��9ᾼG¾m���ͅ�DDX��   �   �uI��%$���	����W�U�޽�Y佪W､�����R�	��{��.���"�~	�3�����tA轤ӽ �m��ݧ��!�Q������ݼ����7������m�<�μ׍+�tO����ý�[	���9�]�r�=���彾w㾵��@��m ��(�+�1(�*���~��D����#���:���9'z��   �   �a�y�7�$O����_���`�������� ����� 
�]��k��
�,��Q���ĳ��޽ؕʽ(|��1���j��:_^��.�^}���Ԫ��hD� � �C� A�9 	����^m��E(�@ڈ��ν>���H��u���G��ͻѾ����_h��$�:-3��k<���?�l'<���2��'$�������t9Ӿ�>������   �   �ct��&G��)'����x�wb��_����Q{�h��T������T; �����ؽ�R½����\��>yw�(�H����u޼�����	�`���p�u;0r�;�3�;�k
;��ջ�H��ۑ'������F׽	��LEU��t������|�ᾋ��1�22��B�T-L�d�O�`L�w�A�22��c�z�����ջ�����   �   �7����P�YX/�f�����g
������<�����H��@��
���������u6̽m���O��������N�� �V�2��T�� ķ����;��<�0<$�<�;�Н��b���5(�?����ݽuU �0~]��U��X������.3���%�V�:�ŒK��IV���Y��AV���K��;�[&��p����0ž$D���   �   J���KT�j'2��h�X��&|���(��K��N���{�����	G�����,*Ƚ�����'��,�r���A�����ͼ��y���ӻ :���; T/<L�G< �.<(��;�]���d����(�2�����߽�8"�\`��`���G���ﾆi�k(���=��N�0�Y�Ӆ]���Y���N�-$>��)�������<jȾ�ڡ��   �   \7����P��W/����t��-g
�F� ���������������������,���5̽ᩲ�������M�N�# �dU缰���������0��;��<�0<`�<��;�̝�pa���4(������ݽ�T �I}]�GU��������뾘2���%���:��K��HV���Y�AV��K��;�cZ&�7p�����/ž{C���   �   �at�/%G�H('����H�Ka��^�n��%z�@��S�������t: �����ؽ�Q½����e[��7xw�[�H�+��t޼����p��x����u;pu�;p7�;Pw
;��ջ
F��ݏ'�:����D׽����CU��s��������o���/��02�)B��+L���O��L���A��2�hb�V����0Ի������   �   /�a�!�7�$M�ҩ������Z���4� �D��$�	��[�"j�0
����;��� ��z޽��ʽB{��t ��
j��f^^��.�D|���Ӫ��fD�� �C� ��9 ��l��\i��(�V؈��νp����H�Jt���E��G�Ѿ�����f��$�+3�Si<�0�?�%<�N�2��%$�1�������6Ӿ�<�����   �   >rI��"$�D�	�m��
S�b�޽�U佺Sｻ���/��s�	��y�P-��
�^!��|	�V�d���b@��ӽ]񺽝l��{���}�Q�i����ݼֲ��<�7�T�����m���μ�+�M����ýZY	���9���r�����⽾�㾔��ش�cj �4}(�@+�h (����M|��B������������#z��   �   �
.�+��T��;ҽi�Ž�Ž(�ͽ�ܽ}��X ��b	��}�yZ����S!���"��!����"��:��� �n�⽖����џ�vS}�c�@�����ͼ�����뒼�A��*@��.%4�8~��kF��EI����)�E�Z�������!�Ǿ�H澬� �[q��)��7�#a�m�	��F��k4ᾰC¾��˅��?X��   �   -�Q콁Yƽh<���槽���$w��+�ʽ A⽤�����b���'��33���=��WE�/�I���I�$/E�~�;���-�yS�^%�j��	#���Γ���c��&.���	��񼘾��e��u�C�(τ�񀳽�7��=�C��4r��2��j���!�ľ�ھ�뾤q��O��V��.]�\FԾH������]�����_���4��   �   �
��弽�	����Hu�����)���ɼ��۽�*����|'��R<��P��	c��Fr���|�῀��d�Gv�u�f��hQ��X8�O��;���ѽ8���tā���O���1�x�)��7�e�[��]�������ὺ���8/��AT�i�{� ��_.��H�����¾vyʾ�̾:Ǿ�n�� ����C����T6]���4�֘��   �   gز��M���"t��0`���c���|��Ȕ�����X۽���ü��;�ɮX��Uv�$��B��蝾�Ȣ�j���n���L���^���xq�SaO��-�����ὢ۲�*P��;'t�h4`�w�c�Ϲ|�Rɔ�a���X۽R������;���X�wSv����i���坾gƢ���Yl���J���\���tq��]O��-�������   �   �����O��1�_�)���7���[�B]�����2��P��:/�MCT���{����-0��j����¾|ʾ�̾�<Ǿzq��l����E������9]���4���|齞輽�����v��'��=��qʼ�U�۽�*���${'�6Q<�#�P�c��Cr��|������`�Cv���f��dQ�hU8�0L� 9���ѽ����   �   ".���	�6��z���w��.�C��΄�����8�l��x�C��6r��3������ľS�ھ���xt��R��A"���_��HԾ�����������_��4��.�C	��[ƽq>���觽@��jx��,�ʽ�A�ܡ��������
'�&23���=�KUE�x�I���I��+E�E�;���-��P��"������]˓��c��   �   ��ͼJ���f撼�=��R=��R$4�(~���F��:J��g�)���Z������ƬǾ�J��� ��r�d+�69��b���	��I���6ᾸE¾���f̅��AX�c.�����	��=ҽ%�Žv	Ž��ͽܽe��Y ��b	��}��Y���UR!���"��!������L8��~ ����J����͟��L}���@�?���   �   8�7������m�j�μ �+�-M���ý�Y	�t�9���r�����㽾]㾆�����k ��~(��+��(�ԁ��}��C��ྖ���򹚾%z��sI�2$$�U�	�:��T���޽�V��Tｸ��������	��y�-�
�� ��{	���-����<�*ӽ��-i��H�����Q�V��.�ݼ�����   �    C� {�9���X��
h��:(�m؈�_ν���b�H��t���F��H�Ѿ���^g���$�,3�oj<�X�?�:&<�l�2��&$� ��T���(8Ӿ�=�������a�8�7�N����P���P��o����� ������	��[�Fj�$
����D�����ｱ޽��ʽ�x������g���Y^�].�t��h̪�8ZD�ڦ��   �   8��; @�;p�
;��ջ.E����'�J����D׽��DU��s������X�����C0�012��B�o,L��O��L���A�v2�c����� ջ�c����bt��%G��('������a�+_�м��z���$T�&�����k: �-���ؽ�P½����Z��^uw�s�H�O���n޼��������;�� �u;�   �   �0<$�<���;0ʝ��`���4(�������ݽ�T �p}]�hU��Ƃ������2�0�%���:�J�K�IV�Z�Y�}AV�T�K�6;��Z&��p�N��^0ž�C���7��1�P��W/�������Vg
�r�N�����2������������=���5̽����������S�N�	 �BS缌 ����� ������;\ <�   �   ���<�r<��+< �/; ����Ӽ��D�l��� ~����R�F���p���ɾ�����2�ت��<����qH��������D;x��ێ���?y��}V�Xy?�^�3�b�1���6��AA�ЋM���X�!a�(d��a�N�W�I�� 6��} �}�	�[��L'��zᑽ��Z��:��mü4�E������;��7<�Ur<�   �   ��s<@a<��<�.�:�!��u׼{}E��P����!w�ٞP�Kl���:��<Aƾ:e�Y��l��LJ����@���������0�ɾ�:���4��,Hu�$S�p<���0���.��4��L>�7wJ���U�q^�>a��^���U���G��55��: �
����&���
k��g�b��"��Լ�;g�(Q���u;��<L|[<�   �   |M7<�,<��;�v��06A����h�G��Q��v�%� 0J�o���`���}���{ܾ8���c���j�9��6B�oM�EU���	ݾui������^����i�+*I�d�3���(�՝&���+���5�	�A���L�;!U�}�X�O"W��O�4C�*�2�,���h�e���Ž/t����{�4$=�P��������$�`Ժ�ƞ;0h<�   �   x$�;���;���:�o����z��y���M������ڽ���Ơ@� Ss��2�����z=;O�徔9����>��Bc������'侃�˾����;i��_���W��9�S�%�������T���Q(���3�L�>�ēG��KL�bL���F��)=�j�/����������Cֽs*��Qϓ���j�s�2�X������l�/��0W���;�   �   �p�� ]J�x:����4�LЩ�����Y������ֽ����5��cb�zi��sO���W��q�Ͼb`�Y�꾘��b���ݾ�˾�4�����FK��'d���@��%���q�
�\�	��[��b��"���-�0�6�I=�_(?�n�<�%�6���-��$"����@��(�Tҽ�����a��`�u���?�����uü�Gu����   �   �����b��.t�,Q��@3輾�'��l�-����Խ%7��*���P�I�y�	���趥�4I����ľ�0;�@Ͼ3�ʾ�D��ٽ��Oѝ�R���j�i:E�!S&����W����T�n��7M���g��_�T��0%%��--��&2�Y�3��r2��X.���'�-�� �:�
��-���n⽶�Žp}��v���m]�))��f���೼�   �   � �J�߼�޼�o���O� �K������^��2׽�$�f�!�0A�
b�ɔ��E?���Ԟ����
��>対x��������1����Wf��D��$�B�
��V�<Wӽ��ƽ��ƽ�Tн��ὢ���R�p���b��&��E-��^1��J3�3��0��
,���$�jz�M���o�<d�½�֠�:���=L�p���   �   mJ�	�1��5+�6�5���P���z��񘽾7���k��m�Cp���4���M�~Yf�]}������?~�����+w�����A>s�fX�@;�9��'���ݽ���7��w��1���CU���J���}ӽ�����:���e�*�Z#5���=���D���H���I��LG�j�@�@�5�}�'�o-����%޽ҷ�����s��   �   ���?}�ap���v��F���j���f��~�н#6�p�	��f��+-���>��N��b]���h�ap�4#r�`dn�`�d��dU���A���*����&���`v̽�@�����:}�Azp���v�9D��ch���d����н�4��	��f�,-��>���N��d]�m�h�Dp�e&r��gn���d�/hU���A�h�*�<������<z̽D���   �   ���*󧽅z�����W��qM���ӽ��x��,;�3�;�*��"5���=��D���H�h�I��IG���@�`�5���'��*�����ݽη�����s�
J�!�1�\1+���5���P�(�z�:𘽊6���j��m��p���4��M�c[f��}�h�����������y��v���As�X��
;����;����ݽ�   �   Z�IZӽq�ƽr�ƽrWн���>�����|��Rc��&��E-��^1��I3��3���0��,���$�x���zm��_��½�Ҡ�����KL�+��k| ���߼�޼�h��TL�T�K�����^���׽�$� �!�IA��b������@���֞�������H篾z��t��ු�Ғ���Zf�WD��$�"�
��   �   ���U���tW�>�� P��Fi�Wa����U&%��.-�4'2���3��r2�3X.�
�'��������
�*��k���Ž�y��튽R]��#)�]��8س�Nz����b�"t��K��R.���'�(l�Я���Խ�7��*�#�P��y�4���Z����J����ľ�2;�BϾ?�ʾ�F�������ҝ�pS��
!j��<E��T&��   �   l�%�t����
���	�,]�/d�g�"�ۥ-�U�6�D=�)?���<�F�6�t�-�$"����/�����Qҽɦ���^����u�2�?����
mü�7u���X���0J�8'��t�4��̩�6���Y�����Nֽ"����5�eb�`j���P���X���Ͼ.b�?�꾋��d�ʝݾ��˾6��P���dL��)d�_�@��   �   I�9���%�Ɓ����{���R(���3�f�>�ƔG��LL� L�h�F�*=�N�/�K����������Aֽ`(��)͓�r�j�4�2�j��:���4�/�PW� ;h6�; ��;���:hc����z�Rx����M�:���.�ڽz����@�XTs��3�������>;��� ;�������d�u���V)���˾΂��,j���`��W��   �   +I�I�3�s�(���&�z�+�޶5���A���L�"U�!�X��"W�/�O�+4C��2����jh�>��:�Ž�r����{�!=�Q��Z�����$� �Ӻ8מ;Xo<�S7<|�,<���;����83A����R�G��Q�� ཝ��0J�케�ើJ���|ܾJ�������k�ֻ��B��M�LV���
ݾ@j��}���_���i��   �   �S��p<�i�0�@�.�z4�'M>��wJ�%�U��^�h>a��^���U���G��55��: ��
�Ҏ�5���
j��k�b�%�"�^�ԼT5g�0E��0�u;��<p�[<t�s<<a<X�<�>�:4!�|u׼�}E��P��#�vw�Q�P��l��0;���Aƾ�e澨������J�d��A�(�����T辙�ɾ;���4���Hu��   �   �}V��y?���3���1��6��AA���M��X�!a�(d��a��W��I�e 6�S} �*�	���彶&��������Z��9�2lü��E�@�����;X�7<�Vr<<��<�r<�+<@�/;��4�Ӽ��D�����=~�;��O�R�b���p���ɾ���)��$2����<����sH��������D;w��ߎ���?y��   �   �S��o<���0���.��4�XL>��vJ�>�U��^�{=a��~^���U�ځG� 55�: �%
���罉����i����b�z�"�t�Լ�3g��B��0�u;h�<<�[<(�s<Ta<��<�K�:�!��s׼�|E�P��,��v�z�P�l���:���@ƾ�d� ��+��J����d@����d��]���ɾ\:��;4���Gu��   �   j)I�ƕ3��(�L�&��+�Q�5�P�A���L�@ U�]�X�!W���O��2C���2����rg������Ž�q��B�{��=�h��������$�`�Ӻpڞ;�p<4U7<@�,<��; ����.A����M�G�uP��!�`~�/J�軀��ߞ�����zܾD���܊�]j�����A��L�:T��	ݾ�h����\^���i��   �   �9�c�%������p���P(�d�3��>�U�G�JL��L�*�F��'=�x�/����,��P���@ֽ'��̓���j���2�z��������/�0�V� ;�:�;P��;�
�:�Z����z�t��̿M�J�����ڽ���j�@��Qs��1��i���<<;���8��K��n��rb�[���}&�9�˾����Fh���]�^�W��   �   ��%����U�
�C�	��Z��a��"��-�l�6�W=�D&?�/�<���6�B�-�4""�b��޴��	�FPҽ{����]��3�u��?�ޱ��kü\5u�l��R��`$J� ��8�4�0ɩ����9�X�r���0ֽ��Q�5��ab�Jh��N���U����Ͼ�^�l�꾢��`��ݾX�˾3������ J��0%d��@��   �   v������R���J��nf�Z^����+#%�\+-� $2���3�p2��U.���'�K��1��l�
�M(���i���Ž y��y슽S
]��")��[���ֳ��x��,�b��t��H��Z*���'�el�A���ԽL5��*�z�P���y�~���0���UG����ľf.;i>Ͼ�ʾ�B�������ϝ��P��j�O8E�YQ&��   �   �S�`Tӽ��ƽ�}ƽ�Qн���#���^�D��`���&��B-� \1�qG3��3�®0��,���$�6w�<���l��^�K½rҠ�v����L�r���{ ���߼�޼�e��PJ�~�K�����w[��u׽j"��!��A�b�&���z=���Ҟ������㯾�u��|��6��������Tf�V�C�ĺ$�m�
��   �   y���]�u��o���XR���G��2zӽ��`��8�6�j�*�# 5�<�=�"�D�'�H�	�I��HG���@���5�+�'�a*����A�ݽ�ͷ�����Fs�AJ�8�1�@0+���5��P�j�z�\�3���gམk��m���4���M�5Vf��}�����.|�����!u������:s�6X�n;�����U�ݽ�   �   ����4}��tp�Y�v�dA��>e��8a����нn0񽝽	��c�)-���>��N��`]�h�h�&p�;"r��cn�Ȩd�vdU�O�A�W�*��������v̽\@������@9}�?yp�j�v�QC�� g��c����н�1��	�4d��(-��>���N�_]�V�h��p�er��`n���d�faU�j�A���*�&������{r̽P=���   �   �J��1�u,+��5���P�G�z��옽�2���f�^k��m�z�4���M��Wf��}�J������}��f���v��r���=s�-X�;�������ݽT���什Lw������xT���I��H|ӽ���D���8�����*��5���=��D���H��I�yFG�B�@�#�5���'��'����+�ݽʷ������s��   �   �w ���߼ ޼�_���G���K�x����Z���׽i"�f�!�UA�Nb�����>��_Ԟ����m
���䯾�w��\����������Wf��D�ʼ$�!�
��V��Vӽ.�ƽ'�ƽTн���d���y�P��	a���&�FC-�$\1�2G3�:3���0�",���$�Mu�5���j��Z㽓½Ϡ�v���GL����   �   Dr����b�<t��C��&��'��l�����TԽv5�~�*�c�P���y�q���j����H����ľ@0;[@Ͼ�ʾ�D��Ľ��=ѝ��Q��|j�L:E�S&�������GT���L���g�~_����L$%�i,-�%2�x�3��p2��U.���'����B��<�
��%���f���Ž�u���銽�]��)�S��fϳ��   �   p>���J� ����4��ũ�P��&�X�*���9ֽU��߅5��bb��h��O��%W��&�Ͼ(`�+��w��b��ݾ�˾�4������9K��'d���@�ت%����Q�
�6�	��[��b���"��-���6�g=�<'?���<�h�6���-�?""� ��X���iNҽa����[��ƿu�͓?�ڭ�Rdü\(u� ��   �   �H�;x��; 8�:�P��(�z�Lr���M�%�����ڽ���@�TRs��2��3���9=;��l9����3��:c������'�z�˾����3i��_���W���9�B�%�������0��YQ(�@�3���>�I�G�	KL��L���F��(=���/����0�����B?ֽ�%���ʓ���j�
�2�����*�����/�p�V�P3;�   �   `Y7<�,<���; 7��,A������G�bP��9ཌྷ~�u/J�.���'���L��{{ܾ���W���j�3��1B�kM�?U���	ݾpi������^����i�*I�W�3���(�ŝ&�~�+�ص5���A���L�� U��X��!W�<�O�D3C�3�2����g�����ŽBq����{�w=������X�$���Ӻ��;�u<�   �   ��s<�a<��< V�:�!�4s׼@|E��O�� ��v���P�,l���:��#Aƾ(e�R��f��GJ�
���@���������-�ɾ�:���4��%Hu� S��o<���0���.��4��L>�(wJ���U�L^��=a�a^�0�U�L�G�g55�q: �k
�]�������i����b�7�"���Լ�1g��>����u;\�<��[<�   �   �Ӑ<��<X@Q<���;�WV�x ������\��X��ཞ��ރ;��f�mg���͞��߱������ʾ��;n�ʾUD��(��2�0ޏ�I�}�ʁa�w�M���C�j-D���N�|�a���z��?���ј�D6��iի�}����ҫ��գ�,Y��ʅ���ek�1^F��("�,^ ���ýh����B�ȥ� �d����x#�; MS<�<�   �   "��<T4|<�?<pB�;hM��X�����
���_�R��b�߽���$:�\d�$އ�nќ�cw��*3��S�Ǿ��ʾ�Ǿ�<���G���c�����`�y���]�7UJ���@��A�8hK�^�<�v�>���p�������8������e`������Vx�����)4i�_�D��y!� N �0�ĽV����F�����|Hz��"b�H�;L??<�4{<�   �   �jW<��D<��< ��:�c�������p���h�|���9�߽�>�HY6�%.^��{��<��*����@���ﾾP����g��/w��������<���3n�5�S��@�4y7���7���A��S��9k�����P����X���������W���L��^������c�XA�Ϸ�%_ �a�ǽ����a�T��t��蝼�m�� ��:�a<�1A<�   �   `f�;�B�;P�!;����H�]�>�ռF6+��y�@��u:὿@�1�@&U���y�����������ᕱ����� W��1ڧ�]��^b��Ly�J�[�5C�W�1�>>)��)���2��vC�iMY�p�q��΄��������,����������b󇾮�v�� Z��;�ǽ�@I�]ν����bm���&���ּt�j��p����:`�;�   �   �������ĻD�N�����p!K��m��Y:��w��=5��+��K��sj�� �����F�����K��D�������I��}k{��_�eqD��U.�2������n�G����.�]|B�b�X�R�n�J���G���<犾qP���腾�_|���g���O��~6�����*��ڽ̯����(�O�.O�d�Ǽԗq��K����K��   �   |�N�@\�|����kżp,
�
b<��lx�z����Ž܀�0��ZM(��A��![�װr��g��%ڊ��莾����3��\�����r�7_Z�:NA�*�)�{��&�����t���	�@�z�(��q<�,DP��a��+o���v���w���r�&h��Y� G��+3�Ǳ��]
�/d���ǽꤽ؈��~�N�ԃ����~���$Cr��   �   ��ڼ����� �AE��?G�s&z�L���v��f޽\��ʤ��)(���;�7*N�n�^�4�l�'�u���y��dw���n��Q`�V~M��8��F"���V���l"�Cx׽�[ؽu>�zk�����7��&1�ҖA�N�N���W�}�[�B�Z�Q�U�,�L�"A��3���$��-�-�����ɽ�%���B��6Xb��14�/B�\���   �   �&2��4��mF�^Bf�=��t����0���t�e ����ړ�^�,���9��mE�O��U��HY�9�X��$S�l&I��;�q�)�����������Ƚ_���r̪�����7����-˽�D���� >���"�2�0��U;�3�B��yF��	G�<�D��?�9�m30���%��L�|z�����gٽ����]��Tl��f�[��_?��   �   v%��f6������ל��[lѽ�$�-{�����"���-���6���=�f$B��D��rD���A��<��d3���'�)S��	����νH��u�>6���"��p3�����^Ԝ�2봽�hѽZ!�y�����"���-���6�h�=��$B�Z�D��sD�9�A�l<��f3�ѭ'�UU��	��#��ν�������H9���   �   �Ϫ�*ë����E1˽�H����@���"��0��W;���B��zF�!
G�P�D���?�:9�@20��%�K��x�Q���dٽ�����Z��Li����[�Z?��!2���4�;hF��<f�c������.��r�,
 ����*���,��9�xnE�O���U��JY�f�X��&S��(I��;���)����������c�Ƚ�����   �   �{׽�^ؽ�A�#o��ء��9��(1��A�Z�N���W��[���Z�%�U���L�A�i�3��$�\,��+�����ɽ�"���?���Rb�t,4�C=����ڼ���%� ��@��:G��!z����Y���޽��o���)(��;�"+N���^���l�K�u���y��gw�M�n�WT`�ʀM��8��H"�x�ڪ���%��   �   4�Hv���	��q�(��s<�XFP�F�a��-o���v�\�w�2�r�'h�_Y�: G��+3�6��#]
�b��ǽ�礽Z�����N�D�F��B����3r�\�N�1\�򖍼Zdż�(
�c^<�_ix������Ž�����M(�0�A��"[�e�r��h��Hۊ��鎾D��I5�������r�yaZ�LPA�
�)�5������   �   ��Cp���W�.�@~B�d�X�i�n�V���K���-芾DQ��y酾�`|���g���O��~6����@*�+ڽAʯ����2�O�HK��Ǽȉq�01�� �K�����p��kĻ��N����K	��K��l���9��/��_5���+�vK��tj�P!��~ ��b����^L������J���
K���m{��	_�sD�`W.�����   �   �?)�h�)�1�2�vxC�OY�1�q��τ�q���������V���=�����/�v�7Z���;�{���H��[νK���!_m���&���ּD�j�[��@k�:��;�x�;8T�;0";�w�� �]��}ռ�4+�ǌy��?��~:��@��1�'U��y�����` �����얱�����X��:ۧ�^��Cc���My���[�l6C���1��   �   3z7���7��A�Y�S��:k�r������dY��)���O����W��HM�����4���c�6A�����^ �b�ǽq����T�>r�䝼�]���=�:�h<�8A<�pW<�E<d�<���:8Y��0����o� �h�c���k�߽?��Y6��.^�,|�����ӌ���A��V� ���^h���w�����P�������Hn�;�S��@��   �   J�@�A��hK��^��v����q���79�������`������fx������3i��D�8y!��M �[�Ľ:U��=�F�L����Bz��b� �;�C?<�8{<��<�7|<�"?<pH�;�G��:���c�
�ň_�_����߽@���$:��\d�nއ��ќ��w���3��ƟǾ0�ʾ�ǾV=��<H��5d��Z�����y�U�]��UJ��   �   ܥC��-D�X�N�ݤa���z�@���ј�^6��uի�z����ҫ��գ��X�������ek��]F�E("��] �9�ýê���B�֣���d�p���(�;�NS<��<LԐ<��<@AQ<���;VV�p ����ӯ\��X��?� �	�;��f��g��Ξ��߱�*�����ʾ��;z�ʾ^D��2��;�;ޏ�d�}��a���M��   �   }�@��A�"hK��^��v�!��~p��B����8��D����_������w��e��3i�R�D��x!�=M ���Ľ�T��Z�F������@z�`b���;�D?<�9{<t��<�8|<�#?<�J�;�D�������
�_������߽���/$:��[d��݇�'ќ�w���2����ǾX�ʾHǾ�<���G���c��Ö���y�f�]��TJ��   �   �x7��7�v�A���S�9k�Z���Չ��X��ԯ������OV��
L��}��0���Gc��A�X���] ���ǽP���b�T��p�2❼�W��@P�:�j<:A<drW<�E<��<`��:�R������n��h������߽�=�ZX6�-^�${�����y���"@��������f��pv��Q��
�������Hn�r�S�j�@��   �   \=)�;�)���2��uC�TLY�*�q��̈́�������� ����������:�b�v���Y���;�׻�tG��Yν�����\m�"�&��ּ,�j��T�����:��;}�;Y�;�";@q����]�lzռ�2+� �y��=��8�v?��1��$U�<�y��~���������Ŕ�������U��$٧�\���a���Jy���[��3C�^�1��   �   ~���m�$��\�.��zB�¥X�t�n�:�������劾O��l煾]|�:�g��O�A|6�����(��ڽXȯ������O��I���Ǽ$�q� +���~K��}�����HdĻ��N�6��p�tK�k��s7��N�彊3�:�+��K�wqj�W��F�����p���I��︞�ϻ���H��gi{�_��oD�eT.�����   �   L�`s���	���ן(��o<�BP���a�')o���v���w���r��"h��Y��F�)3���l[
�k_��ǽ�夽-����N��}�.�⼜����0r�h�N��-\�(���,bż1'
�^\<��fx�"���y�Ž�|� ��#K(��A�[�#�r�:f���؊�&玾s��|2�������r��\Z�4LA�`�)�������   �   ~u׽�Xؽ�;�`h��(���5��$1�P�A���N���W�c�[��Z�
�U���L��A�3���$��*�f*����k�ɽ�!�� ?��FQb�_+4�c<�\���ڼ���<� �t?�q9G��z�����~��(޽~�j��'(���;�n'N���^�.�l��u�h�y��aw���n��N`��{M�E8��D"������{��   �   �ɪ�:���S����*˽~A�����;�?�"�w�0��R;��B��vF�;G�صD���?��9�-00�b�%��I��w������bٽ���Y���h��߁[�VY?�� 2�ݚ4�MgF��;f���������,��Sp�� �0��;����,�)�9��jE�O���U��EY�"�X��!S�#I���:��)�S�����n���}Ƚn����   �   ����0�����Zќ��紽'eѽ� w������"���-���6��=�>!B��|D�jpD�˻A�<�uc3���'�yR�	���k�ν�����5��-"��3��+���Ӝ��괽
hѽ% �x���T�"���-���6���=�u!B��|D��oD���A��<��a3��'��P�5	�|�8�ν���fr3���   �   �2�Ŗ4�cF�G7f�P�����'*���mཻ ���N���,���9�kE��O��U�VGY��X��#S��%I��;� �)�C�������佤�Ƚ���&̪���������V-˽eD潐���=�	�"�F�0��T;���B�xF�@G�s�D���?�r9��/0�b�%��H�:v������_ٽ��@W��8f��)}[�U?��   �   ��ڼ��༙� ��;�}5G��z�����h��>޽H}�ӡ��&(�	�;��'N�w�^���l���u�y�y�$dw�	�n�HQ`��}M�X8��F"�d����("��w׽P[ؽ >�k�����^7�S&1�>�A���N���W�;�[���Z�^�U���L�xA��3�y�$�	*��)����!�ɽV���<���Lb�#'4�m8� ���   �   ��N��"\�4���\ż$
�Y<�ecx������Ž�{�Ή�K(�p�A��[�H�r� g���ي�:莾����3��.���_�r��^Z�NA��)�\����|��t���	��H�(�Iq<��CP���a�0+o���v���w���r�{$h��Y���F��)3�*��2[
�v^�.�ǽa䤽r���a�N�jz����@����$r��   �   @7��P��hRĻ �N�T����	K��i���6�����k3�a�+�K�Grj����	�����~���J�����𼖾�I��Wk{��_�IqD��U.�������n�-��~�.�<|B�8�X��n� �������抾P��T腾�^|���g��O��|6�����(�Yڽ�ǯ�������O�7G���ǼL|q�(���ZK��   �   ���;He�;�5";�c����]��vռ�0+�y�y�>=���7�q?��1�#%U���y�c��+����������t����V��ڧ��\��Pb���Ky�5�[� 5C�F�1�.>)���)���2��vC�NMY�Q�q��΄�l���������_���T����򇾮�v���Y���;�W���G��Yνz����[m���&���ּ��j�H��`��:@�;�   �   �uW<E<�<��:@J��Ԫ���l�*�h�����u�߽�=�~X6�o-^�g{�����򋨾�@��lﾾ7���~g��"w���������2���&n�(�S��@�(y7���7���A��S��9k�����C����X��i��������V���L��������6c��A���(^ �P�ǽs���B�T��p�����0Q���j�:4n<x=A<�   �   �<�9|<%?<`N�;�@������
�+�_�n����߽���0$:��[d��݇�Mќ�Hw��3��B�Ǿ��ʾ�Ǿ�<���G���c�����U�y���]�1UJ���@��A�0hK� ^�3�v�8���p��z����8������Q`������6x������3i���D�y!��M �+�ĽU����F������@z� b�h�;�E?<X:{<�   �   �.�<�)�< �H<��;`Qݺ�gG�ܘͼy&�I#p����0ҽ�.�p����:��eU���l�_O�v����x��5���)����p���^��N��<A�O3;�H4>���K�<d������d��{��˾Zu�Zp��K� ����� ��:����[�Ⱦ����7e����i���6��
�܂ǽ�Շ��(���p,ϻ�#�;�@<@��<�   �    ��<�9m<x1<�r�;_\�8�c�b�ۼ��,�}Av�������ӽ�{��z���9�#�S���j��Y|�Lʃ�"���P���,}|�m���[���J��1>��<8�w/;�fxH� �`� ���7�!��6�Ǿ��޾f�����U��������<޾~�žK�������� g��G5��3	���ƽz"���o*��`��x��P�m;�>0<�p<�   �   0�I<@-<��; �	9�h
�؄�����/B�V����ˬ�\>ٽ{����O7�b�N��c���s�h�}��@���|��oq��kb��~Q��A��U5�Ú/�Mc2�S?��V�H�v��ڏ��ڦ��s��rWԾ.澒��'��Q�&��ʰԾ�Ͻ��'��g����`���0����u�Ž0Q��[s0��iż�u�@5d:���;p<<�   �   pA�; (�;@�`�����^�� ^���)��g�����'���� v���,�3��LH�T�Y�;?g���n��-p��	k��c`�V�Q�	�A���2�*o'�6"�I�$��>0� �E�	�c��Ä�I����Ư�bľW�Ծ��߾(�� yྂ<־�ƾ�g��H4��.����U�S*�ز��ĽRB��� <��1伀e�x����);���;�   �    �'�`���|�;��!��t���*��b�|7�����3�ѽ�j����"v�k31�VA���N��KX���\�a0\���U�� K��,=��.�|* �R�����:���D�\X0��K��Pm�
����2��\^��R���jȾt�̾7+ʾ����$۳��'��.���lr��I�lP#�`� ��ŽS���+O���	�tq���.5�(��p��   �   �h����h�мo���>�l�t��j��ơ���DԽ���b�h��I�$��?1�T<�HD�/9I��-J���F��?���3��&�����
�Z[��h������ă�G%�Q�/� UM��n�EK��/;���|������&ϲ�����q��3������K��� `�b�=�Jc�������ʽ���8l���+�������h�x���U��   �   �I���5e0�(A_��M��N���<8ɽ�D轜��6@�s'�;g&���.�o�5��>:�؉<�r<���8�#�1�A(���
y�D� ������׽�4ϽͬѽE����޵���+�ZH�Ee�a��f����Z��?���D���rZ��#q��U���nZj��rO�sQ4���֋�'ֽ�ޭ�����}�Y���)��R���弄�ټ�   �   fh<�hZ�fO��b����������!���	�|w"��7.�*�6�-�<��t?��?��{=��$9���2��9*�}���|�D��f�Yqսe���X�������f��$�����ɽݑ�*�
�2�"��$;��R��g�ewv�l��6��1�~��u�zg�D�U���B���.�����/�t�轜�Ž�ǥ��ʉ���e�$�D��1��.��   �   ����YW��}ߴ��׽�����B�;x(�.�:��6I�9�S�c0Y�p&Z�R�V��%P���F�`;�.� �~A�3��"T���ǽ��;k�� ����]z��Jz�v����S���۴���׽����+@��u(�i�:�/4I���S�.Y��$Z���V��$P�+�F�b;��.�� ��B�n���V���ǽ��n�������cz��Pz��   �   ����j�ɽ�뽊�
�Ԃ"��';��R��g��zv�e��l7��|�~�yu��g��U�ԷB���.�2��/�v��\�Ž�ť�ȉ���e�4�D��1���.��b<�=Z�L����������1��ԋ�F�6u"��5.�V�6���<��s?�S�?��{=��$9�n�2��:*�ǿ�~����|�jtսn���W�������i���   �   ���
�����+�&H�*He��b����V\��߫�������[��0r�����y[j�TsO��Q4���F��{%ֽ�ܭ�����[�Y���)�>N�҄�p�ټ&@����n_0��:_�^J������4ɽ�@�����>�&�2f&��.�4�5�?:�v�<�h <��8�� 2��B(�+��z��� ������׽�7Ͻ�ѽ�   �   ���A'���/��WM���n��L���<���~��l����в� ������J�������K���`���=�0c������ʽH���4l��+����権���x�`�U���h�8����м�i�]�>���t��g��឵�DBԽ`��a������$��?1��<��HD�S:I��.J�B�F�??�M�3�y&����Z�
��\��k�������   �   UF�<Z0�2�K�Sm�f���;4���_���S���lȾ�̾�,ʾܦ��*ܳ�N(������mr�2�I�cP#�� ���Ž�Q��X)O�'�	��k��@#5�p����0�'��޺��v;����
��;�*�=b�b5�������ѽ�i��K�v��31��VA���N��LX���\��1\�Y�U�Y"K�.=�(.��+ �¦�������   �   J@0���E���c��Ą�~���&ȯ��ľȌԾ#�߾~��2zྍ=־xƾ�h���4��P.���U�S*����P�ĽZA����;�|-伨e�� ���);8�;�T�;�<�;@`�����X���W輬�)��g�>���$��s��v�?����3�uMH�5�Y�N@g���n�*/p�k�be`���Q�U�A���2�ip'�|	"���$��   �   �?�(V���v��ۏ��ۦ��t���XԾ2/澣��(���Q����S�Ծ-н�3(������`���0������ŽYP���q0�dfżo���d:���;<<<�I<TG-< ��; ~9�`
�܀�����wB�����3ˬ�>ٽ�������7���N�9�c���s�\�}�A���|��pq��lb��Q��A��V5���/�bd2��   �   ;yH��`������������ǾF�޾��N�����b���)���<޾��ž@�������7 g�_G5�3	���ƽ�!��qn*�$^��H���m;\C0<T�p<<��<D>m<�1< {�; N\�$�c���ۼ��,��@v�������ӽ�{�{��9���S���j��Z|��ʃ�q��������}|��m��[�5�J�;2>��=8�50;��   �   	�K��<d�����d����+˾�u⾆p��V� ����� ��:��ь�
�ȾH����d���i��6�]
���ǽՇ�̓(��뮼�%ϻ�)�;<@<L��<�/�<�*�<8�H<��;`Kݺ8gG���ͼ�&�y#p�2���?0ҽ�.�����:�
fU�"�l��O������x��D���)����p���^�N�=A��3;��4>��   �   dxH�%�`� ���2����ǾX�޾��?����V���+��<޾��ž����
���Mg��F5��2	��ƽ!���m*��\��8�� �m;�D0<L�p<���<?m<�1<`}�; I\�x�c�x�ۼ7�,��?v������ӽl{��z�<�9���S��j��Y|�ʃ�䚅�����||��m�2�[�[�J�n1>��<8�j/;��   �   �
?�\V���v�cڏ�1ڦ�s���VԾF-澠��&���O���澙�Ծ�ν��&��i���
`�S�0�x���Ž"O���o0��cż,k���d:`��;<<��I<�H-<���; �98^
�<�����B�����ʬ��<ٽ������U7�_�N�q�c���s�O�}��?���|��nq��jb��}Q�B�A�LU5�B�/��b2��   �   >0�0�E��c�Ä������ů�Y ľ#�Ծ_�߾���uw��:־ƾdf���2���,��~�U�Q*���
�Ľ�?��Y�;��)�Te����� *;p	�;hY�;A�; �_�t���V���U�9�)��g��������`�㽴t������3�FKH���Y��=g��n�F,p�/k��b`��Q���A���2�?n'�g"���$��   �   �C�8W0���K�%Om�����1��]���P��ZiȾ��̾e)ʾģ��Uٳ��%�����jr�L�I�N#�R� �A�Ž�O��Q&O���	��h��|5� ������P�'�Hٺ��s;�x������*�~b�<4��������ѽNg����4t�t11�TA���N��IX���\�p.\���U�K��*=�4.�1) �(�����4���   �   ����#���/�2SM��}n�J���9��;{��⩮�;Ͳ�����p��>��ݶ��ZI����_�{�=��`������ʽ
���1l���+�,��2�����x�$�U��h���`�мi�6�>�M�t��f�������@Խ@��:`����$�t=1��<��ED��6I�6+J���F���>���3�&�u��R�
�Z�>f��4����   �   ���/��6����+�H�wBe��_�������X��G���=���fX��!o��g����Vj�joO�^N4��L��s"ֽ�ڭ����܈Y���)��L���弦�ټ�>����^0�:_��I�������3ɽ�?�����=��$�}d&���.���5�)<:�B�<��<�=�8���1��>(�|�.w��� ������׽2Ͻ8�ѽ�   �   j�����ɽ���>�
��}"�1";��R�sg��sv����4��2�~��u��g���U��B�Ծ.�¹�+-����*�Ž�å��Ɖ��e�ܣD���1���.�b<�{Z��K��:������}��a����mt"��4.�
�6��<��q?���?�(y=��!9��2�7*�%��ez�>����nսX�������?��d���   �   ���Q��lش��|׽�����=��r(�Q�:��0I��S�b*Y�� Z��V�� P���F��;�O.�� ��?����R�{�ǽ�쬽jj�������\z�Jz�����S��J۴�9�׽P����?�u(��:�{3I���S��,Y�#Z��V�u"P���F��;�|.�� �:?���GP�z�ǽ�ꬽTh��p����Xz��Ez��   �   �]<�
Z�I��L���ʚ�����V��~�0r"�M2.���6�D�<�"p?��?��x=��!9�O�2��7*����n{�e���bpս����ʹ��~��Xf��Ԛ��T�ɽ�����
��"��$;���R�Ng��vv�����5���~�u��g�"�U� �B�_�.����,������ŽY¥�.ŉ���e�I�D�S�1�$�.��   �   �7�*��CZ0� 5_�G��د��'0ɽ<�1���;�!#�#c&���.��5��;:�d�<�q<��8���1�@(����x��� ���M�׽R4Ͻ}�ѽ���������q�+�/H��De��`��8���fZ��縉�ݜ���Y���p�������Xj��pO�AO4���f��"ֽ�٭�����X�Y��)��I��|�<�ټ�   �   ��h��얼.�мe���>�C�t�Ld��֚���=Խ���_�$��C�$�!=1� <�&FD��7I�4,J���F�� ?��3�b&������
�,[�jh��\������+%�1�/��TM��n�2K��;���|�������β�K���
�����#���eJ��b�_���=�ha�������ʽ�	��Q0l���+�@��¡�� �x��U��   �   �^'�ƺ��h;�,�����*�ib�)2��������ѽ�e�� ��s�\11�BTA�;�N�NJX���\��/\�3�U�S K�9,=�i.�M* �1�����!���D�EX0���K��Pm������2��J^���Q���jȾL�̾+ʾT����ڳ�'������kr���I��N#��� �ɢŽ�O���%O��	�f��`5�`񣻰���   �   �d�;�N�; ~_�`��R��$P�R�)��g�����2��L��Qt�u����3��KH�?�Y�[>g��n�N-p�L	k��c`��Q���A�p�2�o'�""�8�$��>0��E���c��Ä�A����Ư�WľI�Ծ��߾���x�R<־`ƾ�g���3���-��ȟU�R*�±�؎Ľ@����;�8)伸e��񀻠*;p�;�   �   ��I<�L-<���; ]9�W
��{�����&B�����*ɬ��;ٽP��n��]7���N���c�%�s���}�^@���|�doq��kb��~Q�ۀA��U5���/�Ac2�G?��V�>�v��ڏ��ڦ��s��lWԾ.澈��'��Q��澢�Ծ�Ͻ��'��"���3`�:�0�$���Ž�O��}p0�@dż�j�@�d:���;|<<�   �   ���<@m<T1<���;�=\�8�c���ۼ:�,��>v�����r�ӽ?{�fz�/�9���S�0�j��Y|�2ʃ����B���}|�m�|�[���J��1>��<8�q/;�axH��`����6� ��4�Ǿ��޾b�����Q�����ԁ�<޾i�ž/�������: g�jG5�,3	��ƽ�!���n*�"^������m;D0<p�p<�   �   L�e<�N<��<��P;��l&[��üQ��"G�h���U��^��[���o�G���'��-���/���-��4)�a8#�E�l��E�!�S�/���H��n���.�r�վE��������$�#L3�(�<�!�?�J�<��;3�؋$�E�����о�U��9��+�C�,����½
�x���`�s� ƒ�h��;4EN<�   �   <�O<H�4<���; ?�:��ڻ򧂼��ټ�X�8>R�$���F�طý�佁����q+���&��n,�?	.���+�*�&�F� ����Ԇ�)m�� -���E��	k��������&�Ҿ�����h��)"��e0�9�9��<��9�'e0���!�,�������;�
������*�A�l�����5�w�I���y��>�X:�;��<<�   �   py<��;�$�:x����c���¼���'@� Yt�J����@��z�ϽS�콚���\�A���#��C(���(��%��X ������<{���Q%�}�<���_����9᥾��Ⱦ���w�	�5j���'�i�0�t�3���0�[-(�G��)L	����zľGs��s�w��;����ż��u�2��8�� �p�hY�;�G<�   �    �:���~Q��B�ռ�O�g!I�v�{�Nޗ��ձ��˽\��}%����	�����J��^ ��N"�w� ����@a�����C
�vs��j��N���-�-�N���z���븾�E۾����2Y�=��e#��%�1Y#��k����{���ab۾j4��o_���i��\1�^5����$�r�.��.ؚ��}� �b���+;�   �   �?��]�p�������p3�dh�g,�����S�ýP	ܽ����g��l��Pq���NE�l��R��|��t8
�B��^���B��������yM� �8�40`�l����'����þ�X��,���M
����Di�q<��_��� ���徼�ƾƦ�p��$�W�g�%�����E��W�r�;Z�6����lM�`z�ȉ���   �   0﫼���|�"�K8X�������N�Ƚ9�T< �RT�,���T�,P!�/�!�i���>�I���S�Ӓ�����齈�۽�0ս�;ٽ�꽱���[�:�A��ml��ڎ�n\����þ"�۾�n�ni���� �A�����:�ླ�ɾկ�┾lu��E�y)����W��)�w�I�+��4�ࡣ�V���ʇ��   �   ���� E�u(�ޡ�PmǽQ��m�	�Y$���'�^2�j�8��';�HZ:��6��j0�MY(����l�<~������0�̽J����e��%����1ý|�޽�����!���E�v@o��)1��ˋ���#ɾLaԾ/پ�!׾��ξ�O����+���2��>�[�ͼ3����O�������D����B�^����(O�f����   �   Ӗh�����;����⽗	�|� ��q7���J�)�Y��[c��*g��`e�#�^�$�S�u.F��6�G&��B�a���y�*L̽�H��T$��찔�l�$ ��w���f[Խ���ږ��A��if����r]��	?���쭾E����ʱ�ޫ�9���bē��烾)Af�E�D�KM%��f���ݽ����i���Nc���=���*��S+�n@��   �   	�� Ƚ0���mR���4���R��(n�(����	��J����:��猾�/��Q�y�&jc��QK�D�2�%��`����-����Ν����J�o�`md�1	n�冽_����ǽ���}O���4��R��$n�������9����8��a匾J.���y�rhc��PK���2� ������ད���rН������o�Ird��n�C膽�   �   n_Խ������d�A�mf�����_��kA�������)ͱ�૾䁡��œ��胾�Bf�"�D��M%��f��ݽ뎱�h��<Kc���=���*��N+��@�I�h�F���#7��p�⽺	�P� �!n7�Z�J���Y�Xc��'g��]e�ɞ^�R�S�(-F�G�6��&��B�ϥ��z��M̽�J���&��Z���Œ�#��񫱽�   �   ��}�!���E��Co���g3��<���S&ɾ�cԾ�1پ$׾ׇξ�Q��aﭾO���3��D�[�V�3���������rC����B�%�T�F㼮���Y��(E�� ��١��hǽ���	�x!���'��2��8��%;�X:���6�	j0��X(�������~�,�� ��b�̽����|h������%5ý�޽�   �   ^�ƿA��pl�g܎�z^��G�þ��۾�q�l���� �wC��� ���2�ɾD֯��┾!mu�hE��)����%W��P�w���+�d/鼤���2������嫼2��^�"�^1X�@��f�����Ƚ�4�: �6R�-*�~���GO!���!�I���>�Ǳ�cT�����������۽t3ս�>ٽ=�꽄���   �   -�8��2`�ൈ��)����þ�Z�L/��O
�ݬ�wj��=��`�X� ���ǡƾ�Ʀ������W���%�n��UE��ʫr�DX�����LbM�@c��o���0���\�ކ������j3�h�)��;���ý6ܽV���������q����E������d��v9
�X����������������:O��   �   �N�2�z�Y	���츾�G۾����=Z�O��u#��%�Z#��l�> �����0c۾�4���_��;i��\1�?5�)����r�����Ԛ��m� y`���+;�f�:���<���I����ռ*K��I���{�ܗ��ӱ��˽���z$����	�����J�@_ �wO"�2� ����'b�����D
��t��k��O��-��   �   c`�����O⥾قȾ ��<�	�k�Z�'�3�0�0�3�:�0��-(����|L	�3�:{ľgs��{�w��;���ż�Au����5����p��f�;LO<p�<���; t�: ���4c���¼x��&@�!Vt����x?����Ͻ��콄���\�~���#�D(�3�(���%��Y ���\��|���f	%�Ǌ<��   �   �
k�<�������Ҿ����-i�>*"�f0���9�g�<�6�9�`e0���!�=������i;�
��p���ÊA��������w��G���y����C�;��<<P�O<��4<���;�m�:@�ڻФ��b�ټ<W��<R������񣽙�ý�佌��
���+� �&�+o,��	.�)�+���&��� ���j���m��!-���E��   �   ��n��������վ���������$�BL3�6�<� �?�7�<��;3���$������о:U���8��u�C������½d�x����|s� ������;�GN<��e< �N<��<��P;`���%[���üU��"G�8h��V����.\���Do�r��E�'�3�-��/���-��4)��8#�JE������!���/���H��   �   �	k��������'�Ҿx����h��)"�Fe0��9���<�p�9��d0�2�!���������;
��ꎀ���A�n����m�w��F���y� 	�8G�;��<<8�O<T�4<h��;@t�:8�ڻ8�����ټ�V�?<R�3���V��ý����~��+�W�&�xn,��.�o�+���&�� �������!m�� -��E��   �   ��_������ॾ,�Ⱦ���	��i���'���0���3���0��,(�r��\K	�F쾤yľ"r��~�w��;���nü��u����2��@�p�Pl�;HQ<�<���;@�:@����	c�j�¼���)@��Tt�8���|>��r�ϽW�콢���[�X���#��B(�ֽ(�V�%�WX �\����z�g��%�/�<��   �   h�N�	�z�n��D긾�D۾[���vX�a��m
#���%�X#��j�}��t����`۾�2��^��}i��Z1��3�����\�r�~��К�Pc� �_���+;�x�: ��X���H��Z�ռ[J��I�b�{�*ۗ��ұ���˽1��e"��x�	����I��] ��M"�L� ����B`�ʞ��B
��r�j��M���-��   �   �8��.`������&��C�þ�V�+���L
�t��h�(;�?^�B� �l�徢�ƾ;Ħ�����d�W��%�����B����r�JU�n���\M��Y��h��<.�|�\��������j3�!h�u(��w���ý�ܽ����M��f��_o���C���������.7
���R���Z�����&���L��   �   �Z���A��kl�lَ��Z��8�þ�۾�l��f��*� �O>�������:�ɾ�ү�����hu��E��&����T����w���+��*�8�����������`䫼և켺�"��0X����臩�E�Ƚ�3潏9 ��Q�I)�a�����M!�Ԍ!�3���<�`���Q�5������#�۽�.ս�9ٽ�꽊���   �   ���C�!�{�E��=o�2T/������`!ɾ�^Ծ^,پ�׾�ξGM��h뭾����0����[���3�&���{���A��w�B��|���D㼰������sE�Q ��١�&hǽ���Q�	�!�n�'��2� �8��$;� W:��6�*h0��V(�w��L�P|�����_�̽�����c��Ұ���/ý��޽�   �   tXԽ���Ĕ���A��ff�@���f[���<��ꭾ����Lȱ�w۫��}������`僾1=f���D�3J%��c�Ӊݽً���e���Gc�[�=��*��M+��@���h�칑��6���⽊	�� ��m7���J��Y�jWc��&g��\e��^���S�a+F�D�6��&��@�`���u��H̽�E���!��|����������奱��   �   ���z�ǽ&���M���4���R�� n�����_��ף��p6���⌾�+����y�Vdc��LK�J�2��������V����̝������o��kd�n��䆽 ��s�ǽі��VO�^�4���R�k$n�䟂�l��񥏾8���䌾�-����y��fc��NK���2����^�������˝�������o��hd��n��↽�   �   �h�@����3��+��9	�f� ��j7���J���Y��Sc�v#g��Ye���^�U�S�l)F�Ҝ6��&�@�:��.v齱I̽�F��#��򯔽�����������[Խs�������A��if�񆅾X]���>��V쭾����ʱ��ݫ�����Ó��惾�?f���D�kK%��d���ݽ�����e���Fc�_�=�^�*��J+�*@��   �   ����E���+֡�>dǽ���}	�V���'�2�@8�";��T:�;�6��f0��U(�����i|������Ὠ�̽.���e�������1ý%�޽۵�ٶ!�q�E�[@o��1�������#ɾ*aԾ�.پ~!׾h�ξ�O��k����@2��͢[�>�3�*���|�k�&A����B�E{����?㼖����   �   Fޫ�h��.�"�M+X����J���F�Ƚs/�Z7 �LO�+'�t���QL!�؋!����W<�i��.R����Z���L齦�۽<0սV;ٽ��꽎���[�!�A��ml��ڎ�b\����þ�۾�n�Xi��u� ��@��{�����T�ɾ�ԯ��ᔾ�ju��E�&(�%���T����w���+�)�h�������޻���   �    %�0�\��~�����4e3���g�k%��<����ý�ܽ��6����z���n����C����3������7
�̪���������������_M�
�8� 0`�b����'����þ�X��,���M
����:i�c<�t_�f� �z��j�ƾ�Ŧ���2�W�d�%�l���C���r��U�戺��XM��O�`Z���   �   ���: _�t���B��h�ռjF�PI���{��ؗ�6б�~�˽6��� ����	�$���H��] ��M"��� �"���`�\���C
�Hs��j��N�v�-��N���z���븾�E۾����1Y�;��a#���%�)Y#��k�~��M���(b۾'4��"_��<i��[1��4����r��~�vњ�a� �^���+;�   �   L�<���;୼:x���� c�j�¼���6�?��Qt�����=��+�ϽC��<��X[�=���#��B(��(���%��X ���f��{���?%�p�<���_����5᥾��Ⱦ���v�	�4j���'�g�0�q�3���0�T-(�>��L	����zľs���w�1;�d��ļ��u��,4��лp�8m�;PS<�   �   ��O<��4<���;���:Ȋڻꡂ��ټJU��:R�d�����9�ý*����P���*�M�&��n,��.���+��&�+� ����Ć�m�� -���E��	k��������$�Ҿ�����h��)"��e0�8�9��<��9�$e0���!�&������l;�
�������A�0�@���5�w� H�\�y���8D�;H�<<�   �   �u<pT�;P?;��S���0�.����7꼵!�osC��kj��a�����ଽF����˽�!׽>߽����佐��+V�©潍��:*�"���)<��rl��������֫�>���Y2�[RO�BMi��}�|����⇿ϗ����}�;i�^�N��21�����K뾄l���ˈ��E�.H	�v��,BY��0⼬�#�`�:(X�;�   �   �F�;@��;@.:@�Żp^e��仼����,�b'T���z�3�����㲽D½;/ϽqٽkU�#��=�㽇�z���㽔��&&�}6�W49��h�"Z��(�����c�\s/���K�j�e���y�r��۵���v���y�I]e�vxK�zm.�����\³��ᆾTC����a+��N�W����+� ��9PV�;�   �    Y";��P�kۻ(�m�BP¼kA
�A�4�$�^��������৽����uŽ�1ѽ�uڽ��/���7=��(ݽ�ڽy3۽��佶���x8�ܗ0�U�]�^��Y���k�a��	'�0B�}�Z�2�m�glz���~���z�Tn�
�Z�*B�bh&�(
��~ݾ����_��)�;����ݬ���S�
�D_B�`���;�   �   �x�2�bT���q��%�$V�B����͚�߯�� ½�Kѽ�Qݽ7���������3�Δ޽�|ֽA!н�xν:'սEX�B��#�B�L��r��Z��G�оUu �F����2��rI�z[[� �f�jk�2g�M�[���I�6P3����k���R�;�:��o�q��c0�;b���%����N�����n���ֻ �}��   �   �~���oмq��L������;������}|ڽ���\�yu���
������
��d��������ïݽ��Ͻ�Ľm7���*½�UѽW��N����6��i��T��\���A�R	�f����3�!�C��2N���Q���N���D���4��� �w@
��D�nع��z��#�\��`"�
:潈o����J�2b�������!W��YS��   �   �(�j7�uou�Ǟ��|Žfo�g��ψ�3$%�U�-�
�1�92�sc.���'��s�׶�2��1�����Њ˽JP���k��S���������н�G��U2�גI��D����;ƾnF��	��M�6)��L2���5�	�2��r*������`~��ɾL����F���F��\�zԽ_���J��
��q˼�]����̼�   �   7�U�����|���E��t����%� =���P�=H_���g���i�>�e��\��N�H>���+�J��hT��&j˽�r��4��bM������k�����ҽ !��(�(�V��׆�bѥ�K�ƾ��;�����
l��f�Z�k��~���2�;;�A��
ڍ��b��/����LkĽ�����\O����F�m*
�%��   �   �Ԛ�]�Ƚ����]%��@�B�`��P~�
q���"��4����q�������ǋ��.dg��K���/�h��-��r!ѽ�⮽�����2��{Ä�R���v;��D�Խ���yo-�NZ��]�� ���=��) Ӿ�0���[P�����h-뾺>ھ�sľë����JFr��D�;�?����&h��$\���9���1��JD�w�p��   �   K5ҽ!���*��R���|�F���3��n����.����ľˋþ�E�������؟�%d���t���M��G*�aN
���ݽ ��������q��]��'e��$��S���0ҽT���*��R�,�|�uC���0��e����+����ľ�þ(C��8�ן��b��v	t���M�|F*��M
�`�ݽ���������q���]�X,e��'�����   �   n���r-��QZ�$`������@��hӾ�3�a��S��Z���d0�UAھ#vľ�ī�8��0Hr��D��;�������rg���\���9�S�1�GED��p��К�|�Ƚ�����!��@�̒`��K~�xn��  ������xo�������ŋ�S����ag��K�h�/��������!ѽO㮽�����4���ń������>��U�Խ�   �   ��(�{�V��ن��ӥ��ƾP��� �o���m��h��[������4��;\C��ۍ�� b�њ/���SkĽ����ZO����B��%
�t�$�h�U������������0����%�	=�W�P��C_���g���i���e�т\���N�M>�9�+�]���S��꽐j˽�s�����8O��򂝽9���c�ҽJ#��   �   ��I�fF��"��� ƾTI�A�	�`O��7)��N2���5���2�\t*�����3���ɾH����G��^F�.]�zԽ�^��#J�� 
��k˼V����̼�"���6��gu�z��wŽ�i�F������ %��-��1��2�a.���'�*r�ֵ���
1�����z�˽jQ��-m��=��������н	K���4��   �   �i�(V��^��_D��S	������3���C�m4N���Q�P�N��D�:�4��� �IA
��E�Kٹ�{����\�'a"�:�0o��C�J�h^�������W�$KS��u��*eм?����K�����7��۳���wڽ��aZ�>s���
����J�
��c�p�������0�ݽ��Ͻ=�Ľ�8���,½Xѽ�� ��	�6��   �   t������оjv �����2�"tI��\[���f��	k�X3g�|�[���I�Q3�<��Q����;�:����q��c0�b��|%��g�N�^���m�pmֻЬ}�pշ�t�2�4K��.g�%��V�≃��ʚ��ۯ�<½�Hѽ"Oݽ�4�F콸������@3�a�޽�}ֽk"н�yν�(սYZ�\C�#�2�L��   �   _�����5m� b��
'�71B���Z�Z�m��mz���~���z� n���Z��B��h&�b
��~ݾ ���_���;����ܬ�=�S�<弼XB���� ;�";��O��Qۻ��m�xH¼==
�ٹ4���^�ʝ�����ާ�ٖ��OtŽ�0ѽuڽ���7�,��=��)ݽ�ڽ�4۽	��v����9�(�0���]��   �   �Z�������%d�
t/���K�$�e�^�y�jr��!����v��b�y�~]e��xK�m.�������'³��ᆾ�SC�:���*��ԲW�H�⼐+��X�9pa�;�R�;���;��:p�ŻVe�j໼P����,�D%T���z�Z�����ⲽ�½/Ͻqٽ�U�v�㽾��"�:��֮㽪���&�H7�P59�W�h��   �   �X��r�����Y2��RO��Mi�C�}������⇿������}��i��N�421�o��ZK��k��ˈ�F�E��G	�f��w@Y�&.� �#� 4�:@^�;Dx<hY�;�?;p�S���0�����Z7꼣!��sC��kj��a��L���ଽdF����˽B"׽p>߽���I����㽞V�F��1��*�����*<��sl��   �   FZ��K�����c�Os/���K�0�e�V�y��q������5v��\�y��\e��wK��l.�_��Ƚ�k���ᆾ�RC�����)����W����+� ��9�c�;�T�; ��;��:(�ŻXUe�໼��k�,��$T�H�z������ⲽT½h.ϽTpٽ�Tདྷ��Ǯ�$�8��ϭ㽔��8&��6��49�]�h��   �   �]����Pk��`��	'��/B�ӎZ�b�m�vkz���~���z�-n��Z�B�ag&�A
��|ݾ����^��v�;�j���ڬ��S����SB����#;p�";��O��Oۻ��m��G¼�<
�g�4��^�_���r��zݧ����QsŽ�/ѽ�sڽS�དྷ�j��;��'ݽ�ڽ�2۽���8���@8���0��]��   �   `r�����~�о�t ������2��qI�FZ[���f��k�0g���[�)�I��N3�Z��3���r�;�8����q��a0��^��7#��#�N���뼌�m�dֻ��}�Hз�|�2�^J��nf�%�V�����ʚ�ۯ��½�GѽNݽ{3潪
�������U���0�ڒ޽�zֽ�н5wν&ս8W轒A�d#���L��   �   �i��S��[���@徚Q	�M����3���C�1N�9�Q��N��D�E�4��� �?
�BB�Tֹ��x��M�\��^"�F6�ll��X�J��X��؍��4W� GS�<t���cм���x�K�y����6��}���wڽS��Y��r�H�
���T�
��b�0��0���	�"�ݽg�Ͻ�Ľ�5��)½KTѽˎ�v����6��   �   L�I��C������ƾfD�c�	�'L�a4)�K2�ݧ5��2��p*�������a{��ɾ�E���F�TZ��uԽ�[���J���	�Lg˼
S����̼#"� �6��fu�8�nwŽLi���I��� %���-�u�1��2�<`.���'��p�{����-�����˽�M���i��e���詷���нlE��1��   �   <(��V�Rֆ��ϥ�-�ƾ��������<j�
e�2X��~����L/�Ի;Z?���׍��b���/�1��	gĽ𐎽1VO����K@�V$
�N�$���U�,���J���I������%��=��P��C_�V�g�B�i���e��\�z�N�>�ڰ+����PR�l�
g˽5p�����CK���~��K�����ҽ���   �   2��Qm-�NKZ�2\������8;��S�ҾT-�o�L��n����)�P;ھ�pľ<���l��Br��D�8�.�����ld��s\���9�&�1��CD�ݑp��К�*�Ƚ�����!��@���`��K~�[n�����n���6o��E���?ŋ�Ԫ���`g���K���/���J�� ѽ�߮�T����0��Y��� ���9��w�Խ�   �   j-ҽJ����*���R�`�|�6A��B.������k(��N�ľ��þ�?��%�1ԟ�`���t��M�C*��J
�w�ݽP���ӳ���q�)�]��%e��#�����[0ҽ-����*���R��|�fC���0��O���g+��d�ľ��þ�B���򯾛֟�b��Mt���M�E*�[L
�>�ݽJ���*���qq���]�<#e�0"���	���   �   �͚�͖ȽA���'�{@��`�AG~��k��S��Ԉ���l��������ר��]g���K���/����6
���ѽ?߮�T���61��9�s����:��ӤԽ���Vo-��MZ��]��  ���=�� Ӿo0���9P�����--�o>ھ�sľ�«�e��,Er�ED��9�{��-�� e���\���9�Q�1��@D��p��   �    �U�R�����Ѥ�\����%�K=�2�P��?_��g��i�	�e�S~\�O�N�p>���+�C��,Q��
�Lf˽
p��	���K���������f�ҽ� �ʀ(��V��׆�Xѥ�B�ƾ��6�����l��f�Z�U��`��Y2�t�;�A���ٍ��b��/�����hĽ�����VO�����>�"
��$��   �   ��g�6�au����� sŽKd�D��8��U%�`�-�:�1��	2�t].�B�'��n�����J,����཮�˽�M���i�����窷�H�нG��,2���I��D����4ƾhF��	��M� 6)��L2���5���2��r*���{��~���ɾ��~F���F��[�xԽ ]��J���	��e˼�O��v�̼�   �   �n���\м+����K�+����2��4���urڽp�W�Mp��
������
�Za�
������콠�ݽP�Ͻ?�Ľ&6���)½(Uѽ��&����6��i�xT��\���A�|R	�d����3� �C��2N���Q���N���D���4�z� �a@
��D�*ع�?z��y�\�!`"�~8��m��
�J�Z��Z���W��?S��   �   ������2��C��n^��%��V�|����ƚ��ׯ�½FDѽ�Jݽ�0�'����L��;��'0潈�޽{ֽ�н�wν�&ս�W��A��#�,�L��r��S��C�оSu �D����2��rI�z[[� �f�kk�2g�J�[���I�+P3����D���%�;W:����q�c0�a���$���N����`�m�@`ֻ`�}��   �   �";��O��?ۻ�m��A¼^9
�|�4���^�(���0}��Eۧ�󓷽hqŽ&.ѽ[rڽH�����佾;��'ݽ
ڽ�2۽.��l���\8�ȗ0�F�]�^��T���k�a��	'�0B�~�Z�2�m�ilz���~���z�Rn��Z�$B�[h&�
�e~ݾ����_����;�n��Nܬ�ߜS�R�`VB� �� +;�   �   �U�;`��; �:�Ż4Pe��ܻ�:��^�,��"T���z����w���ಽg½�-Ͻ�oٽBT�6��~�����ཪ��b��&�q6�K49��h�Z��&�����c�\s/���K�j�e���y�r��۵���v���y�G]e�wxK�xm.����־�L³��ᆾ�SC�|���*��~�W�&�⼨+��L�9xb�;�   �   ���: ӹ0ʰ�dbK��n����b���?��^�uy�^���Rx��cᖽ���?������}��"���b���ښ��衽�D��Èн���&��]����,�þ ���#�h�J���s�Oʍ�'i���M��W7��bK��}7���B���A���w����r�hAI�0!!��[������$��7S<��@���ڝ��[5� ���j������   �   ����m;��
�nI��j�˼�G��m2��(V���u�b>��㒽�ܚ��;���+��G죽�Т� G�����Ɯ��L���/��u����ͽ�m���Q$��Y�|?�����g����� �ԚG�I�o����sݜ�5����U��[`��b[������Ü�r@����n��F����,����Ϸ�0��4�9����-����4�ȵ����`���   �   �^ǻP�(�jX���%ݼ���1�F���r��<��x/��'���B����������V���{��~����nͤ�䦞����̞�Yj����Ž?u����"�O�ap������T��'�s
>�d�_䄿4w�����������㭿k	������ނ��΄�>�c���<�JW��p�󵯾�~�332�k��nw���}2�8��L9��DŻ�   �   �~��*Y��\P��J;� s��ޕ�����GȽ�C۽ķ�T�FD�S�_s�2�ܽ�aϽ����경�������l*��26��� ��̄�%B���?���Vp��73ݾ�!��/��R��u�~㉿���ם�G���Z���uD���"���gu���R�>�.�{��2پc#��R>m���&��ཷ�����0� �м͂��QX��   �   R���u�(�b�d�X*���`��Y~߽-� �t������!�c+$�ob"�D����B	�LD���:��ɽ�³�r��<����V��t�,hͽ֊��+�Ȓd�-^��rž����R4���;�f�Z��Lv����������%W���t���=w�ߪ[�К<�;��Fc���{þ:X���EW�6'��Ͻ�戽81��D�.	�������   �   t�H��%�����y߽���!�I48�V
K���X���_���`�eK[�xIP�=�@���.�6 ��c�:e齋JȽ.����뛽$y���/��Y:���
�����E����˰����پ���9G"��=�F�T���g�NCt�<�x�n�t��i��WV�ڑ>���#��6�_۾cF���Ɂ��>�b����� 偽�6��`���j���   �   �r��Q�Ľ�;��++�U�@���a���_D��@̔��ߘ��>��m�����c1|�0n`�GC�&&���
����d�������>��'���~���½�����&�(t[��玾 ��������+2�1B�
�L�b�P��eM�ƝC��4��d ��/
��澝���-����_��i&�:���ͬ��z��SA�!},�\�8�g�c��   �   N�н ��p�.��Y�.������׬��缾n�Ǿzs̾��ʾ݉¾���2���Jʏ�r	v��pM��'�	��%�ֽ�������H脽x����[����̽���]�1���g�Br��������۾' ��]��r�0&�dS)��&��B�"��B9����o���)����u��>�>y��Pս������v�yiT�BGU���x������   �   .�M5�'g�$U��Bt���ɾr�⾶������i�{��d���b龘fѾrE���&��?�}���K���,
�� ��䂕��|���o��ك�
��]�ҽJ�xI5�#g�qR��q��E�Ⱦz��}��v���f�n�����S_龿cѾC���$����}�
�K�����������?����|�o�o�B܃������ҽ�   �   ��1���g��t��Ž����۾2
 �-`��t��&��U)�T�&��D����:����q��D+����u�>�z�4Qս����:�v��fT��BU�
�x�����J�н�����.�S{Y����� ��wԬ��㼾ĿǾ�o̾ �ʾ��¾��ʪ��Sȏ�dv�@nM�q�'���*�ֽp��������鄽�≽�^��Z�̽$���   �   �w[��鎾���F�����A�o-2��3B���L��P�;hM���C��!4�df �1
���/���K�����_��j&����ͬ��z�yQA�my,�G�8���c�vn���ĽO5��d'���@���a����}A��Jɔ��ܘ��;�����`���-|�k`��C�Z
&�`�
���zc�������?����������½����S
&��   �   ���������پW��5I"��=���T�b�g��Et�ļx���t��i��YV�z�>�2�#��7��`۾tG���ʁ���>��b�Ɯ��~䁽�6��]��~������H��!��~���s߽���0�!�
08��K��X�6�_�Z�`�kG[��EP�A�@�=�.�Y�fb�xc齚IȽ����6웽2z���1���<��!�����E��   �   �_��Mtž�����5�y�;���Z�Ov����L��㡏�>X���u��P?w�R�[���<����d���|þ�X��BFW�~'��Ͻ戽X61�v?�b�����|�����(�o�d��%��L[��ox߽�� ��� ����!�+($�y_"�������@	��A���8ὶɽu³�*r��৚��W��.󫽈jͽf��(�+�}�d��   �   �q��?5ݾ�"�x /���R��u�䉿
���؝�A���A���BE��V#���hu�ܜR��.���73پ�#���>m���&���8����0��м�ǂ��DX��v��<O���J��C;�us�Nڕ�|����BȽ?۽�轌O�)@��[p�˅ܽ�_Ͻ���&경w���&	��*+��]7���"����⽖C�}�?�����   �   
���
��(��>�l�d�儿�w������i����䭿
��5���N���]΄���c��<�W��p������~�32�����v��?|2����D9�x0Ż�Gǻ��(��P��zݼ�����F���r��9��f,��+���s��	����򼽊��z���ﲽd��-ͤ�����{����̞�dk��p�Ž+w�;����O�pq���   �   ���� ���� ���G�9�o������ݜ�����OV���`���[��G����Ü��@����n��F��������Ϸ������9���
-��4�ŵ�H�� r� $��pM;��
�pD���˼�D��j2��%V���u��<���ᒽ�ۚ��:���*���룽�Т��F����������������u����ͽ8o���R$�a�Y�L@���   �   ��þf �%�#���J��s��ʍ�Si���M��g7��cK��m7��mB���A��lw��R�r��@I�� !�
[��������_R<�4?���ٝ��Y5�^����a���� ��: �ҹHŰ� `K��m���
�pb���?��^�<uy������x���ᖽq��@��򙝽c}�������b��rۚ�,顽|E����н��`�&��]������   �   :��������� �ٚG�:�o�����Mݜ������U���_���Z������TÜ��?����n��F��������η�^���9��	��B,���}4�tõ�8���f� ��pJ;��
�*D����˼�D�tj2��%V���u��<���ᒽ�ۚ�M:��s*��O룽Т�ZF��8��h��������u����ͽn���Q$�u�Y��?���   �   �������&�
>��~d�䄿�v��7������3㭿���楢����J̈́���c�{�<�BV�
o꾕�����~��12����Gu��&z2��꾼�@9� +Ż�Cǻ,�(��O�� ݼ���h�F�V�r��9��%,��ր������������8y���P��̤�����"���c˞��i����Žu������O�Gp���   �   �o��z2ݾ� �F/� �R��u��≿4���֝�M���W���oC���!���eu�L�R�£.�; ��0پ�!���;m���&������ �0��м�Ă��@X�4u��.N��J�{C;�"s�ڕ�G����BȽ�>۽����N�u?���Qo罔�ܽd^Ͻ���貽����?��$)��#5�������⽭A��?�\���   �   d]��qžN���^3�X�;���Z��Jv������������U��ps��K;w���[��<����|`���yþmV���BW��$�H�Ͻ�㈽�21��:������������;�(���d��%��[��Cx߽�� �����x�!��'$�_"�(��:�9@	�@��7��ɽ^����o��s���6U����fͽ��8�+���d��   �   '��������پ����E"���<�Q�T���g��@t���x���t�i�*UV���>���#��4�'\۾	D���ǁ��>��_�ј���ၽ�6�B[��|������H�B!��<����r߽����!��/8��K��X���_��`��F[�dEP���@�x�.�u�ja�Za�TGȽ�����雽9w�� .���8��	佦�{�E��   �   r[�G掾O�����ᾜ��R�)2��.B���L��P�1cM�6�C�l4�}b ��-
����È��ڈ��W�_��f&�]���ɬ��z�iMA��v,�c�8�w�c�n����Ľ5��I'���@���a����kA��2ɔ��ܘ��;��������,|�Aj`��C�\	&�L�
�����`�������<��4�������½���&��   �   @�1�g�zp��r����۾| � \�Xp��&��P)���&�3@����(7�2 㾬l��'��N�u�>�Tv��Kս������v��bT�+@U�3�x������н֠�x�.�<{Y�t��� ��lԬ��㼾��Ǿ�o̾��ʾ{�¾���{����Ǐ��v�QmM�i�'������ֽɬ������/愽hމ��Y����̽���   �   G ��F5��g�\P���n��=�Ⱦ��⾕{��Z���d�6��G��;[��_Ѿ�?���!����}� �K�x��T������>��]
|�E�o�u؃�D	����ҽ�SI5��"g�fR��q��>�Ⱦq��s��n���f�_��t��_�|cѾ�B��^$����}��K�������,�������M|���o�z׃����8�ҽ�   �   ��н�����.��wY�I��E���vѬ��༾*�Ǿl̾W�ʾ��¾~������uŏ�`v��iM���'����ֽ��������儽�މ��Z����̽d��2�1�d�g�6r��������۾$ ��]�~r�+&�^S)���&��B���%9��㾏o��f)����u��>�Dx�aNս:���1�v��bT��>U�E�x�ǟ���   �   Ik���ĽR0��R$�?�@�F�a�����>��UƔ��٘��8�����}��,(|�;f`��C��&�B�
�����^������,<��7���%���½���o&�t[��玾 �������+2�1B�
�L�`�P��eM���C��4��d ��/
����Q���ي��Y�_�i&�g���ˬ��
z��MA��u,��8���c��   �   i�H�U��l���n߽�����!�,8�zK�l�X�Z�_�s�`��B[�WAP���@�\�.���b_�@^�EȽ����蛽�v��I.��C9��;
佉���E����������پ���8G"��=�I�T���g�OCt�=�x�n�t��i��WV�ˑ>���#��6��^۾!F���Ɂ�t�>�ba� ����⁽�6��Z�D{�Ӛ��   �   d�����(�#�d��!���V�� s߽�� �ƙ�����!�p$$��["�!�����=	�%<��4�xɽ�����n��ߤ��
U��D�\gͽ�����+���d�#^��rž����R4���;�f�Z��Lv����������&W���t���=w�ת[�Ě<�*��c���{þX��EW��&���Ͻ�䈽741�;���������   �   �p��
H���E�I>;��s��֕�,���4>Ƚ:۽���*J��:���yk�J�ܽ�[Ͻ����沽�������(���4�� ��9���A�u�?� ��Mp��23ݾ~!��/��R��u��㉿���ם�H���[���vD���"���gu��R�4�.�m�{2پ;#���=m�?�&�%�བ�����0��м8Ă��;X��   �   �:ǻ��(��J���ݼ�����F�%�r��6��!)���}����������E］F��w���첽����ʤ�䤞�����˞��i��p�Ž�t�����O�Xp������R��'�s
>�d�_䄿5w��Ì�������㭿k	������ނ��΄�:�c���<�AW��p�۵����~��22���v���{2��쾼lA9�x'Ż�   �    훹 B;�4�	��A��R�˼�B�h2��"V���u�=;������ٚ��8��)��ꣽϢ�xE��}��Ǜ����������t��F�ͽ�m���Q$��Y�x?������e����� �ӚG�I�o����uݜ�6����U��\`��a[������Ü�q@����n��F����#����Ϸ�"���9�����-���4��ŵ���� n��   �   �^��~��L{ü�n�5o0�IV�	�w�rd����d��nߙ�컗�����D��p���,gt��f��9`��$g��,���Y��N�ͽ�:�	C��뇾Ǫ��~���U(�S$X�UB���-�� ���ѿH��aX��W��W����ѿ����$����[����U��%�{��X�v6z�J�(�m%ٽ߃�kv�~���� ��   �   �(}P�*��^���(�!I�0�q�J}���}���&��$B��.�C�������4������rw���o��[f�;oj�!|���U��;%˽<
�|@��ʅ�r���_����%��T��������/����ο�8�ݚ뿮��S�뿉5��\οe������H��ׄR�*�"�G��j?��"�v��G&��ֽ��ƙ�Vԡ���:��   �   r������5���-��c`��!��P��������ƽ��н6�Խyӽ�#̽�����ݲ�C��������Rmy�r�t�Ʊ�������TĽ���|7��7�Z����k����rrJ�ҡ{��#��s��@�Ŀ>�տ���N��O����տ��Ŀ�S��7˖��xz�x�H�1l�F��"k��Il�9���9Ͻ���Pw�t����䅼�   �   �J�*�,O���<'��e˽�#꽚�?��0�N'��#�px�u������x�ͽ�:���������r!������0���J�������$*�#�k�`f����۾�C���:�:�g��q�� ���H�ſ�ϿTVӿ9�Ͽ��ſA���.���n����g�R�9����TK׾�6����[�PN�*<Ľx�z�P^!�6�伂�˼�   �   O<��Aw�v㡽��ͽ,���:�L*��D;�k[G��xM��LM��G�m�;�,�0�����k��2Ľjj������Uы�����x���b�ὃ\�&�S��8��3Aľ����e&��O��y��Ґ�;ʢ�M�������`��)k���z��7^���T����y��KO��0&��� �tl��̌�r�F�
��j5��:�u��1/�ef�����   �   �ˍ��㹽|,�\��C�6�?SV�-�r������쌾������"D��0��|{j���N��2����b��� �˽�z��\���#*��R@��T�ʽ���)8�/�{�7ĩ���߾����2�NMW�X�z����n��hv���\���ԡ����΍��:|�u�X���3��X�K@�稾 w���/�U:���
��ڜt���D�?�.�]��   �   �oʽ����0*��T������������n���Y5þݜǾ�ž�S��>˯��G��$\��<k���B�����t���5ʽ����?����白ų�p2�Ӫ���S�Q���g���I�X{�T4�r�Q�`l�����Տ����K���hw���On��S�8.6��c�/�ν�������S�a����ٽޞ����y�;�d���y�-횽�   �   BF
��95�|�g��1�������ʾD������H��������8���\��r)Ҿmb��\���ݮ{�P�H��A��������E�����R|��p�½* ���,��7g�X���x�¾�������)�Ħ?���P�
2\�b`��]�b�R���A���,����s�����Ǿ�����n���1����Lg����������*���H����ѽ�   �   ��5�U�n�<����ɽ�;�侷R�Rj��$�j-�>}0�8.��%����<y���F7ž�-��z}�HC����k߽j����Ⓗ0������B�ͽr�R�5���n�L���ƽ���PP��g��$��-�^z0�r.���%����Fw�ҫ뾶4ž�+���}�Z	C�t��D
߽N����㒽�1��s���U�ͽ�t��   �   �;g� ���̠¾��V����)���?���P�E5\�Le`��]�9�R�=�A�˝,�t��H��� �Ǿ�����n��1�8���g�������������Ĺ���ѽ C
��55���g��.��������ʾ���/������J���������x��&Ҿ�_��+�����{���H��?����E���F�����s~����½X, �ғ,��   �   TS���j��&M�}��4�\�Q�1cl�X���������������x��HRn�\�S�06�e�f��%н�����S�!��3�ٽ~���@�y�+�d���y�)隽Vjʽ����,*��T����>���\�������^1þ�Ǿ&�žEP��ȯ�E���Y��8k�
�B���hr��h4ʽ�������B陽vǳ��5�N���S��   �   �Ʃ���߾����2��OW�I�z�/���o��x��h^��֡���[ύ��<|�<�X�G�3��Y��A�	訾jw�V�/��:���
���t�T�D�5?���]�TǍ�N޹��%�}����6�%NV���r������錾������hA���-��Fwj�s�N�+2�z��f���9�˽�y��G����*���A���ʽ����8���{��   �   {Cľ4��tg&��O�^y�Ԑ��ˢ�����x��!b���l��C|��Y_���U��L�y�MO��1&��� �Jm���̌���F�1��5����u�//�yb����bH<�T9w�pޡ���ͽ]}��:6�*�@;��VG�tM�=HM��G�Ϣ;��,�������X罞0Ľ$i�������ы�����3��� ��\^���S�B:���   �   ��۾E�[�:�/ h��r��:����ﵿk�ſS�Ͽ�Wӿe�Ͽ��ſ�A��}/��1o��~�g���9�����K׾�6��ė[�LN��;Ľ��z�	\!��优�˼�@��#��O����S"��� ˽��z����F$�� ��u�(����潭�ͽ�8��~���F���R!������1��5L��y���F&*���k��g���   �   rm����sJ�l�{�x$��t��E�ĿA�տ���9���࿌ ֿT�Ŀ/T���˖�Ryz���H�Yl�f��"k��"l����.9ϽH���Pu������ޅ�d ������,��	-��]`���DL��������ƽ��нi�Խ�ӽ� ̽X���r۲�iA��᱓����ly���t�O�������?VĽ����}7��9������   �   x`��c�%�	�T�{���������R�οI9�k��+�￶���5�	]ο~�����H����R��"���?����v�KG&��ֽ�����С���:�\��(sP����.��U%�x
I�L�q�Q{���{��	%��[@���蛤�����X �����w���o�6\f��oj��|��yV���&˽�<
��@�m˅������   �   �~��aV(��$X��B��.��O ��I�ѿq��yX��W��W�ݷ㿳�ѿI���ـ��A[��A�U���%�?z����a5z�n�(�$ٽރ��t�����, �0W�<�����yü�m��n0��~V���w�kd����d���ߙ�0���w���cE������ht��f��:`��%g��-���Z��]�ͽ<;��	C��쇾x����   �   l_����%�%�T����������~�οc8�y��6��ǡ��4�9\οî��a���G��ރR�V�"���\>��|�v��F&��ֽ���Zϡ�ܦ:���TrP�X�����<%�]
I�=�q�@{���{���$��8@��p����k��� �������v���o�A[f��nj�$|���U���%˽[<
��@��ʅ������   �   rk�ȥ�rJ�W�{�<#���r����Ŀ��տӽ�g��W����տ��Ŀ�R��Vʖ�Lwz��H�k�~���i��)l����F7Ͻ�����s�.��� ݅�V���𘳼t+���-�Y]`����/L������j�ƽ��н*�Խ�ӽa ̽�����ڲ��@��(���?���jy���t� ���/���pTĽ���|7�y7�A����   �   ��۾4C��:�L�g�=q��A���`��ſ��ϿUӿ��Ͽ`�ſ�?���-���m���~g���9�1��8I׾�4���[�bL�9ĽE�z��Y!����J�˼V?�o#��O����2"��� ˽��f������$�� ��u�~���@����ͽ�7��[�������M���/���I��8���$*���k��e���   �   4@ľ
���d&��O�Dy��ѐ�ɢ������_���i��oy���\��xS��B�y��IO�/&�k� �#j��Lʌ���F����1��+�u�,/�q`�o���G<��8w�Aޡ���ͽ:}��-6�*�@;��VG��sM�HM��G�|�;��,�%����$�H/Ľ�g��C����ϋ�<��,����ώ[�$�S��7���   �   �©���߾��9�2�|KW�$�z�P���l���t��[���ҡ����̍��7|�ձX���3��V�B=ྟ䨾lw���/��5������t�
�D�?�4�]��ƍ��ݹ��%�f����6�NV���r������錾�������FA��v-���vj���N��2����������˽�w�����8(���>����ʽ����8�o�{��   �   �O��f��&G��y�n4�+�Q�a]l�2���<���Z�������u��xLn�-�S��+6�ca��{�˽������S�}��
�ٽޚ��=�y�d���y�i蚽�iʽ����,*��T����8���V�������U1þ֘Ǿ�ž%P���ǯ��D���Y���7k�b�B�E���p��~2ʽы������噽ó�0�\��̟S��   �   5g���"�¾�������)�8�?���P��.\��^`��]�4�R���A��,�<��L�����Ǿ����a�n�:�1�����b��q�������������� ѽ�B
��55�e�g��.������~�ʾ���*������D���������S���%Ҿq_��螙��{�1�H�0?������fC�����$z����½�( ���,��   �   ��5�V�n�&���Tý����ON�\e�<$��-�ww0���-���%�����t����1ž�(���}�VC�8���߽Ʌ���ߒ��-�����@�ͽ�q��5���n�@���ƽ���PP��g��$��-�Zz0�l.�x�%����3w����{4žr+��}��C����J߽އ�������-�����H�ͽ4p��   �   �@
��25���g�t,�������ʾ�������r��А���������!Ҿ�[�����>�{���H�m<� ��d����A�����Xz���½�) �k�,��7g�H���n�¾�������)�Ŧ?���P�
2\�b`��]�[�R���A���,����A�����Ǿ:���+�n� �1����#e��Ά�����j������H	ѽ�   �   zfʽ/���)*�	T�l��h����������|-þܔǾ�žRL��]į��A���V��A3k���B�N��El��F/ʽ����ŭ��i噽fó�T1�u����S�Q���g���I�V{�S4�t�Q�`l�����֏����K���fw���On��S�*.6��c� �Sν������S������ٽ����z�y��d�(�y�.暽�   �   .č�Gڹ�� �T����6��IV�s�r������挾怐��P>���*���qj���N��2����M����˽ru��j���P'��Z>����ʽO���8��{�)ĩ�~�߾����2�OMW�Z�z����	n��jv���\���ԡ����΍�z:|�j�X���3��X�!@��樾�w��/��8�����ϗt� �D�J?���]��   �   �C<�3w��ڡ���ͽ�w���2�B*��;;�NRG�_oM�zCM�4G�a�;��,����\�����+Ľ�d��^���L΋��~������\��.\��S�w8��*Aľ����e&��O��y��Ґ�<ʢ�O�������`��)k���z��7^���T����y��KO��0&��� �Ll���ˌ���F�x���3��A�u��,/��_����   �   �9꼌�@O�H��7��"�ʽg�y�֔���� ����r�7��������ͽ�4�������p��K���t.��jI��<���N$*���k�Tf��~�۾�C���:�8�g��q�����J�ſ�ϿWVӿ=�Ͽ��ſA���.���n����g�L�9�|��8K׾`6��4�[��M�;Ľ��z��Z!���l�˼�   �   ����`���0%���-�cX`����H����x�ƽv�н�Խ�ӽ�̽p����ײ�,>�� ���}��0hy���t�T��������SĽZ���{7�w7�R����k����qrJ�ԡ{��#��s��C�Ŀ?�տ���O��Q����տ��Ŀ�S��5˖��xz�s�H�)l�4��k��l����&9Ͻ,����t������ۅ��   �   8���oP�������#��I�"�q��y���y���"��/>��g짽��������j���F���vu��ٶo�iYf�Imj�j{��U���$˽�;
�j@��ʅ�n���_����%�
�T��������/����ο�8�ޚ뿯��T�뿊5��\οe������H��քR�'�"�@��_?���v��G&���ֽ4􂽔�� ѡ� �:��   �   ��6���8{߼#]��7D�ϲq������z��Fd���Գ�J���d������T��LH����z��%]��F��<�;cG���n����%x��"�fk�ʗ������6"�P�W��s��;���{ͿS��HM�����-�����,�®���0�%�̿x�������T�<����렾��Y�d�1���mXW��% ������   �   Ƥ���ü]��D.�_�k)��N؞�h����q���ǽwȽ�ý����&.��:��. ���dn��S��NF�4M� q�J)���޽5P �~�g��𥾬�`���T��8���먿%@ʿ;"�t5��t����P�
��q���ژ�lɿ�ۧ������\Q�7���y�ㄞ���V�i���E���RX�ړ�\d���   �   ��鼼��~F<��"t���������ҽ ��@����5��W����R����ؽ}��D���8����#|��#c�E_���x�6����׽���p�]�=?��*�ݾ���i�I�|������W���}S߿cK��������9������y^��g#߿w`��??���̀�5�G�\h�p1ؾ:���i�M���������[�IN��I��   �   �-0�=^�񙏽�;��ړ߽�/����O�%��0�5�O?4���-�/�"�J�������XQ��G��´��XO��샽�)��P�ͽ�&�Z�M�'H��H�̾D��:�=o������'���nοUi��)�����A� $�������/�ο'!��WC��e&n��8��
��$Ⱦ8���u)@�� �li��Ec�H�*��w��   �   �2�������׽�;�g$�`j@���Y��n�i�|�2Z��A��&`v��_e��'O���5��%��j���Խ��t���MW���-��Mý�;�N�9�`1�� ��t�����%�U�3���Ia���⸿gϿ
+�ک�	��)�D��46п%���pϟ��ᄿ�CU��;%�����ϳ���}���.�$���x��,q�x�O�a Y��   �   A������Ǳ��8C���k����T����⩾�z��g���W��4����ܠ��w��ǲ{� U�ҙ/�H���㽊O���D��齡��|�����_�#���d�����*ؾ�M�Nh8�V�e�����Y��Z���ÿ$�Ϳ�jѿOEο��Ŀ%���Z��)Ԋ��f���8��h�xP׾�����<_�o�;�ڽ]�����h���*ȕ��   �   J���+��[�����x���`��b�ؾ���n����������2���ݾ@bƾL׫��d���k�-�;�|y���,#���k��H���/sֽ�i�x�A�-x��������/�
@�$Bg������[�����3A��qi���ɭ�%���≘��Ƈ�>ui�;�A�����(��r���?��1	�ZZɽ����N8������˽�   �   �1���h����kH���L߾T@�W���] ��()�Ɂ,�Z*��%"�:v�V<������d���u��=�>3����Kh����4*�����̊ ��?Z�h.��\¾���*{�f;��bZ��v�����2������[����ꆿ�wx��]�,>����j���K�žR���V�]��"�r������� ���Ͻ`o��   �   �;h�PƘ���þn�����g+��MA���R�o+^��ob�j$_�X�T�3�C��=.���������Tɾ?�����p���4��m��@ҽ����<�����˽k&�ؓ-�7h�VØ�,�þ�������d+�<JA� �R��'^�lb�� _��T�>�C�J;.����Q���0RɾV����p��4��l�@ҽc���0����˽�(�C�-��   �   1��g_¾.����}�i;�CfZ�iv�����>������M����솿�zx��]��>����D���c�žǾ��:�]��"�8�ｉ����쥽�����Ͻxl��1���h�i����D��H߾�=�t��|Z ��%)��~,�N*�$#"��s�$:���/��&���7�u���=��1�o��(h��2���,����𽕍 ��CZ��   �   ���6��q1��@�mEg������]��9���YC���k���˭��������ȇ��wi�#�A����;����s��"�?�32	�&Zɽn��� 6������ʽ����+�ͨ[�����ʓ��(����ؾ���E����������.��ݾ�^ƾSԫ�7b��[�k�|�;��w��8"���k�������uֽ
l���A�Jz���   �   	ؾyO��j8�7�e�}���[��Z��*�ÿB�Ϳ�lѿGGο��Ŀ�&���[��KՊ���f�N 9��i��Q׾�����=_����ڽ\���	������Dĕ��;���������
4C�Ҩk�£���~��ߩ��v��$c���S������t٠��t��%�{�i�T��/�.�����M��GD��x���0~�����#�&�d�դ���   �   _�����%�t�U������b���丿�hϿ�,�Ы��������῝7пW���kП�gℿ�DU��<%�3���`г���}�,�.�����w���(q��O�=Y�.�����f�׽�7�$��e@���Y�;�n���|�DW��@>���Zv��Ze��#O���5��"��h���Խ��n���2W���.���Ný$=���9��2��Q���   �   ��~
:�8?o������(��pο�j�v+��X���A��$�Ҫ��8���ο�!���C��8'n���8�9 
�%Ⱦg����)@�� ��h���Bc���*�;s��'0��^�q����6��č߽8,���W�%��0��5�f;4���-���"�p�2�����jN��9��z���TN��샽�*��0ν(�x�M��I��P�̾�   �   �����I�[������x����T߿�L��n�����:����b��/_���#߿�`���?���̀�j�G�th�v1ؾ(���&�M�P��Հ����[��K��B漒�鼪��z@<��t����^	��@�ҽ�����3� U�
��E��z�ؽz������~���=!|��"c��D_���x�E ���׽���N�]��@����ݾ�   �   @���T�l9��w쨿�@ʿ
#��5�u����XP�H��0q������!lɿ�ۧ������\Q� ��+y⾄���H�V�ן��D��wPX�����_��������ü��e@.��_�#'���՞�帱�ro���ǽ�tȽ�ýኹ��,����K��~cn�X�S��NF��4M�pq�S*���!޽NQ � �g���
��   �   X7"��W��s������_{Ϳ���lM�����-�����,�������/�ǅ̿�w��(����T�����J렾��Y��c�����vVW�$ �򸦼���0����y߼U\��6D�1�q�����}z��8d���Գ�p�������=U���H����z��&]�.�F�9�<��dG�,�n����ny�Ȏ"�w�k�|�������   �   ����T��8���먿@ʿ"�V5�tt�`���O�����p�,���Wkɿ9ۧ������[Q�\��<x�ۃ��`�V�9��D��YOX�����^��:���@�ü��H@.��_�'���՞�޸��fo��wǽ�tȽ�ý����v,��������bn���S�NF��3M�Pq��)��� ޽�P ��g�����   �   ���+�I�H������������R߿�J��X������8����P��;]��9"߿`_��B>���̀�ɯG�:g��/ؾ爗�k�M���6����[�J�A�Z��Q��5@<��t�𖘽R	��6�ҽ������2�U������+�ؽ�y������ ��� |�A!c�AC_���x�������׽���p�]�4?���ݾ�   �   ��):�=<o�(����&���mο5h�w(�����J@�,#�ۧ����翬�ο��� B��T$n�@�8��
��"Ⱦ����'@�  �ef���?c���*��q��&0�O^�H����6����߽0,�ۨ�N�%��0��5�M;4���-���"�:����I�όM��h�������K�j냽�(����ͽ6&��M��G����̾�   �   2�����%��}U�g���H`���ḿ�eϿl)���%��8�U��Y4пi����͟�C���@AU��9%�(���pͳ�`�}�I�.����<u��T%q��}O��Y�.��?��4�׽�7�$�e@���Y�6�n���|�<W��3>���Zv��Ze�[#O�A�5��"�:h���Խ�������dU��B,���Ký�:�o�9��0��F���   �   �ؾ}L��f8�z�e�����X�����G�ÿ0�Ϳ�hѿ5Cο��Ŀ#���X���Ҋ��f���8��f�xM׾����9_���ĺڽY�����F���pÕ�c;����������3C�èk������~��ߩ��v��c���S������Y٠��t��ҭ{��T��/����΂�ZL��JB��ݻ���z����6�#�k�d������   �   S
��;�ﾙ-�@��?g�<���IZ��@���0?��Wg���ǭ�
��������ć��qi�f�A�Å�X��=ﵾ�p����?��.	��Uɽd����3������ʽ�����+���[�~���Ɠ��(����ؾ���B�����������-��ݾ�^ƾ*ԫ�b����k���;��v���1 ��/i������pֽ�h���A��v���   �   �,���Y¾���Cy��c;��_Z�d v�����@������M����膿�sx�@]�>������ϲž�����]�i"���;����饽���r�Ͻl�һ1�t�h�^����D��H߾�=�v��|Z ��%)��~,�J*�#"��s�:������𿛾��u�%�=�1���Ὓe�������'��ܿ��� �v=Z��   �   �3h�A���p�þ]����	b+�HGA�׻R�,$^�ahb�$_�h�T�оC�(8.��������SNɾ;����p�%�4��i��:ҽ�񲽄���߫˽�%�y�-��6h�DØ�#�þ�������d+�?JA�"�R��'^�lb�� _��T�6�C�>;.�|��*���Rɾ���w�p�V�4��k��=ҽ0�Ķ��ݪ˽�$���-��   �   M�1���h�����A��_D߾�;�����W ��")�p{,�*� "��p�z7�h��4��ۼ����u�{�=�^.����Cc�������'����I� ��?Z�Q.���[¾ެ��){�f;��bZ��v�����3������[����ꆿzwx��]� >����B����ž�����]��"�]��"���%꥽x�����Ͻbj��   �   �����+�٤[�������������ؾ��J�����������(���ݾYZƾ�Ы��^����k��;��s���/��Xg��M���*qֽDi��A�x�����y��/�
@�&Bg������[�� ���5A��ti���ɭ�$���߉���Ƈ�5ui�/�A������񵾾r��a�?��0	��WɽP����3��8��a�ʽ�   �   8��������0C��k�ꠉ�x{��۩��r��_���O�������ՠ��q��.�{�@�T���/����~��H���?��k���z��Q����#���d�����ؾ�M�Nh8�V�e�����Y��]���ÿ'�Ϳ�jѿQEο��Ŀ%���Z��&Ԋ�٥f���8��h�SP׾����<_���F�ڽNZ����H���X����   �   �+�������׽�4��$�Fa@���Y��n�ʏ|�IT��A;��Uv�aUe��O�	�5���Fe�/�ԽQ
��N����S�� +��(Ký;���9�A1����j�����%�U�4���Ja���⸿gϿ+�ݩ���,�E��56п#���oϟ��ᄿ�CU��;%������ϳ�\�}�T�.����v�� &q�z|O��Y��   �   �#0�z^�
���s2����߽<)�}����%��0��5�374���-� �"������&��wI�����د���G��都�'�� �ͽ'&��M�H��<�̾B��:�=o������'���nοWi��)�����A�$�������.�ο&!��UC��a&n��8��
�|$Ⱦ���)@�\ ��g���@c�q�*�&p��   �   ��鼁��O<<�nt�֓�������ҽ^�����]0�tR����:��Ʒؽ�u��)���(���X|�yc�>@_�a�x�����F�׽g��F�]�0?��$�ݾ���h�I�|������X���S߿fK��������9������z^��g#߿y`��??���̀�/�G�Uh�[1ؾ"���(�M�P������S�[��J��?��   �   ����n�üd��0>.�_�u%���Ӟ�����m���ǽ rȽU�ýJ���,*�����4���_n��S��KF��1M�jq��(���޽P �h�g��𥾨�`���T��8���먿$@ʿ<"�t5��t����
P�
��q���ژ�lɿ�ۧ������\Q�4���y�ք����V�@��fE��/QX����h_���   �   {弻� ��b"���P��9��*D��8��_kǽ(�ԽHe۽ؕڽ<�ҽ��Ľu���
f���/����c���E���8��F��y������� �fb@�06��lξ�;��$I�u��� _����ӿ0��.x�n�$��?3��=�Fv@��=��%3�>$�F��d���J=ҿc��������E�.�FZȾ��3��佚a��l�6�}V��   �   � �y�\�8�ol��n��2Ү�E�Ƚ��ݽ�+�*�h��p��*6ٽ�ZĽp_��"����y��|V��HE�S�N��|�0x��a����=����|'˾g��^�E�݉��B����п���6&���!�@D0���9�d1=�J�9�=0�T�!�¿�����?Ͽ6��j���'�B�R���Mž������0�.��я�+�;�x
��   �   �(���H���}���@Ľ���V�������������� -������dݽmǼ�V(�����k��Tg�J���S���y��4`6��ۅ�x���0	��a<�U�z�I�����ƿ��Zr	�J1���'��0���3�:�0���'��=�N	�'��e�ſ\���x�,�9��y��v���O��xO*�c�ݽ�o���8K�%r&��   �   �%o�aO���p����轉.���%��u;�z M���X���]�u�[���R�,~C���/��b����׽0ٱ�09���L���̏��D��t��B +��x�5������~�-��f�K�����g�ۿ���Fg���z�"���%��
#�T����v���ۿ�G�������Ne���+�����4���� o��� �d�ֽ (���g��V��   �   �󪽘�׽~��] *��4M��o��C��ر�����fF���`���{��H����y���X�i7�ؑ�7��1�ƽ����c������׭��p�(�`�愠�ڿ�����N��y���Y��6�Ŀ���K<����
�ب�xA�r��l��0 �>��=]ſ�����U���RM����߾W���LY������Ͻbm��\ǈ��,���   �   ���3h��bD�S�s�Ò�K#������Ҿ�P޾J��@�߾0�վ�9ž?8����������P���&�[K�ֽ֟D����J��m6ڽ����wF��닾 �þ`����1�~e�7[��sɪ��ſ��ݿ%��i>��"� �s����%��^߿�Fǿ�ͫ������e��2��~�=<¾0򉾛AA��`��sʽ��mᦽ ���   �   3%��V�0ሾ����̾�������k�H#�����v�����s�Ҿ�د�-���ha�S/����"z߽{ʽz`Խ��%�+�<�m����m3�f����?�G�n��k��㐦�����)˿��տB�ٿU_ֿZm̿:����������;�p�cA�*��|��N{���*l�S!)�����_9ɽ~7���=Ͻ-~���   �   Z]�{����Q������
��"�J�6��[G��.R�E?V�'S��-I��@9���$�L����v��qZ���)e��R.��)��m��ӽD��J-�JE�9����;���K��:�dA���h�6����s��Cץ������ű�3�����t���w�k�q�C�������&���ч��>F�����潽�ͽ2m׽�b��V'��   �   !菾ȫ���󾖲���6��(U��,p�Xт�'Љ�qk��=a���܃��r�nX��9�HR����9m���U|[�6+$�L��2ڽ��ؽ\����� �J�V�R叾���6�󾼯�{�6��$U��(p� ς��͉�*i��_���ڃ�e�r�>X�o�9�#P�����j��	z[��)$�v���ڽ�ؽB����� �q�V��   �   �>��P�=�>gA�U�h�V���Iv���٥�	���eȱ�r5����q�[��]�k���C�d�����(���҇��?F������� �ͽ�i׽6`�
S'��]�b���N��ʉ�/�
�l"���6� XG��*R�W;V�D#S�*I��=9���$������+s��TX���&e��P.��(�Hm�'�ӽ�꽊/�rME������   �   �6ྴ��v�?���n�n��#���Q��3,˿O�տֈٿ�aֿ�o̿A������(�����p�8A����d�ྍ|��9,l��!)�����
8ɽ�4���9Ͻhx��6/%��V�ވ�����̾l����� �2� � �������Q���~Ҿ�կ�ؓ���da��P/�O���x߽�ʽ�aԽ2���+��m������   �   5��> 2�pe��\��{˪�D�ſ�ݿ����@��h� ������'��`߿FHǿXϫ����<�e� 2�h�b=¾��5BA��`��rʽ�먽ަ�|������>d��]D�R�s�����=��t��L�Ҿ�K޾O��q�߾��վ�5ž�4���|�������P��&��I���ֽd����J��=8ڽX���zF�t틾��þ�   �   ���N�{��F[��$�Ŀ��㿗>����
����B����l��1 ����n^ſꇤ��V���SM�����߾�W���LY����ְϽ�k���Ĉ�)�����׽����*��/M��o�2@��O���w𛾼B��i]��Jx��
E��Y�y�X�X��7���4��}�ƽ����������ۯ㽾r���`�׆������   �   *�-�!�f�QL�������ۿc��Hh�"����"�Ʒ%�r#�&�����w��ўۿXH��:���MOe�N�+�#���w���!o�p� ���ֽ�&���g���V��o��J���k������*���%�@q;��M���X���]���[�0�R�zC�<�/��_�b�@�׽xֱ�o7���K���̏��E������!+���x��������   �   kc<��z�[���5�ƿS��s	�2�f�'�֭0�Z�3���0��'�^>�hN	���쿽�ſ����Xx�K�9��y�wv���O��O*�g�ݽ�n���5K�+n&�6�(���H���}����qĽf��h��}��Z�����ޝ�v*�P���2aݽ|ļ�&��f��@k�lTg�����+T���{���a6�݅����G	��   �   t�E��������ʂп����&�:�!��D0�8�9��1=���9�N=0�z�!�ֿ�����5Ͽ��J�����B����Mž6���T�0��㽘Џ���;��u
�� ��u�i�8��l�|l��oϮ�P�Ƚ��ݽ�(�+�������3ٽ�XĽ�]������o�y��{V��HE�ިN�u�|�Zy���b����=�y���(˾@���   �   p%I�ڲ��o_��I�ӿ���dx���$��?3��=�Fv@��=��%3��=$�������<ҿ���������E��-�jYȾj����3����q`����6�U��x弙� ��a"���P�9���C�����/kǽ�ԽPe۽��ڽ~�ҽ
�Ľ�����f��
0����c��E��8���F��y�֣��M� �fc@��6���lξV<��   �   ��E�����W����п��� &���!�D0�l�9��0=���9��<0�Ԫ!�F������hϿw�������B�~���Lž������0����Ϗ�ی;�Hu
�t �Xu�N�8��l�rl��hϮ�Q�Ƚ��ݽ�(�#�������3ٽ�XĽ�]��͜���y�p{V�HE��N�H�|��x���a���=�����'˾����   �   �a<��z������ƿm�� r	��0� �'�X�0���3�l�0���'�$=�VM	����3�ſS���Xx���9�nx��t���N���M*�}�ݽsm���3K�m&���(�z�H���}����dĽ`��h���z��T�����ϝ�b*�����`ݽ+ļ��%�����# k��Rg������R���y��<`6��ۅ�r���!	��   �   ��-�@�f�~J��W���z�ۿY���f�@����"���%�v	#�J����t��B�ۿ0F��v����Le�2�+����P���/o�s� ���ֽ�$���	g�*�V��o��J��jk��|���*���%�@q;��M���X���]���[��R��yC��/��_�.���׽�ձ��6���J��vˏ��C������+���x�����l����   �   ���N��x���X����Ŀ�㿍:����
����J@�<��<��/ �#��U[ſN����T���PM�4��߾U��hIY�.����Ͻ�i��`È�&(��@6�׽����*��/M��o�2@��P���w𛾺B��c]��Ax���D��0�y�$�X��7�Ў�r�󽉄ƽ����C���k�Y��2p�&�`�0���ξ��   �   n����1��e�Z��Ȫ�U�ſ��ݿ���<���� �����#�\߿]Dǿ�˫�������e�~2��|�p9¾���_>A�^�NoʽR騽�ܦ�������d��]D�E�s�����=��w��N�Ҿ�K޾M��k�߾��վ�5ž�4���|�������P���&��H�.�ֽu���<H��d4ڽ����vF��ꋾ��þ�   �   _1������?���n��j��!������d'˿B�տ��ٿ�\ֿ�j̿Ȉ�����������p�A�ڨ���ྒྷx���&l�)�N���r4ɽw2���7Ͻnw���.%��V��݈����~�̾m����� �3� ���������:���~Ҿ�կ�����;da�%P/�����v߽� ʽ^Խ`���+�(�m������   �   �9��	I�9��aA���h�~����q��ե�,���qñ��0��n��왿{����k�.�C������[#��χ��:F������潆�ͽ�g׽x_��R'�V]�M���N��ŉ�.�
�n"���6�$XG��*R�X;V�B#S�*I��=9���$������s��"X��k&e�P.��'��j�\�ӽ}�꽦+��GE�¤���   �   l㏾����ҋ󾓭���6��!U��$p�͂��ˉ��f���\��D؃�,�r�`X��9�=M�����f��뒾}u[�Q&$�l��wڽz�ؽE���B� ���V�3叾
���.�󾻯�|�6�%U��(p�!ς��͉�,i��_���ڃ�a�r�6X�d�9�P�����j���풾�y[�)$���dڽ۳ؽ����� ���V��   �   B�\�$���K������
��"���6��TG��&R�k7V�OS�7&I��99���$�����o��U���!e��L.��%��g���ӽu��`,��IE�����;���K��:�dA���h�8����s��Gץ������ű�3�����r���n�k�e�C�������&��Zч��=F�������N�ͽ�f׽R^��P'��   �   c,%�P~V��ۈ�� ����̾���}��������������������yҾ�ѯ�����K_a�bL/�����r߽[�ɽ�\Խw�c�+�Ĩm�����Z3�b����?�I�n��k��否�����)˿��տE�ٿW_ֿ[m̿7����������2�p�XA���W��{��$*l�m )�����5ɽ+2��A6Ͻ)t���   �   �~�Ca�%ZD�y�s��������l��ӧҾ�F޾N��k�߾ԕվR1ž�0��Ny�������P���&� F�ȗֽh���]F���3ڽ���awF�T닾�þZ����1�|e�8[��tɪ��ſ��ݿ'��l>��$� �v����%��^߿�Fǿ�ͫ����{�e��2�w~�<¾���@A��_��pʽt騽rۦ�����   �   J몽�׽���:*�&+M��o�6=������웾?���Y���t���A��.�y���X�-7�!������ƽN���ه���񲽣��Bp���`�Ą��ʿ�����N��y���Y��7�Ŀ���L<����
�ڨ�zA�r��n��0 �>��<]ſ�����U���RM�����߾�V���KY����b�Ͻ	j����d&���   �   �o��G��xg��z�轼'��}%�m;��M���X���]�s�[�.�R�XuC���/��[���q�׽�ѱ�>3��H���ɏ�>B�����+�x�������}�-��f�K�����i�ۿ���Fg���z�"���%��
#�T����v���ۿ�G�������Ne���+�������� o�� ���ֽ�%��:	g��V��   �   s�(��H���}�����Ľ�����'�k��&��R�����p'�����%\ݽ���4"����^�j�Og�'����Q���x���_6��ۅ�j���-	��a<�U�z�J�����ƿ���Zr	�J1���'��0���3�:�0���'��=�N	�(��c�ſZ���x�&�9�zy�qv���O��O*�V�ݽgn��a4K�Dl&��   �    �At�w�8�Sl��j��hͮ��Ƚ�ݽ�%��c�����0ٽ�UĽ5[�������y� xV�EE�{�N���|�pw���`��n�=����v'˾f��_�E�݉��B����п���6&���!�@D0���9�d1=�L�9�=0�V�!�¿�����?Ͽ7��i���&�B�O���Mž������0��� я���;��u
��   �   �!��.���T�\ℽ�����5��y۽���<��4�����X��a�彺�ͽ�β�{���%|�+W���G��qX�������ƽ���Ib�M��������o/��q�E��g�̿����*���/�؈F�P�Y���f�.�k�T�f���Y��F���.�H&�"���&�ʿ9\��� n��v,�`]�٣��X�j��+W��#�l�1/��   �   "�-�D�B�/o�����P���Dֽh�	��Ro�����\�
B	�^=���㽋�Ž�&��l ��xk���V��Yb��)����ƽ�&��_��0��̼򾎘,�c�m�˴��A�ɿ��������,�C�:�U��b�d;g���b���U���B�\,��������z�ǿ�훿�ij���)���Cs����U��
�������r��9��   �   ��\����O韽L`ƽ-/𽄶��G�S0.�� 8��8<�#:�d
2�S�$����5 ��aؽ[��l㔽N���h������qǽ�[�ipV�*Ӟ��`�[$�Ab�XA���A���M����Z$��B9���J�\mV�B�Z�x�V�j�J��R9�l'$�@E�1
�r׾�6ה�Ҙ_�E�!����=���z�M�B���J�����Y�Y��   �   7*��.ɷ����z��)+�M�G��Ya���u�vÁ��w���҂���y�� g�W�N�+a3����q��A�ʽ���?	���d���ɽ��
�TcI�2}���վ���P�v�������[ۿ"�����<q*�$�9�"AD�H�4�D��h:�.�*����x����ڿ�ư�٭����N�����Ҿp܏���A�#�����푽�����   �   �ӽW$�j&���M�puw�{"���|��=0��-຾v��� ���q��;���9����<�V���/��*�b��޸½	����;Ͻ-���9�$a������2T��:�e�w�bҞ�_�Ŀ�����`J�t�%��}.��1���.�*^&����h���-�ĿV�����v�P�8�q���������x3���������T1��J ���   �   Ua�6
;�I!m�?㒾������;+辖/��8~�f��/�����H��FҾ�9���{��,v���C��O�b����ڽX�ڽ� �]�(�2�k����b�� �h�U�0���߆��_̿�$��I�,����"������v�v:����WͿ%K���މ��	V�3q ��*龁d����g��>$�R����ν��̽���   �   �iG�^C��(ؤ��̾������n*"���0�o:�s	>��H;��k2��G$�X1������ѾC���<���uN�� �,�Pr���������L��ݍ�wž���3��nf��2��ʫ��ǿ46߿[L�%���n��f������e"��ȿIQ��IO����g��3�[���ž�A��uJ�t�:$�a�~��۞��   �   +߄����6߾��
�UV'��C���[�̜o��y|�L���7�}�<�q�q^���E�6*��S�8g㾇���r䇾�1N���K��-�����j�/��k��I��#�ھG��:�B�h�}׋�su���r���=ƿ��п,WԿSѿw�ǿ�7���?���m��k�+�<��`��lܾ4��5sl��4/��J
�?��g����tDI��   �   ɬ�������6�*\���%$���ڜ�� ���5��˥�����������V	_�L69�,���I��2������]C�����7���E���@�`À��Ŭ���P���6�'\�����!��B؜�-���2��}ȥ���ͨ������ _��39�)���F羵0��E����C�a��1�t��)H��@��ŀ��   �   ��ھ��F�:��h��ً��w���u���@ƿ��пZԿ�Uѿ�ǿ::���A��Co���k�Z�<�#b��nܾ�5���tl��5/��J
�=�������P@I�X܄�G���	߾��
��R'�
C�@�[�;�o��t|�������}� �q�?m^�i�E�l*��Q��c�󸱾�⇾X/N�۵����P�����	�/��k�ZL���   �   7��C	3�rf��4��i̫�oǿ9߿dO�=������S���Y���$�"�ȿS���P���g���3����dž�B���uJ�z��"�^�Jy��w��HeG�`@��^Ԥ�n�̾��������&"���0�(k:��>�	E;�h2��D$��.����� �Ѿ<@���:���rN�1� �@�6r�(��������L��ߍ��ž�   �   G� �B�U�򆉿�����̿u'�FK����"����,��@x��;���YͿvL���߉�WV�Er �,�Xe��w�g��>$�3�����ν�̽��꽼]��;�fm��ߒ�t�����;�%��)��6{�b�-����_��ҾF6���x���v�B�C�;M�����|ڽ��ڽ� �Q�(�S�k�m���e��   �   �:�*�w�Ԟ�^�Ŀ��T���K��%�.���1�\�.�d_&����i�n��J�Ŀ1����v�0�8������@����x3��������T.����ӽ� ��e&�d�M�(ow�����x���+���ۺ�����
���m�����������V�6�/�,(�����½{���f<ϽQ���9��b������U��   �   �P����������]ۿ&��ң�~r*�~�9��BD�^H�j�D��i:��*���� ����ڿGǰ�E�����N����Ҿ�܏���A��"�V��P둽|���&&��ķ�1�彳�%+�L�G�HTa���u�m����t��Ђ�<�y��g��N��]3���m����ʽV���&���d��&�ɽ�
�ReI��~��9�վ����   �   �Bb�fB���B��
O�V���[$��C9���J�rnV�H�Z�^�V�&�J��S9��'$��E��
쿹׾�_ה���_�P�!��������M����oI�����ƟY�?�\�@��(埽][ƽ�)�V��	D��,.�8�,5<��:�2�G�$�@���3 �^ؽ���~ᔽ�L���h��&���rǽ�\�7rV��Ԟ��b�j\$��   �   ��m�����*�ɿ����F����,��C���U���b��;g�,�b�J�U��B�t,��������^�ǿ�훿=ij�]�)�����r��	�U�j�
�T�����r��9���-�Q�B�|*o�Z���`���ֽ�d�:��|m�+��"[�~@	��:����㽡�Ž<%��f���vk�%�V�RZb��*���ƽ�'�_��1��O�򾒙,��   �   N�q��E����̿���n��/��F���Y���f�.�k�:�f���Y��F�H�.�&�������ʿ�[���n��u,�^\�Vأ��X�����U��-�l��/�1 �i.���T��ᄽ ���D5��(۽~��q<��7�����������2�ͽQϲ����&|��W�!�G�7sX�
�����ƽ���vb���������p/��   �   ��m�ﴝ�Z�ɿ���������,��C���U�n�b��:g��b�R�U�.�B��,���������ǿ6훿Jhj���)����&r��(�U���
������r�n�9�\�-��B�^*o�N���[���ֽ�d�>��|m�*�� [�x@	��:����㽊�Ž%��>��jvk���V��Yb�*��2�ƽ�&�$_�	1��K��٘,��   �   �@b�*A��VA��$M�2��rZ$�*B9�ԩJ�vlV�>�Z�h�V�\�J��Q9��&$�tD���;־�/֔�(�_���!����ӆ��\�M�����G�������Y���\�
��埽U[ƽ|)�W��D��,.�8�+5<��:��2�>�$�/��l3 ��]ؽS��ᔽbL���g����Iqǽ�[�tpV�1Ӟ��`�
[$��   �   T�P����c���#[ۿ������Zp*��9��?D��	H�ؗD�Jg:���*����z���ڿ0Ű�������N���UҾ�ڏ�w�A�!�L���鑽�����%���÷��彪�%+�K�G�NTa���u�p����t��	Ђ�4�y��g���N�g]3�m��l��_�ʽ������@c���ɽd�
��bI��|����վ����   �   �:��w�ў�8�Ŀ`��,��PI�6�%�(|.���1�v�.��\&�P�fg�ǅ�7�Ŀ�����v�*�8�������&����u3�D��������,��%���ӽ� ��e&�]�M�'ow�����x�� ,���ۺ�����
���m������	�����V���/��'�(�佰�½�����9ϽX
�ȋ9��`��桿��S��   �   �� ���U�"��������̿�"쿬H�ڠ�����(��fu�9�r��UͿI���܉��V��n �H'�b����g��;$�#�����νP�̽���j]�X;�Om��ߒ�s�����;�%��)��8{�c�-����W���Ҿ16���x��qv��C��L�7���}	ڽ́ڽ� �!�(���k���a��   �   ���3�elf�%1��Hȫ��ǿ�3߿�I�?�����Q�������d�ȿ�N��9M��`�g�D�3�6���ž+?��CqJ�\����[佌w�����dG�H@��SԤ�j�̾��������&"���0�,k:��>�	E;�h2��D$��.�k����Ѿ@���:��frN�� �<�6o�Ǖ��q��ޏL��܍��ž�   �   ��ھ����:�r�h��Ջ�hs��}p��;ƿ��пBTԿ!Pѿ��ǿ5��'=��Fk��5k���<��]��hܾ1���nl�81/��G
�9��:��F���?I�2܄�3��w	߾��
��R'�C�C�[�@�o��t|�������}���q�<m^�b�E�c*��Q��c�ʸ��j⇾�.N������������/���k��G���   �   `ì�~	�H����6���[�������՜����90���ť�s
��K���J���_�:09�O��B�.-�������C���
�`���D�ס@�&À��Ŭ���N���6�)\�����!��E؜�3���2��ȥ���̨������_��39���jF羁0�������C���B����D�.�@������   �   [ڄ�����߾��
�'P'��C�x�[��o�bp|�������}�h�q��h^�v�E��*��N��^�����߇��*N������T}����`�/�u�k�WI���ھA��:�D�h�׋�uu���r���=ƿÃп.WԿSѿw�ǿ�7���?���m��k� �<�u`��lܾ�3��prl��3/�I
�:��κ����c=I��   �   �aG�(>��vѤ���̾�������#"���0�qg:��>�'A;�Id2�A$�d+�ߊ��:ѾR<���7���mN�-� ���Wl�t������ΐL��ݍ�Sž��~3��nf��2��
ʫ��ǿ76߿_L�)���p��i������d"�
�ȿEQ��EO����g���3�H���žLA��tJ�� �q[佀u������   �   [�;��m��ܒ�檰���;� �a$��Ox�`�*�7�����	Ҿ�1��u���v�C�C�0I�����ڽ�ڽB �F�(���k�����b�� �f�U�/���ᆪ�a̿�$��I�.����"������v�v:����WͿ#K���މ��	V�%q �u*�Dd����g��=$����(�ν��̽����   �   ӽ$�Eb&��M��iw����Xu��(��׺�����i���i������l꓾<��k�V���/�T$���佞�½ƶ���7Ͻ�	�ۋ9��`������*T��:�e�w�cҞ�_�Ŀ�����bJ�t�%��}.� �1���.�*^&����h���*�ĿS�����v�H�8�c����������w3�X���<���,�����   �   T#��U���b�彴�u!+���G�\Oa�6�u������q���̂�H�y�g���N��X3���bf��?�ʽ�������`��b�ɽ��
��bI�}����վ���P�v�������[ۿ$�����>q*�&�9�$AD�
H�6�D��h:�.�*����x����ڿ�ư�֭���N����rҾ=܏�Z�A�"�8���鑽h����   �   �\���<⟽�Wƽ%𽬰��@�A).�w8�d1<��:�D2���$�����0 ��Xؽ"���ݔ��I���e��F���oǽ�Z�
pV�Ӟ��`�[$�Ab�XA���A���M����Z$��B9���J�^mV�B�Z�z�V�j�J��R9�j'$�@E�0
�r׾�5ה�͘_�?�!��������M����I��*����Y��   �   ̏-���B�(o�����j����ֽ�a�~��k�V��DY��>	�7��c�㽌�Žv"�����grk��V��Vb��(����ƽ>&�^_��0��Ƽ򾎘,�d�m�˴��A�ɿ��������,�C�:�U��b�f;g���b���U���B�\,��������w�ǿ�훿�ij���)���4s����U���
�λ��I�r�Ą9��   �   �VF��>X�H큽p�������C�� �_����-�vV�������]�t�˽�$����^ q��}_�-�r�Tx���⽻�*�큾��¾��-�K�V)���������x!�Th/�P�M�F�j����������������� ?j���L��?.�����t�뉷�1h��r�H�Ԡ�[达��|�YN$�,Kս�⏽_�Y��   �   ��W���o�m쐽����ֽ�]��W��9�w�#�`_'�K%�D������M��w�r����
���K��U�p��C~�Vs���'�'g)�T5����������wH�i艿����������,���I��Sf�j�~�����������b�~���e�h(I�,�+� �����E���B��ٸE��q
�����xy�M�"���ս���~Qe��   �   \����ݛ�s㾽���(�4c$�Nd9��.J�J?U���Y��V�rM��^=��?)���W��R˽�9��:咽�ې�{Ψ�J
��-%�S�v�7w��� �y�>�m\��"���Q޿�	�d0$�.�?��Y��%p��q������mp�(�Y�L?�>�#�R^��ܿ���X���}�<�����-p�� ��'׽�ڜ������   �   �۴��2ڽ�\�O�&���G�Ѓh��=���b���U���;���G��(����m��M��,�ח����9���pԯ��������
!��g��X��w���v0� Br�����-wͿ�w���z��	0�nG��Z���g��l��Bh��.[��G��T0� q�����I�̿[ß��Rp��:.������e���b�x��j۽Ԇ��f@���   �   &��X'���B��p�k�� ���\Ἶ��;��ؾ�!ݾX�پ�ϾK}�������_��Ǵv��I��M!��[���ݽ(�ӽ9	�)��څU���@޾80��AX�S���(���2㿎���!�v�0�LA�L��7P�
�L��B���1�����bp��ͷ�ZA���*W�R���۾\×�s Q�v ��k�z�ɽ�#ӽ�   �   �I+�+QZ�P/�����$�;R����l>��3�?,�+��s�έ�XR��Ѿ@���S����`�Y�0�}������ġ���-��iB�p���v��h��:�åx�����kiſ���j����bj&��[/���2���/��n'�(��g	� R��Cƿ�럿��x���:������(����?�����������	��   �   Lh�������~w�2���o'�ڿ<�x�M��X���\���Y�FO�.�>���)����8��̓þP�����m���8�����NL��h0�^l��M��P�便���:P�mᅿ�����ƿ�(濣� ����2;�B��8��j����C�̐ȿHJ��U���FQ�y��x���ɣ��j��A.�F���d�t��fZ4��   �   M���ʾ��B�!�l�B��c����+��狒��H�����o0��$ ��>�e�ՁE� $�����;t䜾ͫm�j�7�.��(��@!�VK����l/���Y����(�7SY��$��C���0���ӿ#'�����U����Z��9տ'��.���Mt���.[�*�����5�N҈�R�J��V �������Q&5���i��   �   [�Ⱦ����*�4�T���������.��'����2����¿)￿���!Ҩ�mq���v���W���,�6#�)�ʾ�ޖ�8a�9/��w��#��5.�Xj_��x��r�Ⱦ�����*�?�T�@��6����+��!����/��s�¿0쿿����Ϩ�:o���t���W�[�,�v!���ʾ�ܖ�@6a�f8/��w�B%��8.�Nn_��{���   �    ^����(��VY��&���E���3��ӿt*�]��+Y��E��\���տk)��+����u��c1[��*�@�����Zӈ�=�J��V �q�����#5���i�|����ʾ^���!�u�B� c����{(��1����E��Y���-�����a�e��~E�$�����;U✾�m���7��
��)�>B!�UK�`����2���   �   4���=P�hㅿY����ƿ�+�L� ���� =���������4�fE�͒ȿ�K������0Q����F��ˣ��j�	B.�|��Dc�����V4��Fh�}��E�r����)l'�ʻ<� �M���X��\�R�Y� BO���>�v�)������s�þ֘��8�m�|�8�Ϝ����2M��j0�sal�"P������   �   ��:��x������kſn�뿒k�n��6l&��]/���2���/�Pp'�� ��h	��S�ZEƿ�쟿_�x���:�̉��������?���׍����	��E+��KZ��+��\��1�;��ﾸ�	;�a0��(�����o���^M�Ѿ㻮������{`���0����,������/�%lB�>!���y��N��   �   DDX������[4���l#�&�0�"A��L��9P�ȱL�6B���1���X��q��η�B���+W�����۾�×�� Q�����i�'�ɽӽ���K#���B�`p����ө���ܼ���;h�ؾ�ݾY�پc�Ͼy�������\��ɯv��I��J!��Y�l�ݽr�ӽ
�o��+�U��	���޾2��   �   QDr�0����xͿ�y��|�
0� G�ֆZ���g���l�~Dh�$0[���G�RU0��q�s�����̿�ß�<Sp�;.�����e���b�����۽8����<��&״��,ڽ�X���&���G�~h��삾Ө���^��:R��i8��sD��*%����m���M�y�,�,���|潞���ӯ��������a"�T�g�qZ������70��   �   g]��M#��#S޿b	�`1$�R�?�8�Y�'p�0�����*��np���Y��L?���#��^�/�ܿ;���o�����<�����z-p�
 ��%׽�؜�$���0���	ڛ��޾�������_$�K`9��*J��:U�2�Y�F�V��M�[=��<)� }��R��˽Q7���㒽sې��Ψ���@/%�g�v��x��"���>��   �   '鉿������t��́,���I�lTf�P�~�	��>�������~�<�e��(I�4�+���p������A����E��q
�h��xy���"�1�սW��Ne���W�t�o��鐽�����ֽ�Y��T��7�Z�#�N]'�I%�w��
���L�vuὲ����	��$K����p�#D~�#t��D)�Sh)�46�����j���xH��   �   �)�����m���!��h/���M���j��������������h���>j�d�L�l?.�d��t�g����g����H�?��|羾3�|�hM$��Iս�ᏽ��Y�\UF�{=X��쁽ట�M��zC⽜ �@����-��V�:��.��B^��˽�%������!q�U_� �r��y��Q⽺�*��큾��¾`���K��   �   �艿ͮ��������,���I�NSf���~�P������-����~�(�e��'I���+�������i���\A����E�q
����wy���"�R�ս���rMe�M�W�(�o��鐽�����ֽ�Y��X��7�\�#�M]'�I%�u�����L�nuὤ����	���J��C�p�TC~��s��](⽟g)��5��E���ջ�xH��   �   S\���!��[Q޿H	�0$���?�,�Y��$p����œ������kp���Y��J?�J�#��]�z�ܿޘ��c����<���𳾆+p���T$׽zל�����ɔ���ٛ��޾�އ�����_$�Q`9��*J��:U�6�Y�H�V��M�[=��<)��|��R���˽�6��P㒽�ڐ��ͨ��	��-%�b�v�>w��� �d�>��   �   PAr�:���svͿ�v��6z��0�XG�ƃZ�d�g�(�l�*Ah�-[�\�G�(S0��o�������̿����PPp��8.�����c���b�1��\۽���;���ִ��,ڽ�X��&���G�~h��삾ר���^��=R��j8��rD��'%����m���M�[�,���+|�����ү�봹�L�彋 ���g�YX������0��   �   �@X�����%����0㿸��� �.�0��A�VL��5P�&�L��B��1����:�#n��˷��?��&(W�n��۾L���I�P����g�d�ɽӽ*��#���B�[p����֩���ܼ���;o�ؾ�ݾ\�پc�Ͼy��񸪾�\����v��I��J!�~Y�$�ݽ��ӽ%�:��քU�d��J޾~/��   �   ��:��x�S����gſ����h�^���h&�:Z/�ȴ2��/��l'�t�f	�EO�vAƿ�響V�x�.�:���$�����/	?���֊������	�-E+��KZ��+��X��1�;��ﾽ�;�e0��(�����o���SM�Ѿͻ������r{`�2�0�"���������,��hB�����u����   �   R���8P�"���Y����ƿ%&�C� �4���9�z��j�����&��?��ȿ�G��Z����P�������$ǣ�̳j�}>.�$���a�����U4��Fh�}��;�r����,l'�λ<�#�M���X��\�T�Y� BO���>�p�)����Д�U�þ������m���8����X���J��f0�
\l�2L��O���   �   �V����(��PY�#��A���.��6ӿ,$����sR�������
տ&$����r��!+[�

*�������ψ�0�J�GS �0��$��"5�V�i��{����ʾY���!�x�B� c����}(��4����E��Z���-�����[�e��~E�u$���b�;✾b�m���7�5	�?'��>!�3K�����i-���   �   ��Ⱦ)��C�*�=�T�������=)��f����,��a�¿鿿����̨��l���r���W��,�����ʾ�ٖ�o1a��4/�jt��!��4.��i_��x��R�Ⱦ����*�@�T�C��9����+��%����/��v�¿1쿿����Ϩ�8o���t���W�O�,�f!���ʾ�ܖ�T5a��6/��u�"��3.��g_��v���   �   �y����ʾP��H�!�?�B�I�b�:��&������C�����Y+��n����e��zE��#�E���;�ޜ���m���7�(�8&��>!�.K�����8/��jY����(�6SY��$��	C���0���ӿ''�����U����Z��7տ'��+���Kt���.[��*�f������ш��J��T �������� 5���i��   �   Ch��z���鿾�m�U��i'�+�<��M�@�X���\�ҖY��=O�f�>���)����\���þ5���~�m��8������J�g0�!]l�OM��*�侶���:P�mᅿ�����ƿ�(濥� ����4;�D��8��j����C�ɐȿCJ��Q���;Q�i��D�侞ɣ��j�j@.����a�����S4��   �   xB+��GZ�C)������;������7�-�;%�B���l�����G�zѾ����.���v`��0���׵��N���,��hB����v��Z��:�¥x�����miſ���
j����bj&��[/���2���/��n'�(��g	��Q��Cƿ�럿��x���:��������S?������C��H�	��   �   -��> ���B�cp����2����ؼ�=�;p�ؾpݾ0�پd�Ͼft������Y��n�v��I��F!�[V�r�ݽ0�ӽ	����U����޾/0��AX�U���*���2㿐���!�x�0�PA�L��7P��L��B���1�����`p��ͷ�XA���*W�E���۾×���P����g㽉�ɽ�ӽ�   �   �Ӵ��(ڽ-V��~&���G�yh��邾����[���N���4��A���!����m�t�M���,�^��Lv�J����ί�Z������ �i�g��X��^���r0� Br�����/wͿ�w���z��	0�pG� �Z���g��l��Bh��.[��G��T0� q�����H�̿Xß��Rp��:.�b���^e��b�t��g۽�����:���   �   X����כ�^۾����T��|\$��\9��&J��6U�ՉY��V�8�L��V=��8)��y�M��˽�2��!��� ؐ��˨�Q�L-%��v�w��� �w�>�m\��"���Q޿�	�d0$�0�?��Y��%p�č�r������ mp�(�Y�L?�>�#�R^�߶ܿ	���V���x�<����񳾆-p����%׽�ל�䵄��   �   ��W���o�~落���r�ֽW����6�a�#�4['��F%�W�� ���J��qὙ�������H��Q�p��?~��q���&��f)�:5����������wH�i艿����������,���I��Sf�l�~�����������`�~���e�h(I�,�+� �����G���B��׸E��q
�����xy���"���ս����Me��   �   u�h��f|��,���涽�۽T���V��\�{�%��))���&�,�o��@	��i⽬5��$����߅�H.x��ˆ�֭�O���\>�����Zھ+� �D�d�F5��C�Ͽ2z�"�#��F��j�w��[W��X8�����3��7���&��V�i�Z�D�"�rG� �Ϳ؍��3b�=x�K׾-f��E�9����Iڥ��~��   �   &�{��2���ɦ��Q˽��������yQ.�S�7�QH;�ֲ8�20�F�"�R�����m�ҽ�p��y钽ص���8���.��������<�^.��	׾��� a�p���I�̿f��=!�B�B��f�����(��o���>h���������Zv��He���A�� ��N�8�ʿ�%��v�^�w����ӾI���X&8��3��F��x���   �   cw������ٽ#��U�59�8kP���b�Qo�!�s��!p��e��LS�G�<�Z#����B���ຽ�1��X���`���ƙ���
8�r����x;���nV��i���ÿs�������8�^�Y�¬y�Պ�6}������7���E���&�y��;Y�8C8�����"�����I"���PT�<���ʾ\H����3�~���6���Y���   �   ��ν4*���L�v<�[#a�ʂ��%��J3�����%竾,f���t���ٔ��Ǆ�1he��T@�R���$ ��bֽ��ý��ν� �_1�|Z���������E�����3��I��@���*�L�F�^�b���z�5���Y����݅��j{��Wc��6G�(*�Z�����?������&D�5�	��c��o�~��-�����j_ǽP���   �   �1��Z/�:�[��5��3��⧼�alԾ�d����TX��V���w�辄�־���ź��Ȯ���%`���3�=�I��k����2*�*�n�?t���1����0�6�r��;���οH��T���0�8�G�"o[���h��m�i��s\���H��u1�Nm�F���_�Ϳ�Ҡ��q���/��@��s���y%k���&�t� �Q�����   �   �7A�L�u����^��������w��%�ʍ.�I�1�!/�`�&��j��t�����þ�7��L�z��%E�T5�m2���A$�,:Y�qb��Eپ��j)R��������ݿ����P�+���;��F�J���F��<�-��������ݿP�������Q�}t� �׾ .��0�V���!�b	��*�����   �   ʷ���f��A!ؾM�z�!��<��lT��ag�s�s�L5x��zt���h�zCV���>���#�\��۾�ѫ�9���F:N�(� n�q1!�p9E��O���J���� �0��*j�cc��]I��q�޿�� �xh�~���3%�\M(��%����������yq࿜r��e����j��T0�� �෾ᭃ���C��V�'?�dy%�K��   �   ����	���?��6��`[�Ac�����
I���v��sw��� ��/A���␿����J�]�\(8����1�澃���z߄�՚M�X+��W"��u4��qc�
-��pIҾ/���=��ut�Eؗ���� �ҿZ�*A �z��jG	��O���yT��Կ'�������+v�(?�ʭ�H�Ҿ�^���<c���3�qE!�;�)�O�K�z���   �   8��|^��(@��6o�cя��������`�˿�#ֿ(ڿ��ֿc�̿��ˣ���@��ىq���A�ě��㾩��+|��D��(��D(�\ZC�;�z��秾��ᾗ[��$@�2o��Ώ��������˿c ֿ��ٿQ�ֿM�̿B��W����>��u�q�C�A�ə�������|��D��(�)F(�0]C���z��ꧾ�   �   ��I>��yt��ڗ����4�ҿ�]�C �b��PI	�hQ�q�}W�Կ_������w.v�L?�O��J�Ҿ�_���=c���3�JD!��)���K�`w��Ἥ�2���<��6�f\[�4^�ϧ��F���s��rt������v>��[���n�����]�f%8�<���|�����݄��M��+��X"��w4��tc��/��MҾ�   �   �0�.j��e���K��v�޿�� �Xj�����5%�nO(��%�P��,��>���s�lt�������j�0V0�� �Y᷾x����C��U�L=�kv%��K�ڴ���b��MؾJ���!�΅<�ghT��\g�k�s�C0x��ut��h�\?V���>���#����۾ϫ�D����7N��(��m�f2!��;E��Q���M���� ��   �   H,R�ԫ������xݿ�	����H�+��;�F�LJ���F�Р<��-�F�������ݿfQ������|�Q�pu�D�׾�.��^�V��!����8(�?��3A�I�u�L���������������%�؉.�V�1�0/�̶&��g�r�ռ�C�þ�4���z��"E�u3��1�>��SB$��<Y�td��Gپ@���   �    s�_=���ο�J�����ޮ0�:�G�\q[�F�h�P�m�0�i��u\��H��v1�<n�����y�Ϳ�Ӡ�6�q�e�/��A��ި���%k�Z�&�K� �uM彭��.�bV/��z[�-2���.��+���'gԾ-_���R������1��Ĉ־���L�������$!`�|�3�������d� 4*���n�Jv���4���0��   �   ���Z5��<��j��V*���F�H�b�Юz�R���n����ޅ�2l{�Yc��7G��*���o�}@��+��'D�r�	�d��L�~���-������\ǽs����ν�#���H���;��a��Ƃ�B"��q/�����)㫾Rb��Mq��~֔�*ń�nce�Q@�P���" ��_ֽ�ý��νM ��`1��[���¾���E��   �   �j���ÿ������@�8���Y�\�y��Պ�~���������������y�r<Y��C8�����"��%���f"���PT�7��ǡʾH��C�3�Ʈ�����V���s��a����ٽ�4R��09��fP���b�b�n�9�s�Ap�� e��HS�Ԡ<�u#�d�����]޺�<0����������E����8�����~z;���oV��   �   C���I�̿�f��>!��B��f�A�����������h��S���>���v��BHe���A�� ��N��ʿ�%���^�"��Z�ӾΎ��%8�,2�\E��<v����{�0��"Ǧ�xN˽�������� O.���7��E;���8�00�}�"���R���~�ҽ�o���蒽�����8���/�����@�<�V/��
׾��"a��   �   �5����Ͽ�z�~�#�0F�n�j�Ow���W��m8������2���6��m&���i���D�h�"� G���ͿX���82b��w�P׾ue��;�9�
��٥���}���h�Be|�9,��=涽�۽�����U�h\�i�%��))���&�2,�����	�nj�[6��⽝�Q���0x��̆��׭��P���]>�Y���[ھֆ ��d��   �   ����u�̿$f��=!�4�B��f������������g��p���q���u��2Ge�ړA� �N�C�ʿ�$��.�^�~��{�Ӿ<����$8�:1�D���u��v�{��/��Ǧ�pN˽��������&O.���7�F;���8�00�y�"���F���l�ҽzo��r蒽>���r8��/��$���}�<��.���	׾l��!a��   �   �i��Mÿ���R����8���Y�ԫy�jԊ�w|������U���i�����y�z:Y�B8����� ������:!��OT���� �ʾG����3������ ��V��vs��!����ٽ�
�5R��09��fP���b�k�n�?�s�Fp�� e��HS�Π<�i#�R��v��޺��/����������_���
8�z����x;����mV��   �   ;��-3��|�忶��6*�J�F��b��z�;���E����܅�rh{��Uc�.5G��*�:����_>������$D�ª	��a��H�~���-�@����Zǽv���νc#���H���;��a��Ƃ�G"��w/��&���-㫾Vb��Nq��{֔�&ń�^ce��P@�)��}" ��^ֽއýРν� ��^1�4Z��J���G���E��   �   �r��:���ο�F��`���0���G�Hm[���h���m��|i��q\���H�t1��k���A�Ϳ	Ѡ�H�q���/��=��%����!k��&��� ��K彄�ｶ-�0V/�wz[�)2���.��2���.gԾ6_�'��R������4��È־���C���꫉�� `�5�3���\���	����1*��n��s���0��0�0��   �   �'R�����Q�ݿ�������+��;��F��J�J�F�̜<� -�8��.��i�ݿ�M��Բ��4�Q�Rr���׾�+��v�V�\�!�J��.'�����2A��u�A���������������%�݉.�Z�1�3/�ζ&��g�r�ʼ�2�þ�4����z�Q"E��2�x0�����?$��8Y�va���پ���   �   x0�V(j��a���G��5�޿�� ��f�����1%�PK(���%�������2��qn��o��/����j��Q0�� ��ܷ�����!�C�0S��;�^u%�K������b��BؾJ���!�҅<�mhT��\g�q�s�H0x��ut��h�[?V���>���#����۾�Ϋ����7N��(�<l��/!��7E��N��nI���� ��   �   ����=��rt�v֗����g�ҿW쿁? �����E	��M����P���ԿE���w��w'v��?�6��b�Ҿ�[���7c�#�3��A!�O�)���K�w���������<��6�h\[�:^�ӧ��F���s��ut������w>��[���l�����]�^%8�2���|�堯��݄��M�1+�V"��s4�3oc�p+��-GҾ�   �   ��ᾔY�7"@��.o��̏����~����˿ֿQ�ٿ��ֿ��̿��e���<����q���A�֖����\����|�zD�S|(�cB(��XC�U�z�n秾��ᾏ[��$@�2o��Ώ���ƀ���˿h ֿ��ٿT�ֿN�̿A��V����>��p�q�;�A�����㾅���|�DD��}(��B(�
XC�+�z��姾�   �   O�����㾂:��6��X[��Y�a���jC���p��sq�������;���ݐ���%�]��!8����w�=����ڄ�i�M��+��T"��s4�Ppc��,��8IҾ!���=��ut�Eؗ�����ҿZ�,A �|��lG	��O���xT��Կ%�������+v�?�����ҾH^��<;c���3�iB!�Å)��K��u���   �   �����_��~ؾ�G���!�A�<�VdT�PXg���s�C+x��pt�1�h��:V��>��#����	۾˫�����2N��(�fj��.!��7E�pO���J���� �0��*j�cc��_I��s�޿�� �|h�����3%�^M(��%����������wq࿙r��a����j��T0�� ��߷�V���J�C�T�l;�t%��K��   �   �/A���u�Q������l��"������%��.�f�1�=/���&�d��n�*��v�þ1���{z��E�[/�$.���?$��8Y�
b��پ��e)R��������ݿ����T�+��;��F�J���F��<�-�������
�ݿP�������Q�jt���׾�-��ݽV���!�d��N&�����   �   |+��R/�v[�^/��z+�����wbԾ�Y羅��L�������辂�־��!���l���>`���3��+���콪�1*�-�n��s���1����0�4�r��;���οH��V��"�0�<�G�$o[���h��m�i��s\���H��u1�Lm�E���_�Ϳ�Ҡ�	�q���/��@��&���|$k�X�&�*� ��J�����   �   !�ν ���E���;��a�
Ă����+��L���2߫�X^��qm���Ҕ������]e�L@���: ��Yֽ��ý��ν ��]1�"Z��y������E�����3��K��B���*�N�F�`�b���z�6���Y����݅��j{��Wc��6G�(*�Z�����?������&D�%�	��c����~��-�j����Zǽ����   �   �q�������ٽ��RO��-9��bP���b���n�U�s�Tp���d�6DS���<��#�,��%�ὢٺ�2,�����I��������	8�:����x;���nV��i���ÿu�������8�^�Y�¬y�Պ�5}������6���E���&�y��;Y�:C8�����"�����H"���PT�4��Сʾ$H��9�3�b���0��jU���   �   ��{�	/���Ŧ�xL˽���d����� M.���7��C;�?�8��-0�:�"���}����ҽ�l���咽����6��U-��q����<�C.��	׾��� a�p���K�̿f��=!�B�B��f�����'��p���>h���������Zv��He���A�� ��N�8�ʿ�%��t�^�s����Ӿ-����%8��2�E��
v���   �   ����b���ť�<�Ƚ~𽟈�f����*�N�3��$7�st4��,���%s�)W��rCͽG���������f�������Q��G�M���������8.��Ux�o���>���02�xY���� ,�������B��쥺��=��I���	��H���W��1����_߿����Lv�̫,�uO꾌��܇J����Ҷ�����   �   �⋽���������޽6-������-��6=��$G���J�;�G�s>��/�Ǫ�{\�l��D��T����p������pD��޷���K��皾���q+��Zt����=�ݿ�@�h>/�U��E~��������(��y���.���������}��!T�(@.��V���ۿ����lr���)�r�澨����H���F{����   �   <���y�ĽƤ��Y���-�&�I��}b��Uv�����p���L���C�w�kkd�;�K��0����w�� �ɽt0���ӭ��ʽ>U�4�F����ڸ޾/h#���h�:柿/Tӿz����&��I��o������-��Wu��q�������BR������Dbo��iI��#&���ҿ�ឿ�(g�@"�V�ܾ�M��. D����[�Ž�A���   �   9��4��R'���L��u��B����
��o1��~���ꬷ�U�$������N�w�)�O��	*��I
�~b�'ӽ߽r<
�B�?�<�t�ξ�����V�|����Yÿ�'��B��2K9�� Z��{z�tS�� ��ś���G��_����{�rgZ��A9�l��fm����¿�璿��U����;̄���!=�^���ڽl�ν�   �   �*��0?��o��3��7���DL;�羪����~�)��������R�辛ϾeS���甾�4r���A�B���d��������Q�7�����纾$B���?�����1񮿬h߿��	��&%��@��M[�r��Հ�W��������r��7\�L}A�V�%��	��C߿l�������?�����������5��.����&��   �   �qR��煾�j���ѾC�����2%�1E4���=�%MA��I>��5�E�&���	�����Ӿ�=��2s���	U���+��^�����1��
k��#��J�뾐5&�pnd�ò���)¿c��f>�b2&� q;��*M��3Y���]��Y��N��y<�'�B���p�u¿����a4d�K�%����J��]i���/�|@�r���)��   �   �8��b��sY뾙H��60��IM��-g�X�{�Ur��%Ն�����^�|���h���N���1�[���}���搏���^���5�L�$�iT.�<uU��b���ȾϹ�X}?�$�~�n`��T.ʿ��"�������*���3��?7�[4���+�j������ ˿��w,�n�?����N�Ǿ�񎾧fT� -�a#���3�8�\��   �   � ��i-��uF�@VF���n�늿:,��é��������6���񉪿�$��j틿<�p���G�Ł �����X���ݏ�Fz^��9���/�=lC�H�v�t?��>�����ʿN���Q���ſ���f1 ����A�J�����������k�U ǿ���b����O���N 徽b���cv���B�]�.�28��]�3玾�   �   �����"�G2Q�O'��r`���t���˿0�ܿz,迺A�+��.�ݿ�̿���r������^�R�~�#������A��A����]T�؈6��a6���S����tw��׳����"�N.Q��$���]���q����˿��ܿ�(�>쿖����ݿ�̿x���3������|�R�V�#������?������\T�0�6�Lc6���S�F���z���   �   ���^�N��������ſb��J3 ��!��C�\�����d��>��n濹ǿ����t�O�X���d���dv���B�$�.��8��]�Q䎾����$(��C�'RF���n�J芿<)��ڿ��΃��{��������"��닿E�p�{�G�C ����8V��܏�ex^�9�B�/�DnC�ߋv�9B��>���   �   V�?��~��b��)1ʿ'���������*���3��A7�N]4���+�&��~��\
�"˿:��.��?�մ���ǾB��fT�<-�"_#���3���\��5���]��T�HE��20�zEM��(g��{��o��l҆�����n�|�H�h��N���1�����y�w����/�^�@�5��$�mU.��wU��d���Ⱦ���   �   �qd������+¿A��@�T4&�8s;�-M�&6Y�"�]�~�Y�� N��{<��'�j���r�w¿̼���5d�U�%�2�꾢J��S]i�<�/��>��o�F�)��lR�d䅾�f���Ѿ�<�����Q{%�A4�4�=��HA��E>��5���&�u
������Ӿo:���p���U�x�+�^����1��k��%������7&��   �   r�����j߿��	�P(%���@��O[��r�I׀������ ����r�v9\��~A�`�%���	�E߿M��������?�k���������6�5����D���$�'�,?��o��/������$G;�美����{�����������'��Ͼ�O��r䔾�/r�C�A�ڢ�c��������7����꺾�C��?��   �   ߟ���[ÿ�)������L9��"Z��}z��T��O������H��Y���@{��hZ��B9���<n��I�¿R蒿?�U�T��;����%!=�Z���ڽJ�ν͙⽹���M'�r�L��u�
?������-��'�������iꮾ!������"�w���O�q*��G
�P_�vӽ�߽=
�ҡ?��󋾒�ξW���V��   �   g矿�UӿZ����&�^�I���o������.��bv��l���^����R��1��� co�2jI�$$&�8��ҿ�ឿ�(g�;"�*�ܾ�M��z�C�����Ž�>��������Ľ'�V�̦-���I��xb��Pv�F�����������v�w�gd�|�K��0�@�����X�ɽ�.��ӭ�c�ʽV���F�D�����޾�i#�j�h��   �   ｧ�O�ݿ2A�*?/� U��F~�L��w���)���y��/��c��ݴ���}��!T� @.��V���ۿ���Tlr���)����%����H���{y���퓽����V������D�޽2+�e��z�-�H4=�."G�h�J���G��p>��/���[��i�IC��b���jp��؈��LE�����A�K��蚾*��r+�8\t��   �   �o���Ῐ���02��Y�[���Y,��翩��B��쥺�x=���������G����W�Z1����9_߿s���Kv��,�bN������J�>���Ѷ�� ����������ĥ���Ƚ��[��.��{�*�:�3��$7��t4��,�C��os��W��%Dͽ�G��i������w���ب��/��m�M�g�����쾄9.�pVx��   �   C���m�ݿ�@�l>/�U��E~�z�����x(��~x��.��s�����Њ}�� T�j?.��U���ۿ�~��Wkr���)���澈����H�<��x��\퓽H���9������:�޽/+�e��~�-�M4=�2"G�m�J���G��p>��/���[��i�(C��6���"p��h����D��.��q�K�	蚾4�(r+�6[t��   �   柿�SӿH��z�&���I�X�o�$����,��yt��x���y���?Q�������`o�rhI��"&�,�6ҿ�����&g��"�\�ܾuL����C������Ž0>�������Ľ�V�ͦ-���I��xb��Pv�K�����������{�w�gd�z�K��0�0��c����ɽ:.��Fҭ��ʽU�+�F�����޾,h#�~�h��   �   ���+Yÿ�&�����\J9��Z�zz�xR���������vF��#����{��eZ�L@9�.��Wk����¿�撿��U�|���;���=����T�ڽ7�ν(�⽋���M'�e�L��u�?������ -��-�������lꮾ!�������w��O�M*�NG
��^�Lӽ�߽�;
���?���
�ξv��g�V��   �   H���L�ug߿��	��%%���@��K[��r��Ԁ�����?���r�j5\�X{A���%���	��A߿���������?�9����������5���8���~#��&��+?��o��/������(G;�羘����{���������(��Ͼ�O��g䔾�/r��A�l��nb�����i��;�7����纾�A���?��   �   �ld�����(¿���<=��0&�8o;�p(M�(1Y���]���Y�`N��w<�('����n�Ks¿¹��G1d���%�v��nG��Yi�~�/�*=�wn���)�XlR�H䅾�f���Ѿ�<�����V{%�A4�:�=��HA��E>��5�&�t
�ރ��{�ӾX:���p��U���+��\�� �8�1�:	k��"��ś�v4&��   �   �{?�Ę~��^��],ʿw����.����*�b�3�:=7��X4���+�X��,����@˿M�(�j�?�l���Ǿ�bT�t-�Y]#���3���\�U5���]��T�FE��20�}EM��(g��{��o��o҆�����r�|�I�h��N���1����ry�T������s�^��5�E�$��R.�RsU��a���Ⱦ����   �   E��n�N�;�]����ſ���/ ����?�8����������Fh�9�ƿ����$�����O����侑_���^v���B�|�.�8��]�䎾����(��C�%RF���n�L芿?)��ݿ��҃��}�������"��닿B�p�v�G�8 ����V���ۏ�Gw^�R9���/�'jC���v��=��͈��   �   ������"�k+Q�#��m[��o����˿D�ܿ4%�U:�߾�5�ݿ��̿N���b��u��z�R�"�#������;��9���cXT�$�6�B_6�4�S�j��,w��������"�K.Q��$���]���q����˿��ܿ�(�>쿚����ݿ�̿x���1������t�R�H�#�v���[?������f[T���6��_6�A�S�=��'u���   �   *���T$���@��NF���n��势�&��򼩿����?����ﲿӃ����R苿j�p�V�G��{ �Z���	R���؏�Ts^��9�^�/�!jC��v�?������ÿN���R���ſ���h1 ����A�L�����������k�S ǿ���^����O��� �Pb��9bv���B�#�.�j8��]�K⎾�   �   33���Z���O뾡B�`/0��AM�G$g�-�{��l���φ�C���%�|�M�h���N���1�U��t���T�����^��5�N�$��Q.�|sU�0b��;Ⱦ���N}?� �~�m`��U.ʿ��$�������*���3��?7�[4���+�j������ ˿��n,�`�?������Ǿ
��dT�r-�]#�"�3�+�\��   �   iR��ᅾVc��ͶѾ�7��x���w%�2=4��=��DA�FA>��5�݃&����}��T�Ӿ,6��gm��U��+�dZ�V����1�w	k�B#���뾂5&�jnd�²���)¿e��h>�d2&�q;��*M��3Y���]��Y��N��y<�'�@���p�u¿����X4d�:�%���꾓I���[i���/�J=��m���)��   �   A$�Y(?��o��,������B;������x�����������o���ϾK�������)r��A�����_�����+����7�
��纾B���?�����1񮿭h߿��	��&%��@��M[�r��Հ�X��������r��7\�L}A�X�%��	��C߿j�������?�։�ʟ������5�R��4���"��   �   ��-��WJ'�:�L��u��;��q쟾����(���|��c���:殾&�������w���O��*��C
�Y�&ӽ�߽�:
��?���>�ξ�����V�|����Yÿ�'��D��4K9�� Z��{z�tS����Ǜ���G��`����{�rgZ��A9�l��fm����¿�璿��U� ���;l���� =�����ڽ��ν�   �   J�����Ľ��T���-��~I�\tb��Kv���������D�w�5bd��K��0�������O�ɽp*��Jϭ���ʽT�r�F�������޾'h#���h�:柿0Tӿ|����&��I��o������-��Vu��p�������BR������Fbo��iI��#&���ҿ�ឿ�(g�7"�4�ܾ�M��n�C�l���Žu=���   �   �ߋ�:
�� ���%�޽�)������-�2=��G���J�A�G�Hn>���/�ۦ�Y�Gf�@�������m��k����B��L����K��皾���q+��Zt����=�ݿ�@�f>/�U��E~��������(��y���.���������}��!T�(@.��V���ۿ����lr���)�d�澍��T�H���y���퓽�   �   Ή�"Ĕ������Խ��������$�WM3�ȋ<��?�:�<���3���%����J���:ֽꭱ�l���.鋽���ý��@�V��O�������6�@�������뿢x�.o;���e��3���ڡ�����x��"���u��������:��|�d��:���^��챿د��
�5�r���yW��z[U�FM�׉��cɕ��   �   ʖ��z`���I½�5��K�y�"�L�6�G�F�W�P��{T��,Q�y;G���7���#��Z�d�VxĽ	���h����*��m�ǽ ��vU��%��lT��$�3��,��^ܯ�|!� �L8��Ua��Y���H�����"�������%�������*��!"��@�`�<�7�8���@�N*��H��3�n�!5����S�(r��VŽ����   �   |����8н����4-���6���S�,n�#W�����`a��`5������4�n��U��8��c�)>��~ҽ�޷��h���yӽ�_���O�:Fx�s+� Jt�ݳ��s�ݿE��S/�IU��~��5��}V��b�����Ҭ���l��I;���~�0�T���.���w�ܿ"��Qbs�G�*�b�Q���iN��*��Aѽ�@���   �   F�@*�J0��W��򀾠����.���綾�k��%�þ�����_��ͨ��X��~����Y���1��g���A^ܽ��轢d�fVH����"�ؾ�d�hra��蚿j�̿r����!�YC�l(g��i��h��������{��ǟ�K+��啅��Rg��SC���!�Js�Qr̿	���7�`���!�׾nđ��G��G�'���4ڽ�   �   =o"��XI���{�����gչ�`ؾ
*�bW��J�6��+w��������ؾĺ�֛��L}�żJ���#��S�I ����N@�a����þX��3�I�H��������k�����-�ƥK�&�h�}Ȁ�y_��O���ϋ��J���#i��L�b.�|��qW��n���Z���I�m���Dþ�{���A?��	���^>
��   �   �|]���\����ܾq��ٮ�6.��=�[�G��+K���G�O>�:�.�7N�xo��ݾ�O��K����^���3��(����g�9�8v�v ��
U��v�.��
p��[��9�˿[���0���/��E�f#Y�2f���j���f�v�Y�b�F�0�/�(���'���̿�a��{�o��l.��������8:u���8����N8��2��   �   ���z¾����|�s�9�o)X�Ps��[��!<���gh�������t�bY�e:����?���X�¾Q��gVi��>�T[,��f6���_��T����Ѿ5���WI�Uم�0���)nԿ+�����z%�2�3���=��A���=��N4��%��~������Կ���A���tI�z��-�Ѿ4��5�^��5�i�+�4=�jEh��   �   ��ƾ���Z�'�d�P�ms{�R2���B��Cp������9���oƻ�bಿ%Τ���d{|���Q��f(�����Ǿ������h���A���7���L�eB��S����6𾒱#�وY��܋�{���E�Ͽ�����t7����8]�<��R�� 3��i񿬍пf���=��[ Z�~�#��v�u���V9���L�f�7��9A�-=h��7���   �   �@��'+�2;\����+���7Ͼ�{�տ��5����������ֿ����8)�����y�\�*�+�����6������^��B?��.?��B^�O���]ʿ�K>�N$+�7\�����<����˾���տ��M��3���M�����Ǧֿχ���&���}��r�\��+����4��e���^�C?��0?�F^��⎾�Ϳ��   �   r�#���Y�Aߋ�I�����Ͽ������9�ز�j_�X��B���4��l�+�пu��&?���Z�?�#��x�ڞ���9���L�#�7�<7A�	9h��4����ƾ4��ҷ'��P�[n{�t/��o?���l��8���ӹ��%û�Pݲ�Yˤ�G���>w|�0�Q�d(�����Ǿ,�����h���A�y�7�ʺL�ED��9���;��   �   [I�[ۅ�����!qԿ�������%���3�6�=�"A�<�=��P4�Ƨ%����|�����Կr
��|���vI������Ѿ���d�^�&�5�[�+��0=��@h�Ŝ��¾�����M�9��$X��Js�Y��D9������e�� ���Dt�L�X��a:������� �¾�N���Si�<
>�![,��g6�/�_��V���Ҿ����   �   p�^����˿\�������
/�l�E�&Y��4f���j�,�f�ƶY�P�F���/�b��)��o̿�b���o��m.�3���į��w:u�$�8�V���5�N�2�w]�J�W��I�ܾ=��,���1.���=�סG� 'K�[�G�:>���.� K��l���ݾ_L��ʹ����^���3��'������9��v��"��xX���.��   �   ޓ������Kn�\����-��K���h��ɀ��`��Ё��2���|���%i�pL�~.�R���X��o��0[��fI����cEþ|��_A?�j���v;
�Lk"�nSI�%�{��𚾲й��ؾ
$�*T�QG�޼��s������8�ؾ����қ��G}��J���#�vR���0	�(P@������þ����I��   �   0ꚿ9�̿����!��ZC�z*g�/k������	���}��dȟ�^,������Tg��TC�\�!��s��r̿v�����`�Z��Z�׾]đ�G��F���潰0ڽO@｜&��E0���W�A蠕�p*��m㶾�f����þ�����[��^ɨ��U��ƪ���Y�+�1�Ze����x\ܽP��Pe�XH����W�ؾxf��ta��   �   �����ݿ�E��T/�zJU�ڮ~��6���W������������lm���;����~���T��.�<����ܿ/"��hbs�B�*��a�
��iN��)�5?ѽ{=�������3н�����)���6� �S��m�hT�������^���2�������n��U�8�7��`�:��8{ҽ�ܷ�.h���yӽ�`�+�O���<z�t+��Kt��   �   Kݯ��"����L8��Va��Z���I��5���"��:���&��N����*��9"��N�`�4�7�&��a@�*���G�f3���4����S�Bq��TŽ� ��p����]���F½2��I�!�"�þ6���F���P��xT�D*Q�)9G���7�Ȯ#�8Y��a��vĽ��������*��U�ǽ ���	U��&��V��@�3�h-���   �   ����E��y��o;�z�e��3���ڡ����y��"���u�����|�������d���:������꿇뱿`���J�5�R����V��KZU�dL�}���Fȕ�&͉�NÔ�֍��:Խ��������$�,M3���<��?�P�<���3��%������D;ֽ����Dᖽ ꋽ8�L�ý˘�x�V�|P�������6��@���   �   �ܯ��!�4�L8��Ua��Y���H��-���!������$��I����)���!��B�`�n�7����y?�d)���F��3����3��ƅS��p�TŽD ��1����]���F½2��I�#�"�Ǿ6���F���P��xT�H*Q�*9G���7�Ʈ#�9Y��a�vĽ߅������p*����ǽv��		U� &��U����3��,���   �   ����3�ݿ�D�fS/��HU�D�~�:5���U��r��� �������k��C:��(�~���T���.� ����ܿ� ��l`s�ڽ*��_����dgN��(��=ѽ�<������3нn����)���6��S��m�lT�������^���2�������n��U�2�7��`��9���zҽPܷ�Vg���xӽ�_���O�ENx�s+��It��   �   O蚿��̿����!�2XC�('g�i��S���U���Ez���ş��)�������Pg�8RC�h�!�6r��p̿������`�h����׾���G�E�5�潒/ڽ�?�j&�pE0���W�@정�u*��t㶾g����þ�����[��aɨ��U��ê���Y��1�!e�ۋ�Q[ܽ~���c��UH�O����ؾ�d��qa��   �   ���������j�����-�J�K�8�h�Lǀ�^���~��M������N!i��
L��.�
��U��l���X��I����BBþ�y���>?������:
��j"�5SI�	�{��𚾳й��ؾ$�/T�WG����s������9�ؾ����қ�|G}�׸J���#��Q���|�|M@������þ���G�I��   �   ,	p��Z����˿k������/��E�!Y�p/f���j���f�ʱY���F� �/�b���$��k̿r_��:�o�j.�3���f���6u�A�8����4���2�w]�+�W��D�ܾ<��.���1.���=�ܡG�&'K�`�G�>>���.� K��l���ݾJL�������^��3��&���ٰ9��v�[��tS��M�.��   �   $VI�؅�����lԿ��������%��3�Z�=�A�\�=�NL4���%� }�������ԿV��9 ���qI�����Ѿ�����^�=�5�{�+��/=��?h������¾ �����N�9��$X��Js�Y��H9������e��#���Ht�K�X��a:������� �¾�N���Ri�	>�<Y,�e6���_�?S����Ѿ����   �   ¯#�_�Y�Iۋ�o�����Ͽ�R���5����[�
��0�� 1�f�k�п���/;����Y���#�r�#����6���{L�Z�7�u5A��7h��4����ƾ&��ͷ'��P�\n{�v/��p?���l��=���׹��)û�Sݲ�[ˤ�G���<w|�,�Q��c(�����ǾԴ����h�2�A���7���L�A������>4��   �   �<� "+��3\�������,ɾ���տ_迕��U���f��Ω�.�ֿ�����#��{��@�\���+�o���0��f��=~^��>?�T,?�<A^��ߎ�ʿ�7>�E$+�7\�����;����˾���տ��Q��9���P�����ɦֿЇ���&���}��n�\�ק+���>4�����h�^��@?��,?�>@^��ގ��ǿ��   �   ��ƾ0��+�'���P�<j{�-���<���i������r��������ٲ�5Ȥ�f���'r|�ڴQ�t`(�����Ǿα����h���A�k�7���L��A��牮��6𾂱#�шY��܋�{���G�Ͽ�����x7����:]�@��T�� 3��i񿪍пg���=��Q Z�k�#�Hv�����8���}L�	�7��4A��5h��2���   �   P����¾����1�ߐ9�� X�+Fs�vV���6��=����b��]���t���X�w]:����"�����¾6K���Mi��>�*W,�d6��_��S��;�Ѿ���WI�Sم�1���*nԿ,�����~%�4�3���=��A���=��N4��%��~������Կ���>���tI�b����Ѿ���e�^�G�5�A�+�.=��<h��   �   �s]��댾4T����ܾ������H..��=���G��"K���G��>�u�.�OG��i�I�ݾ�G��8�����^�6�3��#�w��&�9��v� ���T��f�.��
p��[��;�˿]���2���/��E�j#Y�2f���j���f�v�Y�d�F�0�/�(���'���̿�a��t�o�~l.����������8u���8�����3�s�2��   �   dh"��OI��{��횾�̹�Dؾ��-Q�D�����p��������ؾ\����Λ�A}���J���#��N���0��L@����S�þB��*�I�G��������k�����-�ȥK�(�h�}Ȁ�z_��P���Ћ��K���#i��L�b.�|��qW��n���Z��zI�V���Dþf{��<@?�&�&�N9
��   �   O<��#�B0�$�W��쀾�����&��X߶��b��	�þ����HW��DŨ��Q�������Y�{�1�va�$���VܽN���b�,UH�>���ؾ�d�bra��蚿k�̿r����!�YC�l(g��i��h��������{��ǟ�K+��䕅��Rg��SC���!�Ls�Pr̿���0�`� ����׾đ�hG��E�����-ڽ�   �   @����0нT����&���6��S���m��Q�� ����[���/��a�����n�@U��7�P]��3��vҽeط�<d��"vӽ�^���O��"x�s+��It�ݳ��s�ݿE��S/�IU��~��5��}V��b�����Ҭ���l��I;���~�0�T���.���v�ܿ"��Nbs�>�*��a����hN��)�=>ѽ�;���   �   �����\���D½�/�kH�c�"���6�Q�F��P�<vT��'Q��6G�
�7�l�#�W�
^�nsĽ���[���^(��ěǽ���U�t%��]T�� �3��,��_ܯ�|!�"�L8��Ua��Y���H�����"�������%�������*�� "��@�`�:�7�8���@�O*��H��3�^�5��+�S��q��TŽs ���   